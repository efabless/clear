magic
tech sky130A
magscale 1 2
timestamp 1625784287
<< locali >>
rect 8125 20247 8159 20485
rect 13185 19703 13219 19941
rect 10241 18071 10275 18241
rect 10701 14875 10735 15045
rect 18429 13855 18463 14025
rect 9321 11543 9355 11645
rect 15577 11135 15611 11305
rect 17969 11067 18003 11169
rect 19901 9503 19935 9605
rect 19809 9367 19843 9469
<< viali >>
rect 2605 20553 2639 20587
rect 2973 20553 3007 20587
rect 3341 20553 3375 20587
rect 10241 20553 10275 20587
rect 14289 20553 14323 20587
rect 16221 20553 16255 20587
rect 18153 20553 18187 20587
rect 20729 20553 20763 20587
rect 3617 20485 3651 20519
rect 3893 20485 3927 20519
rect 4445 20485 4479 20519
rect 4813 20485 4847 20519
rect 5273 20485 5307 20519
rect 5917 20485 5951 20519
rect 8033 20485 8067 20519
rect 8125 20485 8159 20519
rect 8861 20485 8895 20519
rect 11529 20485 11563 20519
rect 12541 20485 12575 20519
rect 14565 20485 14599 20519
rect 14933 20485 14967 20519
rect 15301 20485 15335 20519
rect 15669 20485 15703 20519
rect 17049 20485 17083 20519
rect 19717 20485 19751 20519
rect 20453 20485 20487 20519
rect 21557 20485 21591 20519
rect 4261 20417 4295 20451
rect 6837 20417 6871 20451
rect 1869 20349 1903 20383
rect 2053 20349 2087 20383
rect 2697 20349 2731 20383
rect 4629 20349 4663 20383
rect 5733 20349 5767 20383
rect 6101 20349 6135 20383
rect 6561 20349 6595 20383
rect 7205 20349 7239 20383
rect 7389 20349 7423 20383
rect 7849 20349 7883 20383
rect 1501 20281 1535 20315
rect 2145 20281 2179 20315
rect 2329 20281 2363 20315
rect 3065 20281 3099 20315
rect 3433 20281 3467 20315
rect 4077 20281 4111 20315
rect 4997 20281 5031 20315
rect 5457 20281 5491 20315
rect 7665 20281 7699 20315
rect 8493 20417 8527 20451
rect 11069 20417 11103 20451
rect 13185 20417 13219 20451
rect 14013 20417 14047 20451
rect 17877 20417 17911 20451
rect 8217 20349 8251 20383
rect 8677 20349 8711 20383
rect 9229 20349 9263 20383
rect 9505 20349 9539 20383
rect 10149 20349 10183 20383
rect 10609 20349 10643 20383
rect 10977 20349 11011 20383
rect 11437 20349 11471 20383
rect 11713 20349 11747 20383
rect 11897 20349 11931 20383
rect 12173 20349 12207 20383
rect 12725 20349 12759 20383
rect 13093 20349 13127 20383
rect 13645 20349 13679 20383
rect 17509 20349 17543 20383
rect 18429 20349 18463 20383
rect 19901 20349 19935 20383
rect 21373 20349 21407 20383
rect 8953 20281 8987 20315
rect 9873 20281 9907 20315
rect 13461 20281 13495 20315
rect 13829 20281 13863 20315
rect 14197 20281 14231 20315
rect 14749 20281 14783 20315
rect 15117 20281 15151 20315
rect 15485 20281 15519 20315
rect 15853 20281 15887 20315
rect 16129 20281 16163 20315
rect 16497 20281 16531 20315
rect 16681 20281 16715 20315
rect 16865 20281 16899 20315
rect 17325 20281 17359 20315
rect 17693 20281 17727 20315
rect 18061 20281 18095 20315
rect 18613 20281 18647 20315
rect 18797 20281 18831 20315
rect 18981 20281 19015 20315
rect 19165 20281 19199 20315
rect 19349 20281 19383 20315
rect 19533 20281 19567 20315
rect 20269 20281 20303 20315
rect 20637 20281 20671 20315
rect 21005 20281 21039 20315
rect 21189 20281 21223 20315
rect 1593 20213 1627 20247
rect 6285 20213 6319 20247
rect 6745 20213 6779 20247
rect 7021 20213 7055 20247
rect 7573 20213 7607 20247
rect 8125 20213 8159 20247
rect 8401 20213 8435 20247
rect 9413 20213 9447 20247
rect 9689 20213 9723 20247
rect 9965 20213 9999 20247
rect 10425 20213 10459 20247
rect 10793 20213 10827 20247
rect 11253 20213 11287 20247
rect 12081 20213 12115 20247
rect 12357 20213 12391 20247
rect 12909 20213 12943 20247
rect 20085 20213 20119 20247
rect 1869 20009 1903 20043
rect 2329 20009 2363 20043
rect 4629 20009 4663 20043
rect 6377 20009 6411 20043
rect 7297 20009 7331 20043
rect 8125 20009 8159 20043
rect 8493 20009 8527 20043
rect 9137 20009 9171 20043
rect 9597 20009 9631 20043
rect 12541 20009 12575 20043
rect 14105 20009 14139 20043
rect 15393 20009 15427 20043
rect 16313 20009 16347 20043
rect 16957 20009 16991 20043
rect 18613 20009 18647 20043
rect 18705 20009 18739 20043
rect 19165 20009 19199 20043
rect 19441 20009 19475 20043
rect 19901 20009 19935 20043
rect 21189 20009 21223 20043
rect 4813 19941 4847 19975
rect 7941 19941 7975 19975
rect 10210 19941 10244 19975
rect 11897 19941 11931 19975
rect 13185 19941 13219 19975
rect 17233 19941 17267 19975
rect 17601 19941 17635 19975
rect 17785 19941 17819 19975
rect 18061 19941 18095 19975
rect 20637 19941 20671 19975
rect 21373 19941 21407 19975
rect 1593 19873 1627 19907
rect 1961 19873 1995 19907
rect 2145 19873 2179 19907
rect 2421 19873 2455 19907
rect 2873 19873 2907 19907
rect 2982 19873 3016 19907
rect 3249 19873 3283 19907
rect 3709 19873 3743 19907
rect 3893 19873 3927 19907
rect 4169 19873 4203 19907
rect 5181 19873 5215 19907
rect 8585 19873 8619 19907
rect 9505 19873 9539 19907
rect 9965 19873 9999 19907
rect 12357 19873 12391 19907
rect 12817 19873 12851 19907
rect 12909 19873 12943 19907
rect 4997 19805 5031 19839
rect 8401 19805 8435 19839
rect 9689 19805 9723 19839
rect 11621 19805 11655 19839
rect 11805 19805 11839 19839
rect 1409 19737 1443 19771
rect 2605 19737 2639 19771
rect 3433 19737 3467 19771
rect 3525 19737 3559 19771
rect 4077 19737 4111 19771
rect 4445 19737 4479 19771
rect 7757 19737 7791 19771
rect 12265 19737 12299 19771
rect 13645 19873 13679 19907
rect 14749 19873 14783 19907
rect 15209 19873 15243 19907
rect 15485 19873 15519 19907
rect 16129 19873 16163 19907
rect 16405 19873 16439 19907
rect 16773 19873 16807 19907
rect 17417 19873 17451 19907
rect 18245 19873 18279 19907
rect 18429 19873 18463 19907
rect 18889 19873 18923 19907
rect 18981 19873 19015 19907
rect 19257 19873 19291 19907
rect 19717 19873 19751 19907
rect 19993 19873 20027 19907
rect 20361 19873 20395 19907
rect 20821 19873 20855 19907
rect 21005 19873 21039 19907
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 14473 19805 14507 19839
rect 14657 19805 14691 19839
rect 16037 19805 16071 19839
rect 15669 19737 15703 19771
rect 20177 19737 20211 19771
rect 21557 19737 21591 19771
rect 2697 19669 2731 19703
rect 3157 19669 3191 19703
rect 4353 19669 4387 19703
rect 5365 19669 5399 19703
rect 8953 19669 8987 19703
rect 11345 19669 11379 19703
rect 12633 19669 12667 19703
rect 13093 19669 13127 19703
rect 13185 19669 13219 19703
rect 14013 19669 14047 19703
rect 15117 19669 15151 19703
rect 15761 19669 15795 19703
rect 16589 19669 16623 19703
rect 17141 19669 17175 19703
rect 20453 19669 20487 19703
rect 2329 19465 2363 19499
rect 2789 19465 2823 19499
rect 3341 19465 3375 19499
rect 7757 19465 7791 19499
rect 10609 19465 10643 19499
rect 11529 19465 11563 19499
rect 15761 19465 15795 19499
rect 18797 19465 18831 19499
rect 2053 19397 2087 19431
rect 3157 19397 3191 19431
rect 11345 19397 11379 19431
rect 14565 19397 14599 19431
rect 15393 19397 15427 19431
rect 16957 19397 16991 19431
rect 18337 19397 18371 19431
rect 14749 19329 14783 19363
rect 17417 19329 17451 19363
rect 19717 19329 19751 19363
rect 20453 19329 20487 19363
rect 1409 19261 1443 19295
rect 1777 19261 1811 19295
rect 2237 19261 2271 19295
rect 2513 19261 2547 19295
rect 2605 19261 2639 19295
rect 2881 19261 2915 19295
rect 3525 19261 3559 19295
rect 3617 19261 3651 19295
rect 3985 19261 4019 19295
rect 6285 19261 6319 19295
rect 9137 19261 9171 19295
rect 9229 19261 9263 19295
rect 11069 19261 11103 19295
rect 13093 19261 13127 19295
rect 13185 19261 13219 19295
rect 13452 19261 13486 19295
rect 14933 19261 14967 19295
rect 15025 19261 15059 19295
rect 15945 19261 15979 19295
rect 16313 19261 16347 19295
rect 16589 19261 16623 19295
rect 17141 19261 17175 19295
rect 18061 19261 18095 19295
rect 18529 19261 18563 19295
rect 18981 19261 19015 19295
rect 19533 19261 19567 19295
rect 21005 19261 21039 19295
rect 21557 19261 21591 19295
rect 1593 19193 1627 19227
rect 4721 19193 4755 19227
rect 8892 19193 8926 19227
rect 9496 19193 9530 19227
rect 12826 19193 12860 19227
rect 17601 19193 17635 19227
rect 20361 19193 20395 19227
rect 21373 19193 21407 19227
rect 1961 19125 1995 19159
rect 3065 19125 3099 19159
rect 3801 19125 3835 19159
rect 4997 19125 5031 19159
rect 6101 19125 6135 19159
rect 10701 19125 10735 19159
rect 11713 19125 11747 19159
rect 15669 19125 15703 19159
rect 16129 19125 16163 19159
rect 16405 19125 16439 19159
rect 16681 19125 16715 19159
rect 17509 19125 17543 19159
rect 17969 19125 18003 19159
rect 18245 19125 18279 19159
rect 18613 19125 18647 19159
rect 19073 19125 19107 19159
rect 19441 19125 19475 19159
rect 19901 19125 19935 19159
rect 20269 19125 20303 19159
rect 20729 19125 20763 19159
rect 21097 19125 21131 19159
rect 1961 18921 1995 18955
rect 2513 18921 2547 18955
rect 2789 18921 2823 18955
rect 3433 18921 3467 18955
rect 6469 18921 6503 18955
rect 9137 18921 9171 18955
rect 9505 18921 9539 18955
rect 12173 18921 12207 18955
rect 13001 18921 13035 18955
rect 14105 18921 14139 18955
rect 17509 18921 17543 18955
rect 17785 18921 17819 18955
rect 10241 18853 10275 18887
rect 10968 18853 11002 18887
rect 14648 18853 14682 18887
rect 19870 18853 19904 18887
rect 1409 18785 1443 18819
rect 1593 18785 1627 18819
rect 1777 18785 1811 18819
rect 2053 18785 2087 18819
rect 2329 18785 2363 18819
rect 2605 18785 2639 18819
rect 6009 18785 6043 18819
rect 6653 18785 6687 18819
rect 8585 18785 8619 18819
rect 9965 18785 9999 18819
rect 12541 18785 12575 18819
rect 12633 18785 12667 18819
rect 13369 18785 13403 18819
rect 13461 18785 13495 18819
rect 16109 18785 16143 18819
rect 17325 18785 17359 18819
rect 17601 18785 17635 18819
rect 18236 18785 18270 18819
rect 21373 18785 21407 18819
rect 21557 18785 21591 18819
rect 3709 18717 3743 18751
rect 8953 18717 8987 18751
rect 9597 18717 9631 18751
rect 9689 18717 9723 18751
rect 10701 18717 10735 18751
rect 12817 18717 12851 18751
rect 13553 18717 13587 18751
rect 14381 18717 14415 18751
rect 15853 18717 15887 18751
rect 17969 18717 18003 18751
rect 19625 18717 19659 18751
rect 2237 18649 2271 18683
rect 2973 18649 3007 18683
rect 8769 18649 8803 18683
rect 10149 18649 10183 18683
rect 12081 18649 12115 18683
rect 3065 18581 3099 18615
rect 3341 18581 3375 18615
rect 6193 18581 6227 18615
rect 10425 18581 10459 18615
rect 15761 18581 15795 18615
rect 17233 18581 17267 18615
rect 19349 18581 19383 18615
rect 21005 18581 21039 18615
rect 21097 18581 21131 18615
rect 1501 18377 1535 18411
rect 2145 18377 2179 18411
rect 5365 18377 5399 18411
rect 8309 18377 8343 18411
rect 12449 18377 12483 18411
rect 12909 18377 12943 18411
rect 18337 18377 18371 18411
rect 20085 18377 20119 18411
rect 20545 18377 20579 18411
rect 2421 18309 2455 18343
rect 21557 18309 21591 18343
rect 7849 18241 7883 18275
rect 10241 18241 10275 18275
rect 10425 18241 10459 18275
rect 10609 18241 10643 18275
rect 11161 18241 11195 18275
rect 11805 18241 11839 18275
rect 12725 18241 12759 18275
rect 13185 18241 13219 18275
rect 14565 18241 14599 18275
rect 16589 18241 16623 18275
rect 16964 18241 16998 18275
rect 19073 18241 19107 18275
rect 19257 18241 19291 18275
rect 2329 18173 2363 18207
rect 2605 18173 2639 18207
rect 2789 18173 2823 18207
rect 5181 18173 5215 18207
rect 8125 18173 8159 18207
rect 1593 18105 1627 18139
rect 1961 18105 1995 18139
rect 2973 18105 3007 18139
rect 7665 18105 7699 18139
rect 14832 18173 14866 18207
rect 16405 18173 16439 18207
rect 19993 18173 20027 18207
rect 20269 18173 20303 18207
rect 20361 18173 20395 18207
rect 20637 18173 20671 18207
rect 11989 18105 12023 18139
rect 14105 18105 14139 18139
rect 17224 18105 17258 18139
rect 18797 18105 18831 18139
rect 21005 18105 21039 18139
rect 21189 18105 21223 18139
rect 21373 18105 21407 18139
rect 1869 18037 1903 18071
rect 3157 18037 3191 18071
rect 7297 18037 7331 18071
rect 7757 18037 7791 18071
rect 10241 18037 10275 18071
rect 10701 18037 10735 18071
rect 11069 18037 11103 18071
rect 12081 18037 12115 18071
rect 13369 18037 13403 18071
rect 15945 18037 15979 18071
rect 16037 18037 16071 18071
rect 16497 18037 16531 18071
rect 18429 18037 18463 18071
rect 19349 18037 19383 18071
rect 19717 18037 19751 18071
rect 20821 18037 20855 18071
rect 2329 17833 2363 17867
rect 7021 17833 7055 17867
rect 7481 17833 7515 17867
rect 8033 17833 8067 17867
rect 8401 17833 8435 17867
rect 11161 17833 11195 17867
rect 11989 17833 12023 17867
rect 14657 17833 14691 17867
rect 15485 17833 15519 17867
rect 15853 17833 15887 17867
rect 15945 17833 15979 17867
rect 16313 17833 16347 17867
rect 17693 17833 17727 17867
rect 17785 17833 17819 17867
rect 18153 17833 18187 17867
rect 19257 17833 19291 17867
rect 5426 17765 5460 17799
rect 15025 17765 15059 17799
rect 19073 17765 19107 17799
rect 21097 17765 21131 17799
rect 1593 17697 1627 17731
rect 2145 17697 2179 17731
rect 5181 17697 5215 17731
rect 7113 17697 7147 17731
rect 7941 17697 7975 17731
rect 10048 17697 10082 17731
rect 11621 17697 11655 17731
rect 12081 17697 12115 17731
rect 14473 17697 14507 17731
rect 15117 17697 15151 17731
rect 17325 17697 17359 17731
rect 18797 17697 18831 17731
rect 19441 17697 19475 17731
rect 20085 17697 20119 17731
rect 20545 17697 20579 17731
rect 20821 17697 20855 17731
rect 21373 17697 21407 17731
rect 6929 17629 6963 17663
rect 8125 17629 8159 17663
rect 9781 17629 9815 17663
rect 11345 17629 11379 17663
rect 11529 17629 11563 17663
rect 14841 17629 14875 17663
rect 15761 17629 15795 17663
rect 17141 17629 17175 17663
rect 17233 17629 17267 17663
rect 18245 17629 18279 17663
rect 18337 17629 18371 17663
rect 20177 17629 20211 17663
rect 20361 17629 20395 17663
rect 21557 17561 21591 17595
rect 1501 17493 1535 17527
rect 6561 17493 6595 17527
rect 7573 17493 7607 17527
rect 16497 17493 16531 17527
rect 18613 17493 18647 17527
rect 19717 17493 19751 17527
rect 21005 17493 21039 17527
rect 1777 17289 1811 17323
rect 2421 17289 2455 17323
rect 5457 17289 5491 17323
rect 8309 17289 8343 17323
rect 11161 17289 11195 17323
rect 13001 17289 13035 17323
rect 16405 17289 16439 17323
rect 17417 17289 17451 17323
rect 18705 17289 18739 17323
rect 19349 17289 19383 17323
rect 2053 17221 2087 17255
rect 5365 17221 5399 17255
rect 9781 17221 9815 17255
rect 17877 17221 17911 17255
rect 18061 17221 18095 17255
rect 18337 17221 18371 17255
rect 19441 17221 19475 17255
rect 3157 17153 3191 17187
rect 6009 17153 6043 17187
rect 10517 17153 10551 17187
rect 13277 17153 13311 17187
rect 13369 17153 13403 17187
rect 15117 17153 15151 17187
rect 1961 17085 1995 17119
rect 2237 17085 2271 17119
rect 2605 17085 2639 17119
rect 3433 17085 3467 17119
rect 3985 17085 4019 17119
rect 6929 17085 6963 17119
rect 8401 17085 8435 17119
rect 8657 17085 8691 17119
rect 10333 17085 10367 17119
rect 12817 17085 12851 17119
rect 13461 17085 13495 17119
rect 14105 17085 14139 17119
rect 16589 17085 16623 17119
rect 17601 17085 17635 17119
rect 18981 17085 19015 17119
rect 19165 17085 19199 17119
rect 20821 17085 20855 17119
rect 21005 17085 21039 17119
rect 1409 17017 1443 17051
rect 1593 17017 1627 17051
rect 4252 17017 4286 17051
rect 5825 17017 5859 17051
rect 7196 17017 7230 17051
rect 10241 17017 10275 17051
rect 15025 17017 15059 17051
rect 18797 17017 18831 17051
rect 20554 17017 20588 17051
rect 21189 17017 21223 17051
rect 21373 17017 21407 17051
rect 3341 16949 3375 16983
rect 3801 16949 3835 16983
rect 5917 16949 5951 16983
rect 9873 16949 9907 16983
rect 13829 16949 13863 16983
rect 13921 16949 13955 16983
rect 14381 16949 14415 16983
rect 14565 16949 14599 16983
rect 14933 16949 14967 16983
rect 15669 16949 15703 16983
rect 17693 16949 17727 16983
rect 18429 16949 18463 16983
rect 21465 16949 21499 16983
rect 3249 16745 3283 16779
rect 3617 16745 3651 16779
rect 5825 16745 5859 16779
rect 10425 16745 10459 16779
rect 11621 16745 11655 16779
rect 12909 16745 12943 16779
rect 13277 16745 13311 16779
rect 13737 16745 13771 16779
rect 14105 16745 14139 16779
rect 16313 16745 16347 16779
rect 16865 16745 16899 16779
rect 18705 16745 18739 16779
rect 19073 16745 19107 16779
rect 19625 16745 19659 16779
rect 21097 16745 21131 16779
rect 6460 16677 6494 16711
rect 12357 16677 12391 16711
rect 12817 16677 12851 16711
rect 13645 16677 13679 16711
rect 17233 16677 17267 16711
rect 18613 16677 18647 16711
rect 1409 16609 1443 16643
rect 1593 16609 1627 16643
rect 2697 16609 2731 16643
rect 3157 16609 3191 16643
rect 4160 16609 4194 16643
rect 5733 16609 5767 16643
rect 8033 16609 8067 16643
rect 9229 16609 9263 16643
rect 11253 16609 11287 16643
rect 14637 16609 14671 16643
rect 16221 16609 16255 16643
rect 17325 16609 17359 16643
rect 19165 16609 19199 16643
rect 20738 16609 20772 16643
rect 21373 16609 21407 16643
rect 21557 16609 21591 16643
rect 3065 16541 3099 16575
rect 3893 16541 3927 16575
rect 6009 16541 6043 16575
rect 6193 16541 6227 16575
rect 8125 16541 8159 16575
rect 8217 16541 8251 16575
rect 9965 16541 9999 16575
rect 10517 16541 10551 16575
rect 10701 16541 10735 16575
rect 11069 16541 11103 16575
rect 11161 16541 11195 16575
rect 12725 16541 12759 16575
rect 13553 16541 13587 16575
rect 14381 16541 14415 16575
rect 16405 16541 16439 16575
rect 17509 16541 17543 16575
rect 19257 16541 19291 16575
rect 21005 16541 21039 16575
rect 7573 16473 7607 16507
rect 7665 16473 7699 16507
rect 15853 16473 15887 16507
rect 2053 16405 2087 16439
rect 5273 16405 5307 16439
rect 5365 16405 5399 16439
rect 9413 16405 9447 16439
rect 10057 16405 10091 16439
rect 15761 16405 15795 16439
rect 17785 16405 17819 16439
rect 1777 16201 1811 16235
rect 2421 16201 2455 16235
rect 5825 16201 5859 16235
rect 6837 16201 6871 16235
rect 9965 16201 9999 16235
rect 11437 16201 11471 16235
rect 14565 16201 14599 16235
rect 16773 16201 16807 16235
rect 20729 16201 20763 16235
rect 4997 16133 5031 16167
rect 16313 16133 16347 16167
rect 20637 16133 20671 16167
rect 1409 16065 1443 16099
rect 4353 16065 4387 16099
rect 5181 16065 5215 16099
rect 7481 16065 7515 16099
rect 8217 16065 8251 16099
rect 9413 16065 9447 16099
rect 9505 16065 9539 16099
rect 10057 16065 10091 16099
rect 14841 16065 14875 16099
rect 17049 16065 17083 16099
rect 17233 16065 17267 16099
rect 17785 16065 17819 16099
rect 21281 16065 21315 16099
rect 1961 15997 1995 16031
rect 2237 15997 2271 16031
rect 3801 15997 3835 16031
rect 4537 15997 4571 16031
rect 4629 15997 4663 16031
rect 9597 15997 9631 16031
rect 11713 15997 11747 16031
rect 13185 15997 13219 16031
rect 14933 15997 14967 16031
rect 15200 15997 15234 16031
rect 16589 15997 16623 16031
rect 19257 15997 19291 16031
rect 1593 15929 1627 15963
rect 3556 15929 3590 15963
rect 7205 15929 7239 15963
rect 8033 15929 8067 15963
rect 10324 15929 10358 15963
rect 11958 15929 11992 15963
rect 13452 15929 13486 15963
rect 16405 15929 16439 15963
rect 18030 15929 18064 15963
rect 19502 15929 19536 15963
rect 21189 15929 21223 15963
rect 2053 15861 2087 15895
rect 5365 15861 5399 15895
rect 5457 15861 5491 15895
rect 6285 15861 6319 15895
rect 7297 15861 7331 15895
rect 7665 15861 7699 15895
rect 8125 15861 8159 15895
rect 13093 15861 13127 15895
rect 17325 15861 17359 15895
rect 17693 15861 17727 15895
rect 19165 15861 19199 15895
rect 21097 15861 21131 15895
rect 1777 15657 1811 15691
rect 2053 15657 2087 15691
rect 2329 15657 2363 15691
rect 2697 15657 2731 15691
rect 4721 15657 4755 15691
rect 5181 15657 5215 15691
rect 7941 15657 7975 15691
rect 8309 15657 8343 15691
rect 8769 15657 8803 15691
rect 11437 15657 11471 15691
rect 11897 15657 11931 15691
rect 13737 15657 13771 15691
rect 14749 15657 14783 15691
rect 17601 15657 17635 15691
rect 19901 15657 19935 15691
rect 20361 15657 20395 15691
rect 20729 15657 20763 15691
rect 21005 15657 21039 15691
rect 4261 15589 4295 15623
rect 5549 15589 5583 15623
rect 7573 15589 7607 15623
rect 13829 15589 13863 15623
rect 15209 15589 15243 15623
rect 15577 15589 15611 15623
rect 16396 15589 16430 15623
rect 21373 15589 21407 15623
rect 1409 15521 1443 15555
rect 1593 15521 1627 15555
rect 1961 15521 1995 15555
rect 2237 15521 2271 15555
rect 2513 15521 2547 15555
rect 6193 15521 6227 15555
rect 9496 15521 9530 15555
rect 11069 15521 11103 15555
rect 15117 15521 15151 15555
rect 18714 15521 18748 15555
rect 18981 15521 19015 15555
rect 19993 15521 20027 15555
rect 20545 15521 20579 15555
rect 20821 15521 20855 15555
rect 21557 15521 21591 15555
rect 4813 15453 4847 15487
rect 4997 15453 5031 15487
rect 5641 15453 5675 15487
rect 5825 15453 5859 15487
rect 8401 15453 8435 15487
rect 8493 15453 8527 15487
rect 9229 15453 9263 15487
rect 10793 15453 10827 15487
rect 10977 15453 11011 15487
rect 11989 15453 12023 15487
rect 12081 15453 12115 15487
rect 13645 15453 13679 15487
rect 15301 15453 15335 15487
rect 16129 15453 16163 15487
rect 19073 15453 19107 15487
rect 19717 15453 19751 15487
rect 4353 15385 4387 15419
rect 11529 15385 11563 15419
rect 14197 15385 14231 15419
rect 17509 15385 17543 15419
rect 21097 15385 21131 15419
rect 2881 15317 2915 15351
rect 6009 15317 6043 15351
rect 10609 15317 10643 15351
rect 19441 15317 19475 15351
rect 1501 15113 1535 15147
rect 3709 15113 3743 15147
rect 5641 15113 5675 15147
rect 7481 15113 7515 15147
rect 8309 15113 8343 15147
rect 11529 15113 11563 15147
rect 15761 15113 15795 15147
rect 17141 15113 17175 15147
rect 17969 15113 18003 15147
rect 19349 15113 19383 15147
rect 20545 15113 20579 15147
rect 10701 15045 10735 15079
rect 15485 15045 15519 15079
rect 19993 15045 20027 15079
rect 20269 15045 20303 15079
rect 21189 15045 21223 15079
rect 3065 14977 3099 15011
rect 7021 14977 7055 15011
rect 8033 14977 8067 15011
rect 8953 14977 8987 15011
rect 1961 14909 1995 14943
rect 4261 14909 4295 14943
rect 6929 14909 6963 14943
rect 8501 14909 8535 14943
rect 10885 14977 10919 15011
rect 11713 14977 11747 15011
rect 12357 14977 12391 15011
rect 13185 14977 13219 15011
rect 14933 14977 14967 15011
rect 17601 14977 17635 15011
rect 17785 14977 17819 15011
rect 18521 14977 18555 15011
rect 11161 14909 11195 14943
rect 12449 14909 12483 14943
rect 15577 14909 15611 14943
rect 18337 14909 18371 14943
rect 19625 14909 19659 14943
rect 19809 14909 19843 14943
rect 20085 14909 20119 14943
rect 20361 14909 20395 14943
rect 20637 14909 20671 14943
rect 1593 14841 1627 14875
rect 2145 14841 2179 14875
rect 3249 14841 3283 14875
rect 4506 14841 4540 14875
rect 8861 14841 8895 14875
rect 10701 14841 10735 14875
rect 12541 14841 12575 14875
rect 15117 14841 15151 14875
rect 21005 14841 21039 14875
rect 21373 14841 21407 14875
rect 21557 14841 21591 14875
rect 1777 14773 1811 14807
rect 3341 14773 3375 14807
rect 3801 14773 3835 14807
rect 5825 14773 5859 14807
rect 6469 14773 6503 14807
rect 6837 14773 6871 14807
rect 7849 14773 7883 14807
rect 7941 14773 7975 14807
rect 10609 14773 10643 14807
rect 11069 14773 11103 14807
rect 11989 14773 12023 14807
rect 12909 14773 12943 14807
rect 13277 14773 13311 14807
rect 13369 14773 13403 14807
rect 13737 14773 13771 14807
rect 15025 14773 15059 14807
rect 15853 14773 15887 14807
rect 17509 14773 17543 14807
rect 18429 14773 18463 14807
rect 19441 14773 19475 14807
rect 20821 14773 20855 14807
rect 1869 14569 1903 14603
rect 2145 14569 2179 14603
rect 15761 14569 15795 14603
rect 16313 14569 16347 14603
rect 19441 14569 19475 14603
rect 20821 14569 20855 14603
rect 5794 14501 5828 14535
rect 9413 14501 9447 14535
rect 9505 14501 9539 14535
rect 12878 14501 12912 14535
rect 14626 14501 14660 14535
rect 1593 14433 1627 14467
rect 2053 14433 2087 14467
rect 2329 14433 2363 14467
rect 2605 14433 2639 14467
rect 5017 14433 5051 14467
rect 7564 14433 7598 14467
rect 12633 14433 12667 14467
rect 16221 14433 16255 14467
rect 19257 14433 19291 14467
rect 20085 14433 20119 14467
rect 20637 14433 20671 14467
rect 21005 14433 21039 14467
rect 21373 14433 21407 14467
rect 5273 14365 5307 14399
rect 5549 14365 5583 14399
rect 7297 14365 7331 14399
rect 9229 14365 9263 14399
rect 14381 14365 14415 14399
rect 16405 14365 16439 14399
rect 19809 14365 19843 14399
rect 19993 14365 20027 14399
rect 2421 14297 2455 14331
rect 6929 14297 6963 14331
rect 14013 14297 14047 14331
rect 21189 14297 21223 14331
rect 21557 14297 21591 14331
rect 1501 14229 1535 14263
rect 3893 14229 3927 14263
rect 8677 14229 8711 14263
rect 9873 14229 9907 14263
rect 10057 14229 10091 14263
rect 15853 14229 15887 14263
rect 17785 14229 17819 14263
rect 20453 14229 20487 14263
rect 2145 14025 2179 14059
rect 2881 14025 2915 14059
rect 4261 14025 4295 14059
rect 5181 14025 5215 14059
rect 9965 14025 9999 14059
rect 13553 14025 13587 14059
rect 14933 14025 14967 14059
rect 18429 14025 18463 14059
rect 18521 14025 18555 14059
rect 1685 13957 1719 13991
rect 2421 13957 2455 13991
rect 7481 13957 7515 13991
rect 11529 13957 11563 13991
rect 12725 13957 12759 13991
rect 15761 13957 15795 13991
rect 16957 13957 16991 13991
rect 3709 13889 3743 13923
rect 4905 13889 4939 13923
rect 5641 13889 5675 13923
rect 5733 13889 5767 13923
rect 6929 13889 6963 13923
rect 7021 13889 7055 13923
rect 9229 13889 9263 13923
rect 9413 13889 9447 13923
rect 10425 13889 10459 13923
rect 10517 13889 10551 13923
rect 10977 13889 11011 13923
rect 12173 13889 12207 13923
rect 12265 13889 12299 13923
rect 12909 13889 12943 13923
rect 15393 13889 15427 13923
rect 15577 13889 15611 13923
rect 16313 13889 16347 13923
rect 20729 13957 20763 13991
rect 20085 13889 20119 13923
rect 21281 13889 21315 13923
rect 21373 13889 21407 13923
rect 1501 13821 1535 13855
rect 1777 13821 1811 13855
rect 1961 13821 1995 13855
rect 2329 13821 2363 13855
rect 2605 13821 2639 13855
rect 3801 13821 3835 13855
rect 4813 13821 4847 13855
rect 7297 13821 7331 13855
rect 8605 13821 8639 13855
rect 8861 13821 8895 13855
rect 11161 13821 11195 13855
rect 13093 13821 13127 13855
rect 14841 13821 14875 13855
rect 15301 13821 15335 13855
rect 16221 13821 16255 13855
rect 18081 13821 18115 13855
rect 18337 13821 18371 13855
rect 18429 13821 18463 13855
rect 19634 13821 19668 13855
rect 19901 13821 19935 13855
rect 20269 13821 20303 13855
rect 3893 13753 3927 13787
rect 5549 13753 5583 13787
rect 16589 13753 16623 13787
rect 21189 13753 21223 13787
rect 2697 13685 2731 13719
rect 4353 13685 4387 13719
rect 4721 13685 4755 13719
rect 6469 13685 6503 13719
rect 6837 13685 6871 13719
rect 9505 13685 9539 13719
rect 9873 13685 9907 13719
rect 10333 13685 10367 13719
rect 11069 13685 11103 13719
rect 12357 13685 12391 13719
rect 13185 13685 13219 13719
rect 13645 13685 13679 13719
rect 16129 13685 16163 13719
rect 20361 13685 20395 13719
rect 20821 13685 20855 13719
rect 4629 13481 4663 13515
rect 5457 13481 5491 13515
rect 7205 13481 7239 13515
rect 7757 13481 7791 13515
rect 8769 13481 8803 13515
rect 14197 13481 14231 13515
rect 18981 13481 19015 13515
rect 19809 13481 19843 13515
rect 20177 13481 20211 13515
rect 20637 13481 20671 13515
rect 21189 13481 21223 13515
rect 1501 13413 1535 13447
rect 2145 13413 2179 13447
rect 9864 13413 9898 13447
rect 13093 13413 13127 13447
rect 15862 13413 15896 13447
rect 1869 13345 1903 13379
rect 2053 13345 2087 13379
rect 2596 13345 2630 13379
rect 4997 13345 5031 13379
rect 5089 13345 5123 13379
rect 7297 13345 7331 13379
rect 8125 13345 8159 13379
rect 8953 13345 8987 13379
rect 11345 13345 11379 13379
rect 13829 13345 13863 13379
rect 14381 13345 14415 13379
rect 17857 13345 17891 13379
rect 19625 13345 19659 13379
rect 19901 13345 19935 13379
rect 20545 13345 20579 13379
rect 21005 13345 21039 13379
rect 21557 13345 21591 13379
rect 2329 13277 2363 13311
rect 5181 13277 5215 13311
rect 7021 13277 7055 13311
rect 8217 13277 8251 13311
rect 8401 13277 8435 13311
rect 9597 13277 9631 13311
rect 13553 13277 13587 13311
rect 13737 13277 13771 13311
rect 16129 13277 16163 13311
rect 17601 13277 17635 13311
rect 20729 13277 20763 13311
rect 1685 13209 1719 13243
rect 3709 13209 3743 13243
rect 7665 13209 7699 13243
rect 14565 13209 14599 13243
rect 20085 13209 20119 13243
rect 21373 13209 21407 13243
rect 5825 13141 5859 13175
rect 8585 13141 8619 13175
rect 10977 13141 11011 13175
rect 14749 13141 14783 13175
rect 19165 13141 19199 13175
rect 19441 13141 19475 13175
rect 1593 12937 1627 12971
rect 2421 12937 2455 12971
rect 3525 12937 3559 12971
rect 3801 12937 3835 12971
rect 7573 12937 7607 12971
rect 13093 12937 13127 12971
rect 13645 12937 13679 12971
rect 20177 12937 20211 12971
rect 21373 12937 21407 12971
rect 3341 12869 3375 12903
rect 16957 12869 16991 12903
rect 1869 12801 1903 12835
rect 2605 12801 2639 12835
rect 2789 12801 2823 12835
rect 5365 12801 5399 12835
rect 6929 12801 6963 12835
rect 10241 12801 10275 12835
rect 10701 12801 10735 12835
rect 11713 12801 11747 12835
rect 14289 12801 14323 12835
rect 15209 12801 15243 12835
rect 18981 12801 19015 12835
rect 20729 12801 20763 12835
rect 21005 12801 21039 12835
rect 1409 12733 1443 12767
rect 2053 12733 2087 12767
rect 8217 12733 8251 12767
rect 10057 12733 10091 12767
rect 10885 12733 10919 12767
rect 11969 12733 12003 12767
rect 18337 12733 18371 12767
rect 20085 12733 20119 12767
rect 21465 12733 21499 12767
rect 1961 12665 1995 12699
rect 7113 12665 7147 12699
rect 7205 12665 7239 12699
rect 7665 12665 7699 12699
rect 8462 12665 8496 12699
rect 14105 12665 14139 12699
rect 14841 12665 14875 12699
rect 15301 12665 15335 12699
rect 15393 12665 15427 12699
rect 15853 12665 15887 12699
rect 18092 12665 18126 12699
rect 20637 12665 20671 12699
rect 2881 12597 2915 12631
rect 3249 12597 3283 12631
rect 4721 12597 4755 12631
rect 5089 12597 5123 12631
rect 5181 12597 5215 12631
rect 9597 12597 9631 12631
rect 9689 12597 9723 12631
rect 10149 12597 10183 12631
rect 10793 12597 10827 12631
rect 11253 12597 11287 12631
rect 14013 12597 14047 12631
rect 15761 12597 15795 12631
rect 18429 12597 18463 12631
rect 18797 12597 18831 12631
rect 18889 12597 18923 12631
rect 19901 12597 19935 12631
rect 20545 12597 20579 12631
rect 1593 12393 1627 12427
rect 3985 12393 4019 12427
rect 4445 12393 4479 12427
rect 8309 12393 8343 12427
rect 14381 12393 14415 12427
rect 17141 12393 17175 12427
rect 17693 12393 17727 12427
rect 18521 12393 18555 12427
rect 18889 12393 18923 12427
rect 20177 12393 20211 12427
rect 21005 12393 21039 12427
rect 14841 12325 14875 12359
rect 17233 12325 17267 12359
rect 19717 12325 19751 12359
rect 20545 12325 20579 12359
rect 21281 12325 21315 12359
rect 2706 12257 2740 12291
rect 4353 12257 4387 12291
rect 5172 12257 5206 12291
rect 7185 12257 7219 12291
rect 10342 12257 10376 12291
rect 11713 12257 11747 12291
rect 11969 12257 12003 12291
rect 14749 12257 14783 12291
rect 15669 12257 15703 12291
rect 18061 12257 18095 12291
rect 21189 12257 21223 12291
rect 21465 12257 21499 12291
rect 2973 12189 3007 12223
rect 4629 12189 4663 12223
rect 4905 12189 4939 12223
rect 6929 12189 6963 12223
rect 10609 12189 10643 12223
rect 14933 12189 14967 12223
rect 15393 12189 15427 12223
rect 15577 12189 15611 12223
rect 16957 12189 16991 12223
rect 18153 12189 18187 12223
rect 18337 12189 18371 12223
rect 18981 12189 19015 12223
rect 19165 12189 19199 12223
rect 20637 12189 20671 12223
rect 20729 12189 20763 12223
rect 19901 12121 19935 12155
rect 1501 12053 1535 12087
rect 6285 12053 6319 12087
rect 9229 12053 9263 12087
rect 13093 12053 13127 12087
rect 16037 12053 16071 12087
rect 16129 12053 16163 12087
rect 17601 12053 17635 12087
rect 20085 12053 20119 12087
rect 1593 11849 1627 11883
rect 6561 11849 6595 11883
rect 14105 11849 14139 11883
rect 15669 11849 15703 11883
rect 18337 11849 18371 11883
rect 20361 11849 20395 11883
rect 20821 11849 20855 11883
rect 21373 11849 21407 11883
rect 3065 11781 3099 11815
rect 5365 11781 5399 11815
rect 8309 11781 8343 11815
rect 15577 11781 15611 11815
rect 3617 11713 3651 11747
rect 3985 11713 4019 11747
rect 5917 11713 5951 11747
rect 6101 11713 6135 11747
rect 7113 11713 7147 11747
rect 7941 11713 7975 11747
rect 8125 11713 8159 11747
rect 9873 11713 9907 11747
rect 9965 11713 9999 11747
rect 10701 11713 10735 11747
rect 10793 11713 10827 11747
rect 11989 11713 12023 11747
rect 16129 11713 16163 11747
rect 16221 11713 16255 11747
rect 19257 11713 19291 11747
rect 19901 11713 19935 11747
rect 19993 11713 20027 11747
rect 2973 11645 3007 11679
rect 3433 11645 3467 11679
rect 8493 11645 8527 11679
rect 9321 11645 9355 11679
rect 10885 11645 10919 11679
rect 12725 11645 12759 11679
rect 12992 11645 13026 11679
rect 14197 11645 14231 11679
rect 14453 11645 14487 11679
rect 16037 11645 16071 11679
rect 16957 11645 16991 11679
rect 20545 11645 20579 11679
rect 21005 11645 21039 11679
rect 21465 11645 21499 11679
rect 2728 11577 2762 11611
rect 4252 11577 4286 11611
rect 9781 11577 9815 11611
rect 17202 11577 17236 11611
rect 18981 11577 19015 11611
rect 20729 11577 20763 11611
rect 1409 11509 1443 11543
rect 3525 11509 3559 11543
rect 5457 11509 5491 11543
rect 5825 11509 5859 11543
rect 6929 11509 6963 11543
rect 7021 11509 7055 11543
rect 7481 11509 7515 11543
rect 7849 11509 7883 11543
rect 9321 11509 9355 11543
rect 9413 11509 9447 11543
rect 11253 11509 11287 11543
rect 12173 11509 12207 11543
rect 12265 11509 12299 11543
rect 12633 11509 12667 11543
rect 18613 11509 18647 11543
rect 19073 11509 19107 11543
rect 19441 11509 19475 11543
rect 19809 11509 19843 11543
rect 21189 11509 21223 11543
rect 1593 11305 1627 11339
rect 1961 11305 1995 11339
rect 2789 11305 2823 11339
rect 3249 11305 3283 11339
rect 4721 11305 4755 11339
rect 4813 11305 4847 11339
rect 5273 11305 5307 11339
rect 5641 11305 5675 11339
rect 6101 11305 6135 11339
rect 7297 11305 7331 11339
rect 7757 11305 7791 11339
rect 9689 11305 9723 11339
rect 12265 11305 12299 11339
rect 12633 11305 12667 11339
rect 13093 11305 13127 11339
rect 13553 11305 13587 11339
rect 15485 11305 15519 11339
rect 15577 11305 15611 11339
rect 17049 11305 17083 11339
rect 18613 11305 18647 11339
rect 19625 11305 19659 11339
rect 21373 11305 21407 11339
rect 5181 11237 5215 11271
rect 7665 11237 7699 11271
rect 8217 11237 8251 11271
rect 9597 11237 9631 11271
rect 12725 11237 12759 11271
rect 13461 11237 13495 11271
rect 1501 11169 1535 11203
rect 1777 11169 1811 11203
rect 2421 11169 2455 11203
rect 4353 11169 4387 11203
rect 6009 11169 6043 11203
rect 8677 11169 8711 11203
rect 11060 11169 11094 11203
rect 13921 11169 13955 11203
rect 14657 11169 14691 11203
rect 15914 11237 15948 11271
rect 17601 11237 17635 11271
rect 19993 11237 20027 11271
rect 20085 11237 20119 11271
rect 20913 11237 20947 11271
rect 17509 11169 17543 11203
rect 17969 11169 18003 11203
rect 18061 11169 18095 11203
rect 19073 11169 19107 11203
rect 20821 11169 20855 11203
rect 21465 11169 21499 11203
rect 2237 11101 2271 11135
rect 2329 11101 2363 11135
rect 3341 11101 3375 11135
rect 3525 11101 3559 11135
rect 4077 11101 4111 11135
rect 4261 11101 4295 11135
rect 5457 11101 5491 11135
rect 6285 11101 6319 11135
rect 7113 11101 7147 11135
rect 7941 11101 7975 11135
rect 9781 11101 9815 11135
rect 10793 11101 10827 11135
rect 12817 11101 12851 11135
rect 13737 11101 13771 11135
rect 15025 11101 15059 11135
rect 15577 11101 15611 11135
rect 15669 11101 15703 11135
rect 17693 11101 17727 11135
rect 18245 11101 18279 11135
rect 19165 11101 19199 11135
rect 19257 11101 19291 11135
rect 20177 11101 20211 11135
rect 21005 11101 21039 11135
rect 2881 11033 2915 11067
rect 8861 11033 8895 11067
rect 17969 11033 18003 11067
rect 18705 11033 18739 11067
rect 6653 10965 6687 10999
rect 9229 10965 9263 10999
rect 12173 10965 12207 10999
rect 14841 10965 14875 10999
rect 17141 10965 17175 10999
rect 20453 10965 20487 10999
rect 2789 10761 2823 10795
rect 4261 10761 4295 10795
rect 5181 10761 5215 10795
rect 6745 10761 6779 10795
rect 7113 10761 7147 10795
rect 11713 10761 11747 10795
rect 17693 10761 17727 10795
rect 18521 10761 18555 10795
rect 20177 10761 20211 10795
rect 21005 10761 21039 10795
rect 3157 10693 3191 10727
rect 11069 10693 11103 10727
rect 13461 10693 13495 10727
rect 20085 10693 20119 10727
rect 1777 10625 1811 10659
rect 2237 10625 2271 10659
rect 2881 10625 2915 10659
rect 3709 10625 3743 10659
rect 4997 10625 5031 10659
rect 5733 10625 5767 10659
rect 7665 10625 7699 10659
rect 9965 10625 9999 10659
rect 10057 10625 10091 10659
rect 10517 10625 10551 10659
rect 10609 10625 10643 10659
rect 14289 10625 14323 10659
rect 15577 10625 15611 10659
rect 16313 10625 16347 10659
rect 17049 10625 17083 10659
rect 17233 10625 17267 10659
rect 19165 10625 19199 10659
rect 19441 10625 19475 10659
rect 20729 10625 20763 10659
rect 6653 10557 6687 10591
rect 7941 10557 7975 10591
rect 11253 10557 11287 10591
rect 12826 10557 12860 10591
rect 13093 10557 13127 10591
rect 13645 10557 13679 10591
rect 14197 10557 14231 10591
rect 16589 10557 16623 10591
rect 17325 10557 17359 10591
rect 18981 10557 19015 10591
rect 19625 10557 19659 10591
rect 20545 10557 20579 10591
rect 21189 10557 21223 10591
rect 1501 10489 1535 10523
rect 1685 10489 1719 10523
rect 2421 10489 2455 10523
rect 4813 10489 4847 10523
rect 8186 10489 8220 10523
rect 15393 10489 15427 10523
rect 16129 10489 16163 10523
rect 18889 10489 18923 10523
rect 21281 10489 21315 10523
rect 21465 10489 21499 10523
rect 2329 10421 2363 10455
rect 3801 10421 3835 10455
rect 3893 10421 3927 10455
rect 4353 10421 4387 10455
rect 4721 10421 4755 10455
rect 5549 10421 5583 10455
rect 5641 10421 5675 10455
rect 6469 10421 6503 10455
rect 7481 10421 7515 10455
rect 7573 10421 7607 10455
rect 9321 10421 9355 10455
rect 9505 10421 9539 10455
rect 9873 10421 9907 10455
rect 10701 10421 10735 10455
rect 13185 10421 13219 10455
rect 13737 10421 13771 10455
rect 14105 10421 14139 10455
rect 14933 10421 14967 10455
rect 15301 10421 15335 10455
rect 15761 10421 15795 10455
rect 16221 10421 16255 10455
rect 16773 10421 16807 10455
rect 19717 10421 19751 10455
rect 20637 10421 20671 10455
rect 1777 10217 1811 10251
rect 2237 10217 2271 10251
rect 4537 10217 4571 10251
rect 5457 10217 5491 10251
rect 7113 10217 7147 10251
rect 9137 10217 9171 10251
rect 9505 10217 9539 10251
rect 9597 10217 9631 10251
rect 12449 10217 12483 10251
rect 13277 10217 13311 10251
rect 13737 10217 13771 10251
rect 14749 10217 14783 10251
rect 17601 10217 17635 10251
rect 19625 10217 19659 10251
rect 21005 10217 21039 10251
rect 4445 10149 4479 10183
rect 6592 10149 6626 10183
rect 11100 10149 11134 10183
rect 11989 10149 12023 10183
rect 13829 10149 13863 10183
rect 16466 10149 16500 10183
rect 1501 10081 1535 10115
rect 1961 10081 1995 10115
rect 2053 10081 2087 10115
rect 2329 10081 2363 10115
rect 4905 10081 4939 10115
rect 8329 10081 8363 10115
rect 12081 10081 12115 10115
rect 12909 10081 12943 10115
rect 15862 10081 15896 10115
rect 16129 10081 16163 10115
rect 16221 10081 16255 10115
rect 19993 10081 20027 10115
rect 20821 10081 20855 10115
rect 21281 10081 21315 10115
rect 21465 10081 21499 10115
rect 4997 10013 5031 10047
rect 5181 10013 5215 10047
rect 6837 10013 6871 10047
rect 8585 10013 8619 10047
rect 9689 10013 9723 10047
rect 11345 10013 11379 10047
rect 11897 10013 11931 10047
rect 12633 10013 12667 10047
rect 12817 10013 12851 10047
rect 13645 10013 13679 10047
rect 20085 10013 20119 10047
rect 20269 10013 20303 10047
rect 20729 10013 20763 10047
rect 1685 9945 1719 9979
rect 21189 9945 21223 9979
rect 2513 9877 2547 9911
rect 7205 9877 7239 9911
rect 9965 9877 9999 9911
rect 14197 9877 14231 9911
rect 20545 9877 20579 9911
rect 2421 9673 2455 9707
rect 8033 9673 8067 9707
rect 15485 9673 15519 9707
rect 21005 9673 21039 9707
rect 2145 9605 2179 9639
rect 5365 9605 5399 9639
rect 14841 9605 14875 9639
rect 16681 9605 16715 9639
rect 16957 9605 16991 9639
rect 19901 9605 19935 9639
rect 19993 9605 20027 9639
rect 21373 9605 21407 9639
rect 2697 9537 2731 9571
rect 2881 9537 2915 9571
rect 4537 9537 4571 9571
rect 4767 9537 4801 9571
rect 4905 9537 4939 9571
rect 7389 9537 7423 9571
rect 8677 9537 8711 9571
rect 10333 9537 10367 9571
rect 10793 9537 10827 9571
rect 13461 9537 13495 9571
rect 16129 9537 16163 9571
rect 17509 9537 17543 9571
rect 20729 9537 20763 9571
rect 2329 9469 2363 9503
rect 2605 9469 2639 9503
rect 3157 9469 3191 9503
rect 7481 9469 7515 9503
rect 8401 9469 8435 9503
rect 10149 9469 10183 9503
rect 10977 9469 11011 9503
rect 11897 9469 11931 9503
rect 13728 9469 13762 9503
rect 15853 9469 15887 9503
rect 17417 9469 17451 9503
rect 19717 9469 19751 9503
rect 19809 9469 19843 9503
rect 19901 9469 19935 9503
rect 20637 9469 20671 9503
rect 21189 9469 21223 9503
rect 21557 9469 21591 9503
rect 1501 9401 1535 9435
rect 1869 9401 1903 9435
rect 2053 9401 2087 9435
rect 4997 9401 5031 9435
rect 8493 9401 8527 9435
rect 10241 9401 10275 9435
rect 10885 9401 10919 9435
rect 12164 9401 12198 9435
rect 16497 9401 16531 9435
rect 17325 9401 17359 9435
rect 19472 9401 19506 9435
rect 1593 9333 1627 9367
rect 7573 9333 7607 9367
rect 7941 9333 7975 9367
rect 9781 9333 9815 9367
rect 11345 9333 11379 9367
rect 13277 9333 13311 9367
rect 15945 9333 15979 9367
rect 18337 9333 18371 9367
rect 19809 9333 19843 9367
rect 20177 9333 20211 9367
rect 20545 9333 20579 9367
rect 1593 9129 1627 9163
rect 3893 9129 3927 9163
rect 5457 9129 5491 9163
rect 5825 9129 5859 9163
rect 6193 9129 6227 9163
rect 6285 9129 6319 9163
rect 9321 9129 9355 9163
rect 9781 9129 9815 9163
rect 10425 9129 10459 9163
rect 10885 9129 10919 9163
rect 13369 9129 13403 9163
rect 13737 9129 13771 9163
rect 14473 9129 14507 9163
rect 15577 9129 15611 9163
rect 16037 9129 16071 9163
rect 18981 9129 19015 9163
rect 21005 9129 21039 9163
rect 21373 9129 21407 9163
rect 7113 9061 7147 9095
rect 9137 9061 9171 9095
rect 9689 9061 9723 9095
rect 13829 9061 13863 9095
rect 19901 9061 19935 9095
rect 20085 9061 20119 9095
rect 1409 8993 1443 9027
rect 1952 8993 1986 9027
rect 4261 8993 4295 9027
rect 5365 8993 5399 9027
rect 8401 8993 8435 9027
rect 10793 8993 10827 9027
rect 13021 8993 13055 9027
rect 15669 8993 15703 9027
rect 17049 8993 17083 9027
rect 17601 8993 17635 9027
rect 17868 8993 17902 9027
rect 20545 8993 20579 9027
rect 21465 8993 21499 9027
rect 1685 8925 1719 8959
rect 4353 8925 4387 8959
rect 4445 8925 4479 8959
rect 5641 8925 5675 8959
rect 6377 8925 6411 8959
rect 7205 8925 7239 8959
rect 7389 8925 7423 8959
rect 8493 8925 8527 8959
rect 8585 8925 8619 8959
rect 9873 8925 9907 8959
rect 10977 8925 11011 8959
rect 11345 8925 11379 8959
rect 13277 8925 13311 8959
rect 13921 8925 13955 8959
rect 15485 8925 15519 8959
rect 16865 8925 16899 8959
rect 16957 8925 16991 8959
rect 20637 8925 20671 8959
rect 20729 8925 20763 8959
rect 3065 8857 3099 8891
rect 4997 8857 5031 8891
rect 7665 8857 7699 8891
rect 8953 8857 8987 8891
rect 6745 8789 6779 8823
rect 8033 8789 8067 8823
rect 11897 8789 11931 8823
rect 15209 8789 15243 8823
rect 16313 8789 16347 8823
rect 16589 8789 16623 8823
rect 17417 8789 17451 8823
rect 20177 8789 20211 8823
rect 2421 8585 2455 8619
rect 3341 8585 3375 8619
rect 4169 8585 4203 8619
rect 5457 8585 5491 8619
rect 6285 8585 6319 8619
rect 7941 8585 7975 8619
rect 19349 8585 19383 8619
rect 20085 8585 20119 8619
rect 21005 8585 21039 8619
rect 21373 8585 21407 8619
rect 3249 8517 3283 8551
rect 8401 8517 8435 8551
rect 18521 8517 18555 8551
rect 1869 8449 1903 8483
rect 2605 8449 2639 8483
rect 2789 8449 2823 8483
rect 3893 8449 3927 8483
rect 4905 8449 4939 8483
rect 5641 8449 5675 8483
rect 5825 8449 5859 8483
rect 17141 8449 17175 8483
rect 18705 8449 18739 8483
rect 18889 8449 18923 8483
rect 19993 8449 20027 8483
rect 20637 8449 20671 8483
rect 2053 8381 2087 8415
rect 2881 8381 2915 8415
rect 3801 8381 3835 8415
rect 6561 8381 6595 8415
rect 9514 8381 9548 8415
rect 9781 8381 9815 8415
rect 19809 8381 19843 8415
rect 1961 8313 1995 8347
rect 6806 8313 6840 8347
rect 17386 8313 17420 8347
rect 19625 8313 19659 8347
rect 21097 8313 21131 8347
rect 21465 8313 21499 8347
rect 1409 8245 1443 8279
rect 3709 8245 3743 8279
rect 4997 8245 5031 8279
rect 5089 8245 5123 8279
rect 5917 8245 5951 8279
rect 18981 8245 19015 8279
rect 20453 8245 20487 8279
rect 20545 8245 20579 8279
rect 2053 8041 2087 8075
rect 17969 8041 18003 8075
rect 18337 8041 18371 8075
rect 19717 8041 19751 8075
rect 20177 8041 20211 8075
rect 20545 8041 20579 8075
rect 21373 8041 21407 8075
rect 1501 7973 1535 8007
rect 1685 7973 1719 8007
rect 4988 7973 5022 8007
rect 6438 7973 6472 8007
rect 8125 7973 8159 8007
rect 8585 7973 8619 8007
rect 20085 7973 20119 8007
rect 1777 7905 1811 7939
rect 3177 7905 3211 7939
rect 4261 7905 4295 7939
rect 4721 7905 4755 7939
rect 8033 7905 8067 7939
rect 20729 7905 20763 7939
rect 21189 7905 21223 7939
rect 21465 7905 21499 7939
rect 3433 7837 3467 7871
rect 4353 7837 4387 7871
rect 4537 7837 4571 7871
rect 6193 7837 6227 7871
rect 8217 7837 8251 7871
rect 17693 7837 17727 7871
rect 17877 7837 17911 7871
rect 20361 7837 20395 7871
rect 20913 7837 20947 7871
rect 6101 7769 6135 7803
rect 7665 7769 7699 7803
rect 21005 7769 21039 7803
rect 1961 7701 1995 7735
rect 3893 7701 3927 7735
rect 7573 7701 7607 7735
rect 2145 7497 2179 7531
rect 16957 7497 16991 7531
rect 20821 7497 20855 7531
rect 1685 7429 1719 7463
rect 2881 7429 2915 7463
rect 4905 7429 4939 7463
rect 7389 7429 7423 7463
rect 1777 7361 1811 7395
rect 3525 7361 3559 7395
rect 3893 7361 3927 7395
rect 5457 7361 5491 7395
rect 8769 7361 8803 7395
rect 21373 7361 21407 7395
rect 5365 7293 5399 7327
rect 18337 7293 18371 7327
rect 19349 7293 19383 7327
rect 1501 7225 1535 7259
rect 1961 7225 1995 7259
rect 3249 7225 3283 7259
rect 8524 7225 8558 7259
rect 18092 7225 18126 7259
rect 19616 7225 19650 7259
rect 3341 7157 3375 7191
rect 5273 7157 5307 7191
rect 5733 7157 5767 7191
rect 20729 7157 20763 7191
rect 21189 7157 21223 7191
rect 21281 7157 21315 7191
rect 5273 6953 5307 6987
rect 21005 6953 21039 6987
rect 1501 6817 1535 6851
rect 2982 6817 3016 6851
rect 3249 6817 3283 6851
rect 19625 6817 19659 6851
rect 19892 6817 19926 6851
rect 21189 6817 21223 6851
rect 21465 6817 21499 6851
rect 5365 6749 5399 6783
rect 5457 6749 5491 6783
rect 4905 6681 4939 6715
rect 21281 6681 21315 6715
rect 1593 6613 1627 6647
rect 1869 6613 1903 6647
rect 21281 6341 21315 6375
rect 20729 6273 20763 6307
rect 1501 6137 1535 6171
rect 1685 6137 1719 6171
rect 21189 6137 21223 6171
rect 21465 6137 21499 6171
rect 1777 6069 1811 6103
rect 1593 5865 1627 5899
rect 21097 5865 21131 5899
rect 21373 5865 21407 5899
rect 1409 5729 1443 5763
rect 1685 5729 1719 5763
rect 20729 5729 20763 5763
rect 21281 5729 21315 5763
rect 21557 5729 21591 5763
rect 20545 5661 20579 5695
rect 20637 5661 20671 5695
rect 20177 5525 20211 5559
rect 1685 5253 1719 5287
rect 21281 5253 21315 5287
rect 1501 5117 1535 5151
rect 1777 5117 1811 5151
rect 21189 5117 21223 5151
rect 21465 5117 21499 5151
rect 1593 4777 1627 4811
rect 21373 4777 21407 4811
rect 1961 4709 1995 4743
rect 1409 4641 1443 4675
rect 1685 4641 1719 4675
rect 2145 4641 2179 4675
rect 20821 4641 20855 4675
rect 21281 4641 21315 4675
rect 21557 4641 21591 4675
rect 21005 4573 21039 4607
rect 1869 4505 1903 4539
rect 21097 4505 21131 4539
rect 1593 4233 1627 4267
rect 1409 4029 1443 4063
rect 1685 4029 1719 4063
rect 21281 4029 21315 4063
rect 21557 4029 21591 4063
rect 21373 3893 21407 3927
rect 1593 3689 1627 3723
rect 21373 3689 21407 3723
rect 1409 3553 1443 3587
rect 1869 3553 1903 3587
rect 21097 3553 21131 3587
rect 21557 3553 21591 3587
rect 20913 3485 20947 3519
rect 1685 3417 1719 3451
rect 2237 3417 2271 3451
rect 21281 3417 21315 3451
rect 2053 3349 2087 3383
rect 20637 3349 20671 3383
rect 2145 3145 2179 3179
rect 4813 3145 4847 3179
rect 5641 3145 5675 3179
rect 20821 3145 20855 3179
rect 21373 3145 21407 3179
rect 1593 3077 1627 3111
rect 20545 3077 20579 3111
rect 1409 2941 1443 2975
rect 1685 2941 1719 2975
rect 1961 2941 1995 2975
rect 4997 2941 5031 2975
rect 5825 2941 5859 2975
rect 20729 2941 20763 2975
rect 21005 2941 21039 2975
rect 21281 2941 21315 2975
rect 21557 2941 21591 2975
rect 2237 2873 2271 2907
rect 2513 2873 2547 2907
rect 15393 2873 15427 2907
rect 15577 2873 15611 2907
rect 20361 2873 20395 2907
rect 1869 2805 1903 2839
rect 2697 2805 2731 2839
rect 21097 2805 21131 2839
rect 1869 2601 1903 2635
rect 2145 2601 2179 2635
rect 2973 2601 3007 2635
rect 3341 2601 3375 2635
rect 11529 2601 11563 2635
rect 16129 2601 16163 2635
rect 20177 2601 20211 2635
rect 20453 2601 20487 2635
rect 21005 2601 21039 2635
rect 7113 2533 7147 2567
rect 1409 2465 1443 2499
rect 1685 2465 1719 2499
rect 1961 2465 1995 2499
rect 2329 2465 2363 2499
rect 3249 2465 3283 2499
rect 3525 2465 3559 2499
rect 3893 2465 3927 2499
rect 11713 2465 11747 2499
rect 11897 2465 11931 2499
rect 16313 2465 16347 2499
rect 19717 2465 19751 2499
rect 20361 2465 20395 2499
rect 20637 2465 20671 2499
rect 20913 2465 20947 2499
rect 21189 2465 21223 2499
rect 21465 2465 21499 2499
rect 3617 2397 3651 2431
rect 20085 2397 20119 2431
rect 3065 2329 3099 2363
rect 6929 2329 6963 2363
rect 20729 2329 20763 2363
rect 1593 2261 1627 2295
rect 16405 2261 16439 2295
rect 21373 2261 21407 2295
<< metal1 >>
rect 2682 20884 2688 20936
rect 2740 20924 2746 20936
rect 3510 20924 3516 20936
rect 2740 20896 3516 20924
rect 2740 20884 2746 20896
rect 3510 20884 3516 20896
rect 3568 20884 3574 20936
rect 1854 20816 1860 20868
rect 1912 20856 1918 20868
rect 3418 20856 3424 20868
rect 1912 20828 3424 20856
rect 1912 20816 1918 20828
rect 3418 20816 3424 20828
rect 3476 20816 3482 20868
rect 1394 20748 1400 20800
rect 1452 20788 1458 20800
rect 2866 20788 2872 20800
rect 1452 20760 2872 20788
rect 1452 20748 1458 20760
rect 2866 20748 2872 20760
rect 2924 20748 2930 20800
rect 17954 20748 17960 20800
rect 18012 20788 18018 20800
rect 21450 20788 21456 20800
rect 18012 20760 21456 20788
rect 18012 20748 18018 20760
rect 21450 20748 21456 20760
rect 21508 20748 21514 20800
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 2593 20587 2651 20593
rect 2593 20553 2605 20587
rect 2639 20584 2651 20587
rect 2774 20584 2780 20596
rect 2639 20556 2780 20584
rect 2639 20553 2651 20556
rect 2593 20547 2651 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 2958 20584 2964 20596
rect 2919 20556 2964 20584
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 3326 20584 3332 20596
rect 3287 20556 3332 20584
rect 3326 20544 3332 20556
rect 3384 20544 3390 20596
rect 3786 20544 3792 20596
rect 3844 20584 3850 20596
rect 9398 20584 9404 20596
rect 3844 20556 9404 20584
rect 3844 20544 3850 20556
rect 9398 20544 9404 20556
rect 9456 20544 9462 20596
rect 9950 20544 9956 20596
rect 10008 20584 10014 20596
rect 10229 20587 10287 20593
rect 10229 20584 10241 20587
rect 10008 20556 10241 20584
rect 10008 20544 10014 20556
rect 1486 20476 1492 20528
rect 1544 20516 1550 20528
rect 3605 20519 3663 20525
rect 3605 20516 3617 20519
rect 1544 20488 3617 20516
rect 1544 20476 1550 20488
rect 3605 20485 3617 20488
rect 3651 20485 3663 20519
rect 3878 20516 3884 20528
rect 3839 20488 3884 20516
rect 3605 20479 3663 20485
rect 3878 20476 3884 20488
rect 3936 20476 3942 20528
rect 4338 20476 4344 20528
rect 4396 20516 4402 20528
rect 4433 20519 4491 20525
rect 4433 20516 4445 20519
rect 4396 20488 4445 20516
rect 4396 20476 4402 20488
rect 4433 20485 4445 20488
rect 4479 20485 4491 20519
rect 4798 20516 4804 20528
rect 4759 20488 4804 20516
rect 4433 20479 4491 20485
rect 4798 20476 4804 20488
rect 4856 20476 4862 20528
rect 5258 20516 5264 20528
rect 5219 20488 5264 20516
rect 5258 20476 5264 20488
rect 5316 20476 5322 20528
rect 5905 20519 5963 20525
rect 5905 20485 5917 20519
rect 5951 20516 5963 20519
rect 6730 20516 6736 20528
rect 5951 20488 6736 20516
rect 5951 20485 5963 20488
rect 5905 20479 5963 20485
rect 6730 20476 6736 20488
rect 6788 20476 6794 20528
rect 7466 20476 7472 20528
rect 7524 20516 7530 20528
rect 8021 20519 8079 20525
rect 8021 20516 8033 20519
rect 7524 20488 8033 20516
rect 7524 20476 7530 20488
rect 8021 20485 8033 20488
rect 8067 20485 8079 20519
rect 8021 20479 8079 20485
rect 8113 20519 8171 20525
rect 8113 20485 8125 20519
rect 8159 20516 8171 20519
rect 8849 20519 8907 20525
rect 8159 20488 8800 20516
rect 8159 20485 8171 20488
rect 8113 20479 8171 20485
rect 2590 20448 2596 20460
rect 1872 20420 2596 20448
rect 1026 20340 1032 20392
rect 1084 20380 1090 20392
rect 1872 20389 1900 20420
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 2774 20408 2780 20460
rect 2832 20448 2838 20460
rect 4249 20451 4307 20457
rect 4249 20448 4261 20451
rect 2832 20420 4261 20448
rect 2832 20408 2838 20420
rect 4249 20417 4261 20420
rect 4295 20417 4307 20451
rect 6825 20451 6883 20457
rect 6825 20448 6837 20451
rect 4249 20411 4307 20417
rect 5736 20420 6837 20448
rect 5736 20392 5764 20420
rect 6825 20417 6837 20420
rect 6871 20417 6883 20451
rect 8481 20451 8539 20457
rect 8481 20448 8493 20451
rect 6825 20411 6883 20417
rect 7392 20420 8493 20448
rect 7392 20392 7420 20420
rect 8481 20417 8493 20420
rect 8527 20417 8539 20451
rect 8772 20448 8800 20488
rect 8849 20485 8861 20519
rect 8895 20516 8907 20519
rect 10042 20516 10048 20528
rect 8895 20488 10048 20516
rect 8895 20485 8907 20488
rect 8849 20479 8907 20485
rect 10042 20476 10048 20488
rect 10100 20476 10106 20528
rect 9858 20448 9864 20460
rect 8772 20420 9864 20448
rect 8481 20411 8539 20417
rect 9858 20408 9864 20420
rect 9916 20408 9922 20460
rect 1857 20383 1915 20389
rect 1857 20380 1869 20383
rect 1084 20352 1869 20380
rect 1084 20340 1090 20352
rect 1857 20349 1869 20352
rect 1903 20349 1915 20383
rect 1857 20343 1915 20349
rect 2041 20383 2099 20389
rect 2041 20349 2053 20383
rect 2087 20380 2099 20383
rect 2685 20383 2743 20389
rect 2087 20352 2636 20380
rect 2087 20349 2099 20352
rect 2041 20343 2099 20349
rect 566 20272 572 20324
rect 624 20312 630 20324
rect 1486 20312 1492 20324
rect 624 20284 1492 20312
rect 624 20272 630 20284
rect 1486 20272 1492 20284
rect 1544 20272 1550 20324
rect 2130 20312 2136 20324
rect 2091 20284 2136 20312
rect 2130 20272 2136 20284
rect 2188 20272 2194 20324
rect 2317 20315 2375 20321
rect 2317 20281 2329 20315
rect 2363 20312 2375 20315
rect 2498 20312 2504 20324
rect 2363 20284 2504 20312
rect 2363 20281 2375 20284
rect 2317 20275 2375 20281
rect 2498 20272 2504 20284
rect 2556 20272 2562 20324
rect 1581 20247 1639 20253
rect 1581 20213 1593 20247
rect 1627 20244 1639 20247
rect 2222 20244 2228 20256
rect 1627 20216 2228 20244
rect 1627 20213 1639 20216
rect 1581 20207 1639 20213
rect 2222 20204 2228 20216
rect 2280 20204 2286 20256
rect 2608 20244 2636 20352
rect 2685 20349 2697 20383
rect 2731 20380 2743 20383
rect 3878 20380 3884 20392
rect 2731 20352 3884 20380
rect 2731 20349 2743 20352
rect 2685 20343 2743 20349
rect 3878 20340 3884 20352
rect 3936 20340 3942 20392
rect 4617 20383 4675 20389
rect 4617 20349 4629 20383
rect 4663 20380 4675 20383
rect 5074 20380 5080 20392
rect 4663 20352 5080 20380
rect 4663 20349 4675 20352
rect 4617 20343 4675 20349
rect 5074 20340 5080 20352
rect 5132 20340 5138 20392
rect 5718 20380 5724 20392
rect 5679 20352 5724 20380
rect 5718 20340 5724 20352
rect 5776 20340 5782 20392
rect 6086 20380 6092 20392
rect 6047 20352 6092 20380
rect 6086 20340 6092 20352
rect 6144 20340 6150 20392
rect 6546 20380 6552 20392
rect 6507 20352 6552 20380
rect 6546 20340 6552 20352
rect 6604 20340 6610 20392
rect 7006 20340 7012 20392
rect 7064 20380 7070 20392
rect 7193 20383 7251 20389
rect 7193 20380 7205 20383
rect 7064 20352 7205 20380
rect 7064 20340 7070 20352
rect 7193 20349 7205 20352
rect 7239 20349 7251 20383
rect 7374 20380 7380 20392
rect 7335 20352 7380 20380
rect 7193 20343 7251 20349
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 7834 20380 7840 20392
rect 7795 20352 7840 20380
rect 7834 20340 7840 20352
rect 7892 20340 7898 20392
rect 8202 20380 8208 20392
rect 8163 20352 8208 20380
rect 8202 20340 8208 20352
rect 8260 20340 8266 20392
rect 8662 20380 8668 20392
rect 8623 20352 8668 20380
rect 8662 20340 8668 20352
rect 8720 20340 8726 20392
rect 9122 20340 9128 20392
rect 9180 20380 9186 20392
rect 9217 20383 9275 20389
rect 9217 20380 9229 20383
rect 9180 20352 9229 20380
rect 9180 20340 9186 20352
rect 9217 20349 9229 20352
rect 9263 20349 9275 20383
rect 9490 20380 9496 20392
rect 9451 20352 9496 20380
rect 9217 20343 9275 20349
rect 9490 20340 9496 20352
rect 9548 20340 9554 20392
rect 10152 20389 10180 20556
rect 10229 20553 10241 20556
rect 10275 20553 10287 20587
rect 10229 20547 10287 20553
rect 11974 20544 11980 20596
rect 12032 20584 12038 20596
rect 13354 20584 13360 20596
rect 12032 20556 13360 20584
rect 12032 20544 12038 20556
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 14277 20587 14335 20593
rect 14277 20553 14289 20587
rect 14323 20584 14335 20587
rect 15930 20584 15936 20596
rect 14323 20556 15936 20584
rect 14323 20553 14335 20556
rect 14277 20547 14335 20553
rect 15930 20544 15936 20556
rect 15988 20544 15994 20596
rect 16209 20587 16267 20593
rect 16209 20553 16221 20587
rect 16255 20584 16267 20587
rect 17954 20584 17960 20596
rect 16255 20556 17960 20584
rect 16255 20553 16267 20556
rect 16209 20547 16267 20553
rect 17954 20544 17960 20556
rect 18012 20544 18018 20596
rect 18141 20587 18199 20593
rect 18141 20553 18153 20587
rect 18187 20584 18199 20587
rect 18874 20584 18880 20596
rect 18187 20556 18880 20584
rect 18187 20553 18199 20556
rect 18141 20547 18199 20553
rect 18874 20544 18880 20556
rect 18932 20544 18938 20596
rect 20162 20584 20168 20596
rect 18984 20556 20168 20584
rect 11517 20519 11575 20525
rect 11517 20485 11529 20519
rect 11563 20516 11575 20519
rect 12158 20516 12164 20528
rect 11563 20488 12164 20516
rect 11563 20485 11575 20488
rect 11517 20479 11575 20485
rect 12158 20476 12164 20488
rect 12216 20476 12222 20528
rect 12250 20476 12256 20528
rect 12308 20516 12314 20528
rect 12529 20519 12587 20525
rect 12529 20516 12541 20519
rect 12308 20488 12541 20516
rect 12308 20476 12314 20488
rect 12529 20485 12541 20488
rect 12575 20485 12587 20519
rect 12529 20479 12587 20485
rect 12802 20476 12808 20528
rect 12860 20516 12866 20528
rect 13722 20516 13728 20528
rect 12860 20488 13728 20516
rect 12860 20476 12866 20488
rect 13722 20476 13728 20488
rect 13780 20476 13786 20528
rect 14182 20476 14188 20528
rect 14240 20516 14246 20528
rect 14553 20519 14611 20525
rect 14553 20516 14565 20519
rect 14240 20488 14565 20516
rect 14240 20476 14246 20488
rect 14553 20485 14565 20488
rect 14599 20485 14611 20519
rect 14553 20479 14611 20485
rect 14642 20476 14648 20528
rect 14700 20516 14706 20528
rect 14921 20519 14979 20525
rect 14921 20516 14933 20519
rect 14700 20488 14933 20516
rect 14700 20476 14706 20488
rect 14921 20485 14933 20488
rect 14967 20485 14979 20519
rect 14921 20479 14979 20485
rect 15194 20476 15200 20528
rect 15252 20516 15258 20528
rect 15289 20519 15347 20525
rect 15289 20516 15301 20519
rect 15252 20488 15301 20516
rect 15252 20476 15258 20488
rect 15289 20485 15301 20488
rect 15335 20485 15347 20519
rect 15289 20479 15347 20485
rect 15470 20476 15476 20528
rect 15528 20516 15534 20528
rect 15657 20519 15715 20525
rect 15657 20516 15669 20519
rect 15528 20488 15669 20516
rect 15528 20476 15534 20488
rect 15657 20485 15669 20488
rect 15703 20485 15715 20519
rect 15657 20479 15715 20485
rect 17037 20519 17095 20525
rect 17037 20485 17049 20519
rect 17083 20516 17095 20519
rect 18984 20516 19012 20556
rect 20162 20544 20168 20556
rect 20220 20544 20226 20596
rect 20530 20544 20536 20596
rect 20588 20584 20594 20596
rect 20717 20587 20775 20593
rect 20717 20584 20729 20587
rect 20588 20556 20729 20584
rect 20588 20544 20594 20556
rect 20717 20553 20729 20556
rect 20763 20553 20775 20587
rect 20717 20547 20775 20553
rect 19702 20516 19708 20528
rect 17083 20488 19012 20516
rect 19663 20488 19708 20516
rect 17083 20485 17095 20488
rect 17037 20479 17095 20485
rect 19702 20476 19708 20488
rect 19760 20476 19766 20528
rect 20438 20516 20444 20528
rect 20399 20488 20444 20516
rect 20438 20476 20444 20488
rect 20496 20476 20502 20528
rect 21545 20519 21603 20525
rect 21545 20485 21557 20519
rect 21591 20516 21603 20519
rect 22738 20516 22744 20528
rect 21591 20488 22744 20516
rect 21591 20485 21603 20488
rect 21545 20479 21603 20485
rect 22738 20476 22744 20488
rect 22796 20476 22802 20528
rect 11057 20451 11115 20457
rect 11057 20448 11069 20451
rect 10612 20420 11069 20448
rect 10137 20383 10195 20389
rect 10137 20349 10149 20383
rect 10183 20349 10195 20383
rect 10137 20343 10195 20349
rect 10410 20340 10416 20392
rect 10468 20380 10474 20392
rect 10612 20389 10640 20420
rect 11057 20417 11069 20420
rect 11103 20417 11115 20451
rect 13173 20451 13231 20457
rect 13173 20448 13185 20451
rect 11057 20411 11115 20417
rect 11440 20420 13185 20448
rect 10597 20383 10655 20389
rect 10597 20380 10609 20383
rect 10468 20352 10609 20380
rect 10468 20340 10474 20352
rect 10597 20349 10609 20352
rect 10643 20349 10655 20383
rect 10597 20343 10655 20349
rect 10778 20340 10784 20392
rect 10836 20380 10842 20392
rect 10965 20383 11023 20389
rect 10965 20380 10977 20383
rect 10836 20352 10977 20380
rect 10836 20340 10842 20352
rect 10965 20349 10977 20352
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 11238 20340 11244 20392
rect 11296 20380 11302 20392
rect 11440 20389 11468 20420
rect 13173 20417 13185 20420
rect 13219 20417 13231 20451
rect 13173 20411 13231 20417
rect 14001 20451 14059 20457
rect 14001 20417 14013 20451
rect 14047 20448 14059 20451
rect 16298 20448 16304 20460
rect 14047 20420 16304 20448
rect 14047 20417 14059 20420
rect 14001 20411 14059 20417
rect 16298 20408 16304 20420
rect 16356 20408 16362 20460
rect 17865 20451 17923 20457
rect 17865 20417 17877 20451
rect 17911 20448 17923 20451
rect 19334 20448 19340 20460
rect 17911 20420 19340 20448
rect 17911 20417 17923 20420
rect 17865 20411 17923 20417
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 11425 20383 11483 20389
rect 11425 20380 11437 20383
rect 11296 20352 11437 20380
rect 11296 20340 11302 20352
rect 11425 20349 11437 20352
rect 11471 20349 11483 20383
rect 11425 20343 11483 20349
rect 11701 20383 11759 20389
rect 11701 20349 11713 20383
rect 11747 20349 11759 20383
rect 11701 20343 11759 20349
rect 3050 20312 3056 20324
rect 3011 20284 3056 20312
rect 3050 20272 3056 20284
rect 3108 20272 3114 20324
rect 3326 20272 3332 20324
rect 3384 20312 3390 20324
rect 3421 20315 3479 20321
rect 3421 20312 3433 20315
rect 3384 20284 3433 20312
rect 3384 20272 3390 20284
rect 3421 20281 3433 20284
rect 3467 20281 3479 20315
rect 3694 20312 3700 20324
rect 3421 20275 3479 20281
rect 3528 20284 3700 20312
rect 3528 20244 3556 20284
rect 3694 20272 3700 20284
rect 3752 20272 3758 20324
rect 4062 20312 4068 20324
rect 4023 20284 4068 20312
rect 4062 20272 4068 20284
rect 4120 20272 4126 20324
rect 4890 20272 4896 20324
rect 4948 20312 4954 20324
rect 4985 20315 5043 20321
rect 4985 20312 4997 20315
rect 4948 20284 4997 20312
rect 4948 20272 4954 20284
rect 4985 20281 4997 20284
rect 5031 20281 5043 20315
rect 4985 20275 5043 20281
rect 5445 20315 5503 20321
rect 5445 20281 5457 20315
rect 5491 20312 5503 20315
rect 6564 20312 6592 20340
rect 7653 20315 7711 20321
rect 7653 20312 7665 20315
rect 5491 20284 6500 20312
rect 6564 20284 7665 20312
rect 5491 20281 5503 20284
rect 5445 20275 5503 20281
rect 2608 20216 3556 20244
rect 3602 20204 3608 20256
rect 3660 20244 3666 20256
rect 4246 20244 4252 20256
rect 3660 20216 4252 20244
rect 3660 20204 3666 20216
rect 4246 20204 4252 20216
rect 4304 20204 4310 20256
rect 6270 20244 6276 20256
rect 6231 20216 6276 20244
rect 6270 20204 6276 20216
rect 6328 20204 6334 20256
rect 6472 20244 6500 20284
rect 7653 20281 7665 20284
rect 7699 20281 7711 20315
rect 7852 20312 7880 20340
rect 8941 20315 8999 20321
rect 8941 20312 8953 20315
rect 7852 20284 8953 20312
rect 7653 20275 7711 20281
rect 8941 20281 8953 20284
rect 8987 20281 8999 20315
rect 8941 20275 8999 20281
rect 9861 20315 9919 20321
rect 9861 20281 9873 20315
rect 9907 20312 9919 20315
rect 11716 20312 11744 20343
rect 11790 20340 11796 20392
rect 11848 20380 11854 20392
rect 11885 20383 11943 20389
rect 11885 20380 11897 20383
rect 11848 20352 11897 20380
rect 11848 20340 11854 20352
rect 11885 20349 11897 20352
rect 11931 20349 11943 20383
rect 11885 20343 11943 20349
rect 12066 20340 12072 20392
rect 12124 20380 12130 20392
rect 12161 20383 12219 20389
rect 12161 20380 12173 20383
rect 12124 20352 12173 20380
rect 12124 20340 12130 20352
rect 12161 20349 12173 20352
rect 12207 20349 12219 20383
rect 12161 20343 12219 20349
rect 12526 20340 12532 20392
rect 12584 20380 12590 20392
rect 12710 20380 12716 20392
rect 12584 20352 12716 20380
rect 12584 20340 12590 20352
rect 12710 20340 12716 20352
rect 12768 20340 12774 20392
rect 12894 20340 12900 20392
rect 12952 20380 12958 20392
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 12952 20352 13093 20380
rect 12952 20340 12958 20352
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 13633 20383 13691 20389
rect 13633 20349 13645 20383
rect 13679 20380 13691 20383
rect 16758 20380 16764 20392
rect 13679 20352 16764 20380
rect 13679 20349 13691 20352
rect 13633 20343 13691 20349
rect 16758 20340 16764 20352
rect 16816 20340 16822 20392
rect 17497 20383 17555 20389
rect 17497 20349 17509 20383
rect 17543 20380 17555 20383
rect 18414 20380 18420 20392
rect 17543 20352 18276 20380
rect 18375 20352 18420 20380
rect 17543 20349 17555 20352
rect 17497 20343 17555 20349
rect 11974 20312 11980 20324
rect 9907 20284 11980 20312
rect 9907 20281 9919 20284
rect 9861 20275 9919 20281
rect 11974 20272 11980 20284
rect 12032 20272 12038 20324
rect 13449 20315 13507 20321
rect 13449 20281 13461 20315
rect 13495 20281 13507 20315
rect 13449 20275 13507 20281
rect 13817 20315 13875 20321
rect 13817 20281 13829 20315
rect 13863 20312 13875 20315
rect 13998 20312 14004 20324
rect 13863 20284 14004 20312
rect 13863 20281 13875 20284
rect 13817 20275 13875 20281
rect 6638 20244 6644 20256
rect 6472 20216 6644 20244
rect 6638 20204 6644 20216
rect 6696 20204 6702 20256
rect 6733 20247 6791 20253
rect 6733 20213 6745 20247
rect 6779 20244 6791 20247
rect 6914 20244 6920 20256
rect 6779 20216 6920 20244
rect 6779 20213 6791 20216
rect 6733 20207 6791 20213
rect 6914 20204 6920 20216
rect 6972 20204 6978 20256
rect 7009 20247 7067 20253
rect 7009 20213 7021 20247
rect 7055 20244 7067 20247
rect 7190 20244 7196 20256
rect 7055 20216 7196 20244
rect 7055 20213 7067 20216
rect 7009 20207 7067 20213
rect 7190 20204 7196 20216
rect 7248 20204 7254 20256
rect 7561 20247 7619 20253
rect 7561 20213 7573 20247
rect 7607 20244 7619 20247
rect 8113 20247 8171 20253
rect 8113 20244 8125 20247
rect 7607 20216 8125 20244
rect 7607 20213 7619 20216
rect 7561 20207 7619 20213
rect 8113 20213 8125 20216
rect 8159 20213 8171 20247
rect 8113 20207 8171 20213
rect 8389 20247 8447 20253
rect 8389 20213 8401 20247
rect 8435 20244 8447 20247
rect 8754 20244 8760 20256
rect 8435 20216 8760 20244
rect 8435 20213 8447 20216
rect 8389 20207 8447 20213
rect 8754 20204 8760 20216
rect 8812 20204 8818 20256
rect 9030 20204 9036 20256
rect 9088 20244 9094 20256
rect 9401 20247 9459 20253
rect 9401 20244 9413 20247
rect 9088 20216 9413 20244
rect 9088 20204 9094 20216
rect 9401 20213 9413 20216
rect 9447 20213 9459 20247
rect 9674 20244 9680 20256
rect 9635 20216 9680 20244
rect 9401 20207 9459 20213
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 9950 20244 9956 20256
rect 9911 20216 9956 20244
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 10042 20204 10048 20256
rect 10100 20244 10106 20256
rect 10413 20247 10471 20253
rect 10413 20244 10425 20247
rect 10100 20216 10425 20244
rect 10100 20204 10106 20216
rect 10413 20213 10425 20216
rect 10459 20213 10471 20247
rect 10413 20207 10471 20213
rect 10502 20204 10508 20256
rect 10560 20244 10566 20256
rect 10781 20247 10839 20253
rect 10781 20244 10793 20247
rect 10560 20216 10793 20244
rect 10560 20204 10566 20216
rect 10781 20213 10793 20216
rect 10827 20213 10839 20247
rect 10781 20207 10839 20213
rect 11146 20204 11152 20256
rect 11204 20244 11210 20256
rect 11241 20247 11299 20253
rect 11241 20244 11253 20247
rect 11204 20216 11253 20244
rect 11204 20204 11210 20216
rect 11241 20213 11253 20216
rect 11287 20213 11299 20247
rect 11241 20207 11299 20213
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 12069 20247 12127 20253
rect 12069 20244 12081 20247
rect 11940 20216 12081 20244
rect 11940 20204 11946 20216
rect 12069 20213 12081 20216
rect 12115 20213 12127 20247
rect 12342 20244 12348 20256
rect 12303 20216 12348 20244
rect 12069 20207 12127 20213
rect 12342 20204 12348 20216
rect 12400 20204 12406 20256
rect 12618 20204 12624 20256
rect 12676 20244 12682 20256
rect 12897 20247 12955 20253
rect 12897 20244 12909 20247
rect 12676 20216 12909 20244
rect 12676 20204 12682 20216
rect 12897 20213 12909 20216
rect 12943 20213 12955 20247
rect 13464 20244 13492 20275
rect 13998 20272 14004 20284
rect 14056 20272 14062 20324
rect 14185 20315 14243 20321
rect 14185 20281 14197 20315
rect 14231 20281 14243 20315
rect 14185 20275 14243 20281
rect 14090 20244 14096 20256
rect 13464 20216 14096 20244
rect 12897 20207 12955 20213
rect 14090 20204 14096 20216
rect 14148 20204 14154 20256
rect 14200 20244 14228 20275
rect 14274 20272 14280 20324
rect 14332 20312 14338 20324
rect 14737 20315 14795 20321
rect 14737 20312 14749 20315
rect 14332 20284 14749 20312
rect 14332 20272 14338 20284
rect 14737 20281 14749 20284
rect 14783 20281 14795 20315
rect 14737 20275 14795 20281
rect 14826 20272 14832 20324
rect 14884 20312 14890 20324
rect 15105 20315 15163 20321
rect 15105 20312 15117 20315
rect 14884 20284 15117 20312
rect 14884 20272 14890 20284
rect 15105 20281 15117 20284
rect 15151 20281 15163 20315
rect 15470 20312 15476 20324
rect 15431 20284 15476 20312
rect 15105 20275 15163 20281
rect 15470 20272 15476 20284
rect 15528 20272 15534 20324
rect 15838 20312 15844 20324
rect 15799 20284 15844 20312
rect 15838 20272 15844 20284
rect 15896 20272 15902 20324
rect 15930 20272 15936 20324
rect 15988 20312 15994 20324
rect 16117 20315 16175 20321
rect 16117 20312 16129 20315
rect 15988 20284 16129 20312
rect 15988 20272 15994 20284
rect 16117 20281 16129 20284
rect 16163 20281 16175 20315
rect 16117 20275 16175 20281
rect 16206 20272 16212 20324
rect 16264 20312 16270 20324
rect 16485 20315 16543 20321
rect 16485 20312 16497 20315
rect 16264 20284 16497 20312
rect 16264 20272 16270 20284
rect 16485 20281 16497 20284
rect 16531 20281 16543 20315
rect 16666 20312 16672 20324
rect 16627 20284 16672 20312
rect 16485 20275 16543 20281
rect 16666 20272 16672 20284
rect 16724 20272 16730 20324
rect 16853 20315 16911 20321
rect 16853 20281 16865 20315
rect 16899 20281 16911 20315
rect 16853 20275 16911 20281
rect 17313 20315 17371 20321
rect 17313 20281 17325 20315
rect 17359 20281 17371 20315
rect 17313 20275 17371 20281
rect 16022 20244 16028 20256
rect 14200 20216 16028 20244
rect 16022 20204 16028 20216
rect 16080 20204 16086 20256
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 16868 20244 16896 20275
rect 16816 20216 16896 20244
rect 17328 20244 17356 20275
rect 17678 20272 17684 20324
rect 17736 20312 17742 20324
rect 18049 20315 18107 20321
rect 17736 20284 17781 20312
rect 17736 20272 17742 20284
rect 18049 20281 18061 20315
rect 18095 20312 18107 20315
rect 18138 20312 18144 20324
rect 18095 20284 18144 20312
rect 18095 20281 18107 20284
rect 18049 20275 18107 20281
rect 18138 20272 18144 20284
rect 18196 20272 18202 20324
rect 18248 20312 18276 20352
rect 18414 20340 18420 20352
rect 18472 20340 18478 20392
rect 19610 20380 19616 20392
rect 18524 20352 19616 20380
rect 18524 20312 18552 20352
rect 19610 20340 19616 20352
rect 19668 20340 19674 20392
rect 19702 20340 19708 20392
rect 19760 20380 19766 20392
rect 19889 20383 19947 20389
rect 19889 20380 19901 20383
rect 19760 20352 19901 20380
rect 19760 20340 19766 20352
rect 19889 20349 19901 20352
rect 19935 20349 19947 20383
rect 19889 20343 19947 20349
rect 20714 20340 20720 20392
rect 20772 20380 20778 20392
rect 21361 20383 21419 20389
rect 21361 20380 21373 20383
rect 20772 20352 21373 20380
rect 20772 20340 20778 20352
rect 21361 20349 21373 20352
rect 21407 20349 21419 20383
rect 21361 20343 21419 20349
rect 18248 20284 18552 20312
rect 18598 20272 18604 20324
rect 18656 20312 18662 20324
rect 18785 20315 18843 20321
rect 18656 20284 18701 20312
rect 18656 20272 18662 20284
rect 18785 20281 18797 20315
rect 18831 20281 18843 20315
rect 18966 20312 18972 20324
rect 18927 20284 18972 20312
rect 18785 20275 18843 20281
rect 18690 20244 18696 20256
rect 17328 20216 18696 20244
rect 16816 20204 16822 20216
rect 18690 20204 18696 20216
rect 18748 20204 18754 20256
rect 18800 20244 18828 20275
rect 18966 20272 18972 20284
rect 19024 20272 19030 20324
rect 19150 20312 19156 20324
rect 19111 20284 19156 20312
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 19337 20315 19395 20321
rect 19337 20281 19349 20315
rect 19383 20281 19395 20315
rect 19337 20275 19395 20281
rect 19242 20244 19248 20256
rect 18800 20216 19248 20244
rect 19242 20204 19248 20216
rect 19300 20204 19306 20256
rect 19352 20244 19380 20275
rect 19426 20272 19432 20324
rect 19484 20312 19490 20324
rect 19521 20315 19579 20321
rect 19521 20312 19533 20315
rect 19484 20284 19533 20312
rect 19484 20272 19490 20284
rect 19521 20281 19533 20284
rect 19567 20281 19579 20315
rect 19521 20275 19579 20281
rect 20257 20315 20315 20321
rect 20257 20281 20269 20315
rect 20303 20281 20315 20315
rect 20257 20275 20315 20281
rect 19794 20244 19800 20256
rect 19352 20216 19800 20244
rect 19794 20204 19800 20216
rect 19852 20204 19858 20256
rect 20073 20247 20131 20253
rect 20073 20213 20085 20247
rect 20119 20244 20131 20247
rect 20272 20244 20300 20275
rect 20438 20272 20444 20324
rect 20496 20312 20502 20324
rect 20625 20315 20683 20321
rect 20625 20312 20637 20315
rect 20496 20284 20637 20312
rect 20496 20272 20502 20284
rect 20625 20281 20637 20284
rect 20671 20281 20683 20315
rect 20990 20312 20996 20324
rect 20951 20284 20996 20312
rect 20625 20275 20683 20281
rect 20990 20272 20996 20284
rect 21048 20272 21054 20324
rect 21174 20312 21180 20324
rect 21135 20284 21180 20312
rect 21174 20272 21180 20284
rect 21232 20272 21238 20324
rect 20119 20216 20300 20244
rect 20119 20213 20131 20216
rect 20073 20207 20131 20213
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 1854 20040 1860 20052
rect 1815 20012 1860 20040
rect 1854 20000 1860 20012
rect 1912 20000 1918 20052
rect 2317 20043 2375 20049
rect 2317 20009 2329 20043
rect 2363 20040 2375 20043
rect 4062 20040 4068 20052
rect 2363 20012 4068 20040
rect 2363 20009 2375 20012
rect 2317 20003 2375 20009
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4617 20043 4675 20049
rect 4617 20040 4629 20043
rect 4212 20012 4629 20040
rect 4212 20000 4218 20012
rect 4617 20009 4629 20012
rect 4663 20009 4675 20043
rect 4617 20003 4675 20009
rect 6086 20000 6092 20052
rect 6144 20040 6150 20052
rect 6365 20043 6423 20049
rect 6365 20040 6377 20043
rect 6144 20012 6377 20040
rect 6144 20000 6150 20012
rect 6365 20009 6377 20012
rect 6411 20009 6423 20043
rect 6365 20003 6423 20009
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 7285 20043 7343 20049
rect 7285 20040 7297 20043
rect 7064 20012 7297 20040
rect 7064 20000 7070 20012
rect 7285 20009 7297 20012
rect 7331 20009 7343 20043
rect 7285 20003 7343 20009
rect 8113 20043 8171 20049
rect 8113 20009 8125 20043
rect 8159 20040 8171 20043
rect 8202 20040 8208 20052
rect 8159 20012 8208 20040
rect 8159 20009 8171 20012
rect 8113 20003 8171 20009
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 8481 20043 8539 20049
rect 8481 20009 8493 20043
rect 8527 20040 8539 20043
rect 9125 20043 9183 20049
rect 9125 20040 9137 20043
rect 8527 20012 9137 20040
rect 8527 20009 8539 20012
rect 8481 20003 8539 20009
rect 9125 20009 9137 20012
rect 9171 20009 9183 20043
rect 9125 20003 9183 20009
rect 9398 20000 9404 20052
rect 9456 20040 9462 20052
rect 9585 20043 9643 20049
rect 9585 20040 9597 20043
rect 9456 20012 9597 20040
rect 9456 20000 9462 20012
rect 9585 20009 9597 20012
rect 9631 20009 9643 20043
rect 9585 20003 9643 20009
rect 9950 20000 9956 20052
rect 10008 20040 10014 20052
rect 10870 20040 10876 20052
rect 10008 20012 10876 20040
rect 10008 20000 10014 20012
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 12529 20043 12587 20049
rect 12529 20009 12541 20043
rect 12575 20009 12587 20043
rect 12529 20003 12587 20009
rect 2038 19932 2044 19984
rect 2096 19972 2102 19984
rect 2096 19944 2452 19972
rect 2096 19932 2102 19944
rect 1578 19904 1584 19916
rect 1539 19876 1584 19904
rect 1578 19864 1584 19876
rect 1636 19864 1642 19916
rect 1946 19904 1952 19916
rect 1907 19876 1952 19904
rect 1946 19864 1952 19876
rect 2004 19864 2010 19916
rect 2130 19904 2136 19916
rect 2091 19876 2136 19904
rect 2130 19864 2136 19876
rect 2188 19864 2194 19916
rect 2424 19913 2452 19944
rect 2498 19932 2504 19984
rect 2556 19972 2562 19984
rect 4801 19975 4859 19981
rect 4801 19972 4813 19975
rect 2556 19944 4813 19972
rect 2556 19932 2562 19944
rect 2409 19907 2467 19913
rect 2409 19873 2421 19907
rect 2455 19873 2467 19907
rect 2409 19867 2467 19873
rect 2861 19907 2919 19913
rect 2861 19873 2873 19907
rect 2907 19873 2919 19907
rect 2861 19867 2919 19873
rect 2970 19907 3028 19913
rect 2970 19873 2982 19907
rect 3016 19873 3028 19907
rect 2970 19867 3028 19873
rect 3237 19907 3295 19913
rect 3237 19873 3249 19907
rect 3283 19904 3295 19907
rect 3418 19904 3424 19916
rect 3283 19876 3424 19904
rect 3283 19873 3295 19876
rect 3237 19867 3295 19873
rect 198 19796 204 19848
rect 256 19836 262 19848
rect 2682 19836 2688 19848
rect 256 19808 2688 19836
rect 256 19796 262 19808
rect 2682 19796 2688 19808
rect 2740 19796 2746 19848
rect 1394 19768 1400 19780
rect 1355 19740 1400 19768
rect 1394 19728 1400 19740
rect 1452 19728 1458 19780
rect 1762 19728 1768 19780
rect 1820 19768 1826 19780
rect 2590 19768 2596 19780
rect 1820 19740 2452 19768
rect 2551 19740 2596 19768
rect 1820 19728 1826 19740
rect 2424 19700 2452 19740
rect 2590 19728 2596 19740
rect 2648 19728 2654 19780
rect 2700 19768 2728 19796
rect 2884 19768 2912 19867
rect 2976 19780 3004 19867
rect 3418 19864 3424 19876
rect 3476 19864 3482 19916
rect 3510 19864 3516 19916
rect 3568 19904 3574 19916
rect 3712 19913 3740 19944
rect 4801 19941 4813 19944
rect 4847 19941 4859 19975
rect 4801 19935 4859 19941
rect 7929 19975 7987 19981
rect 7929 19941 7941 19975
rect 7975 19972 7987 19975
rect 8662 19972 8668 19984
rect 7975 19944 8668 19972
rect 7975 19941 7987 19944
rect 7929 19935 7987 19941
rect 8662 19932 8668 19944
rect 8720 19932 8726 19984
rect 8846 19932 8852 19984
rect 8904 19972 8910 19984
rect 9306 19972 9312 19984
rect 8904 19944 9312 19972
rect 8904 19932 8910 19944
rect 9306 19932 9312 19944
rect 9364 19932 9370 19984
rect 10198 19975 10256 19981
rect 10198 19972 10210 19975
rect 9600 19944 10210 19972
rect 3697 19907 3755 19913
rect 3568 19876 3648 19904
rect 3568 19864 3574 19876
rect 3620 19836 3648 19876
rect 3697 19873 3709 19907
rect 3743 19873 3755 19907
rect 3697 19867 3755 19873
rect 3881 19907 3939 19913
rect 3881 19873 3893 19907
rect 3927 19873 3939 19907
rect 3881 19867 3939 19873
rect 4157 19907 4215 19913
rect 4157 19873 4169 19907
rect 4203 19904 4215 19907
rect 4246 19904 4252 19916
rect 4203 19876 4252 19904
rect 4203 19873 4215 19876
rect 4157 19867 4215 19873
rect 3896 19836 3924 19867
rect 4246 19864 4252 19876
rect 4304 19904 4310 19916
rect 5169 19907 5227 19913
rect 5169 19904 5181 19907
rect 4304 19876 5181 19904
rect 4304 19864 4310 19876
rect 5169 19873 5181 19876
rect 5215 19873 5227 19907
rect 8570 19904 8576 19916
rect 8531 19876 8576 19904
rect 5169 19867 5227 19873
rect 8570 19864 8576 19876
rect 8628 19864 8634 19916
rect 8754 19864 8760 19916
rect 8812 19904 8818 19916
rect 9030 19904 9036 19916
rect 8812 19876 9036 19904
rect 8812 19864 8818 19876
rect 9030 19864 9036 19876
rect 9088 19864 9094 19916
rect 9214 19864 9220 19916
rect 9272 19904 9278 19916
rect 9493 19907 9551 19913
rect 9493 19904 9505 19907
rect 9272 19876 9505 19904
rect 9272 19864 9278 19876
rect 9493 19873 9505 19876
rect 9539 19873 9551 19907
rect 9493 19867 9551 19873
rect 4985 19839 5043 19845
rect 4985 19836 4997 19839
rect 3620 19808 4997 19836
rect 4985 19805 4997 19808
rect 5031 19805 5043 19839
rect 4985 19799 5043 19805
rect 8389 19839 8447 19845
rect 8389 19805 8401 19839
rect 8435 19836 8447 19839
rect 9600 19836 9628 19944
rect 10198 19941 10210 19944
rect 10244 19972 10256 19975
rect 10594 19972 10600 19984
rect 10244 19944 10600 19972
rect 10244 19941 10256 19944
rect 10198 19935 10256 19941
rect 10594 19932 10600 19944
rect 10652 19932 10658 19984
rect 11885 19975 11943 19981
rect 11885 19941 11897 19975
rect 11931 19972 11943 19975
rect 12434 19972 12440 19984
rect 11931 19944 12440 19972
rect 11931 19941 11943 19944
rect 11885 19935 11943 19941
rect 12434 19932 12440 19944
rect 12492 19932 12498 19984
rect 12544 19972 12572 20003
rect 12710 20000 12716 20052
rect 12768 20040 12774 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 12768 20012 14105 20040
rect 12768 20000 12774 20012
rect 14093 20009 14105 20012
rect 14139 20009 14151 20043
rect 14093 20003 14151 20009
rect 14182 20000 14188 20052
rect 14240 20040 14246 20052
rect 15194 20040 15200 20052
rect 14240 20012 15200 20040
rect 14240 20000 14246 20012
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 15381 20043 15439 20049
rect 15381 20009 15393 20043
rect 15427 20040 15439 20043
rect 15838 20040 15844 20052
rect 15427 20012 15844 20040
rect 15427 20009 15439 20012
rect 15381 20003 15439 20009
rect 15838 20000 15844 20012
rect 15896 20000 15902 20052
rect 16301 20043 16359 20049
rect 16301 20009 16313 20043
rect 16347 20040 16359 20043
rect 16850 20040 16856 20052
rect 16347 20012 16856 20040
rect 16347 20009 16359 20012
rect 16301 20003 16359 20009
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 16945 20043 17003 20049
rect 16945 20009 16957 20043
rect 16991 20040 17003 20043
rect 18601 20043 18659 20049
rect 16991 20012 17816 20040
rect 16991 20009 17003 20012
rect 16945 20003 17003 20009
rect 13173 19975 13231 19981
rect 12544 19944 12940 19972
rect 9953 19907 10011 19913
rect 9953 19873 9965 19907
rect 9999 19904 10011 19907
rect 10686 19904 10692 19916
rect 9999 19876 10692 19904
rect 9999 19873 10011 19876
rect 9953 19867 10011 19873
rect 10686 19864 10692 19876
rect 10744 19864 10750 19916
rect 12345 19907 12403 19913
rect 12345 19904 12357 19907
rect 12268 19876 12357 19904
rect 8435 19808 9628 19836
rect 9677 19839 9735 19845
rect 8435 19805 8447 19808
rect 8389 19799 8447 19805
rect 9677 19805 9689 19839
rect 9723 19805 9735 19839
rect 9677 19799 9735 19805
rect 2700 19740 2912 19768
rect 2958 19728 2964 19780
rect 3016 19728 3022 19780
rect 3418 19768 3424 19780
rect 3379 19740 3424 19768
rect 3418 19728 3424 19740
rect 3476 19728 3482 19780
rect 3513 19771 3571 19777
rect 3513 19737 3525 19771
rect 3559 19768 3571 19771
rect 3786 19768 3792 19780
rect 3559 19740 3792 19768
rect 3559 19737 3571 19740
rect 3513 19731 3571 19737
rect 3786 19728 3792 19740
rect 3844 19728 3850 19780
rect 4062 19768 4068 19780
rect 4023 19740 4068 19768
rect 4062 19728 4068 19740
rect 4120 19728 4126 19780
rect 4246 19728 4252 19780
rect 4304 19768 4310 19780
rect 4433 19771 4491 19777
rect 4433 19768 4445 19771
rect 4304 19740 4445 19768
rect 4304 19728 4310 19740
rect 4433 19737 4445 19740
rect 4479 19737 4491 19771
rect 6914 19768 6920 19780
rect 4433 19731 4491 19737
rect 4816 19740 6920 19768
rect 2685 19703 2743 19709
rect 2685 19700 2697 19703
rect 2424 19672 2697 19700
rect 2685 19669 2697 19672
rect 2731 19669 2743 19703
rect 2685 19663 2743 19669
rect 2774 19660 2780 19712
rect 2832 19700 2838 19712
rect 3145 19703 3203 19709
rect 3145 19700 3157 19703
rect 2832 19672 3157 19700
rect 2832 19660 2838 19672
rect 3145 19669 3157 19672
rect 3191 19669 3203 19703
rect 3145 19663 3203 19669
rect 4341 19703 4399 19709
rect 4341 19669 4353 19703
rect 4387 19700 4399 19703
rect 4816 19700 4844 19740
rect 6914 19728 6920 19740
rect 6972 19728 6978 19780
rect 7745 19771 7803 19777
rect 7745 19737 7757 19771
rect 7791 19768 7803 19771
rect 9122 19768 9128 19780
rect 7791 19740 9128 19768
rect 7791 19737 7803 19740
rect 7745 19731 7803 19737
rect 9122 19728 9128 19740
rect 9180 19728 9186 19780
rect 9490 19728 9496 19780
rect 9548 19768 9554 19780
rect 9692 19768 9720 19799
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11609 19839 11667 19845
rect 11609 19836 11621 19839
rect 11296 19808 11621 19836
rect 11296 19796 11302 19808
rect 11609 19805 11621 19808
rect 11655 19805 11667 19839
rect 11790 19836 11796 19848
rect 11751 19808 11796 19836
rect 11609 19799 11667 19805
rect 11790 19796 11796 19808
rect 11848 19796 11854 19848
rect 12268 19777 12296 19876
rect 12345 19873 12357 19876
rect 12391 19873 12403 19907
rect 12802 19904 12808 19916
rect 12763 19876 12808 19904
rect 12345 19867 12403 19873
rect 12802 19864 12808 19876
rect 12860 19864 12866 19916
rect 12912 19913 12940 19944
rect 13173 19941 13185 19975
rect 13219 19972 13231 19975
rect 17218 19972 17224 19984
rect 13219 19944 16896 19972
rect 17179 19944 17224 19972
rect 13219 19941 13231 19944
rect 13173 19935 13231 19941
rect 12897 19907 12955 19913
rect 12897 19873 12909 19907
rect 12943 19873 12955 19907
rect 13630 19904 13636 19916
rect 13591 19876 13636 19904
rect 12897 19867 12955 19873
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 14734 19904 14740 19916
rect 14695 19876 14740 19904
rect 14734 19864 14740 19876
rect 14792 19864 14798 19916
rect 14826 19864 14832 19916
rect 14884 19904 14890 19916
rect 15197 19907 15255 19913
rect 15197 19904 15209 19907
rect 14884 19876 15209 19904
rect 14884 19864 14890 19876
rect 15197 19873 15209 19876
rect 15243 19873 15255 19907
rect 15197 19867 15255 19873
rect 15378 19864 15384 19916
rect 15436 19904 15442 19916
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 15436 19876 15485 19904
rect 15436 19864 15442 19876
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 16114 19904 16120 19916
rect 16075 19876 16120 19904
rect 15473 19867 15531 19873
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 16390 19904 16396 19916
rect 16351 19876 16396 19904
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 16482 19864 16488 19916
rect 16540 19904 16546 19916
rect 16761 19907 16819 19913
rect 16761 19904 16773 19907
rect 16540 19876 16773 19904
rect 16540 19864 16546 19876
rect 16761 19873 16773 19876
rect 16807 19873 16819 19907
rect 16868 19904 16896 19944
rect 17218 19932 17224 19944
rect 17276 19932 17282 19984
rect 17586 19972 17592 19984
rect 17547 19944 17592 19972
rect 17586 19932 17592 19944
rect 17644 19932 17650 19984
rect 17788 19981 17816 20012
rect 18601 20009 18613 20043
rect 18647 20009 18659 20043
rect 18601 20003 18659 20009
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 18782 20040 18788 20052
rect 18739 20012 18788 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 17773 19975 17831 19981
rect 17773 19941 17785 19975
rect 17819 19941 17831 19975
rect 18046 19972 18052 19984
rect 18007 19944 18052 19972
rect 17773 19935 17831 19941
rect 18046 19932 18052 19944
rect 18104 19932 18110 19984
rect 18616 19972 18644 20003
rect 18782 20000 18788 20012
rect 18840 20000 18846 20052
rect 19150 20040 19156 20052
rect 19111 20012 19156 20040
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 19426 20040 19432 20052
rect 19387 20012 19432 20040
rect 19426 20000 19432 20012
rect 19484 20000 19490 20052
rect 19889 20043 19947 20049
rect 19889 20009 19901 20043
rect 19935 20040 19947 20043
rect 20438 20040 20444 20052
rect 19935 20012 20444 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 20438 20000 20444 20012
rect 20496 20000 20502 20052
rect 21177 20043 21235 20049
rect 21177 20009 21189 20043
rect 21223 20009 21235 20043
rect 21177 20003 21235 20009
rect 18616 19944 18736 19972
rect 17405 19907 17463 19913
rect 17405 19904 17417 19907
rect 16868 19876 17417 19904
rect 16761 19867 16819 19873
rect 17405 19873 17417 19876
rect 17451 19873 17463 19907
rect 17405 19867 17463 19873
rect 17954 19864 17960 19916
rect 18012 19904 18018 19916
rect 18233 19907 18291 19913
rect 18233 19904 18245 19907
rect 18012 19876 18245 19904
rect 18012 19864 18018 19876
rect 18233 19873 18245 19876
rect 18279 19873 18291 19907
rect 18233 19867 18291 19873
rect 18417 19907 18475 19913
rect 18417 19873 18429 19907
rect 18463 19873 18475 19907
rect 18417 19867 18475 19873
rect 13354 19836 13360 19848
rect 12544 19808 13360 19836
rect 9548 19740 9720 19768
rect 12253 19771 12311 19777
rect 9548 19728 9554 19740
rect 12253 19737 12265 19771
rect 12299 19737 12311 19771
rect 12253 19731 12311 19737
rect 4387 19672 4844 19700
rect 4387 19669 4399 19672
rect 4341 19663 4399 19669
rect 4890 19660 4896 19712
rect 4948 19700 4954 19712
rect 5353 19703 5411 19709
rect 5353 19700 5365 19703
rect 4948 19672 5365 19700
rect 4948 19660 4954 19672
rect 5353 19669 5365 19672
rect 5399 19669 5411 19703
rect 5353 19663 5411 19669
rect 6270 19660 6276 19712
rect 6328 19700 6334 19712
rect 8846 19700 8852 19712
rect 6328 19672 8852 19700
rect 6328 19660 6334 19672
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 8941 19703 8999 19709
rect 8941 19669 8953 19703
rect 8987 19700 8999 19703
rect 9950 19700 9956 19712
rect 8987 19672 9956 19700
rect 8987 19669 8999 19672
rect 8941 19663 8999 19669
rect 9950 19660 9956 19672
rect 10008 19660 10014 19712
rect 11333 19703 11391 19709
rect 11333 19669 11345 19703
rect 11379 19700 11391 19703
rect 12544 19700 12572 19808
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13538 19796 13544 19848
rect 13596 19836 13602 19848
rect 14461 19839 14519 19845
rect 13596 19808 13641 19836
rect 13596 19796 13602 19808
rect 14461 19805 14473 19839
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19836 14703 19839
rect 14691 19808 15148 19836
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 13372 19768 13400 19796
rect 14476 19768 14504 19799
rect 13372 19740 14504 19768
rect 14550 19728 14556 19780
rect 14608 19768 14614 19780
rect 14826 19768 14832 19780
rect 14608 19740 14832 19768
rect 14608 19728 14614 19740
rect 14826 19728 14832 19740
rect 14884 19728 14890 19780
rect 15120 19768 15148 19808
rect 15562 19796 15568 19848
rect 15620 19836 15626 19848
rect 16025 19839 16083 19845
rect 16025 19836 16037 19839
rect 15620 19808 16037 19836
rect 15620 19796 15626 19808
rect 16025 19805 16037 19808
rect 16071 19836 16083 19839
rect 17126 19836 17132 19848
rect 16071 19808 17132 19836
rect 16071 19805 16083 19808
rect 16025 19799 16083 19805
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 15580 19768 15608 19796
rect 15120 19740 15608 19768
rect 15657 19771 15715 19777
rect 15657 19737 15669 19771
rect 15703 19768 15715 19771
rect 16666 19768 16672 19780
rect 15703 19740 16672 19768
rect 15703 19737 15715 19740
rect 15657 19731 15715 19737
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 18046 19768 18052 19780
rect 16960 19740 18052 19768
rect 11379 19672 12572 19700
rect 12621 19703 12679 19709
rect 11379 19669 11391 19672
rect 11333 19663 11391 19669
rect 12621 19669 12633 19703
rect 12667 19700 12679 19703
rect 12986 19700 12992 19712
rect 12667 19672 12992 19700
rect 12667 19669 12679 19672
rect 12621 19663 12679 19669
rect 12986 19660 12992 19672
rect 13044 19660 13050 19712
rect 13081 19703 13139 19709
rect 13081 19669 13093 19703
rect 13127 19700 13139 19703
rect 13173 19703 13231 19709
rect 13173 19700 13185 19703
rect 13127 19672 13185 19700
rect 13127 19669 13139 19672
rect 13081 19663 13139 19669
rect 13173 19669 13185 19672
rect 13219 19669 13231 19703
rect 13998 19700 14004 19712
rect 13959 19672 14004 19700
rect 13173 19663 13231 19669
rect 13998 19660 14004 19672
rect 14056 19660 14062 19712
rect 14090 19660 14096 19712
rect 14148 19700 14154 19712
rect 14918 19700 14924 19712
rect 14148 19672 14924 19700
rect 14148 19660 14154 19672
rect 14918 19660 14924 19672
rect 14976 19660 14982 19712
rect 15102 19700 15108 19712
rect 15063 19672 15108 19700
rect 15102 19660 15108 19672
rect 15160 19660 15166 19712
rect 15286 19660 15292 19712
rect 15344 19700 15350 19712
rect 15749 19703 15807 19709
rect 15749 19700 15761 19703
rect 15344 19672 15761 19700
rect 15344 19660 15350 19672
rect 15749 19669 15761 19672
rect 15795 19669 15807 19703
rect 15749 19663 15807 19669
rect 16577 19703 16635 19709
rect 16577 19669 16589 19703
rect 16623 19700 16635 19703
rect 16960 19700 16988 19740
rect 18046 19728 18052 19740
rect 18104 19728 18110 19780
rect 18432 19768 18460 19867
rect 18708 19836 18736 19944
rect 19058 19932 19064 19984
rect 19116 19972 19122 19984
rect 20622 19972 20628 19984
rect 19116 19944 20484 19972
rect 20583 19944 20628 19972
rect 19116 19932 19122 19944
rect 18874 19904 18880 19916
rect 18835 19876 18880 19904
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 18969 19907 19027 19913
rect 18969 19873 18981 19907
rect 19015 19904 19027 19907
rect 19150 19904 19156 19916
rect 19015 19876 19156 19904
rect 19015 19873 19027 19876
rect 18969 19867 19027 19873
rect 19150 19864 19156 19876
rect 19208 19864 19214 19916
rect 19242 19864 19248 19916
rect 19300 19904 19306 19916
rect 19300 19876 19345 19904
rect 19300 19864 19306 19876
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 19705 19907 19763 19913
rect 19705 19904 19717 19907
rect 19668 19876 19717 19904
rect 19668 19864 19674 19876
rect 19705 19873 19717 19876
rect 19751 19873 19763 19907
rect 19978 19904 19984 19916
rect 19939 19876 19984 19904
rect 19705 19867 19763 19873
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 20346 19904 20352 19916
rect 20307 19876 20352 19904
rect 20346 19864 20352 19876
rect 20404 19864 20410 19916
rect 20456 19904 20484 19944
rect 20622 19932 20628 19944
rect 20680 19932 20686 19984
rect 20898 19972 20904 19984
rect 20732 19944 20904 19972
rect 20732 19904 20760 19944
rect 20898 19932 20904 19944
rect 20956 19932 20962 19984
rect 21192 19972 21220 20003
rect 21361 19975 21419 19981
rect 21361 19972 21373 19975
rect 21192 19944 21373 19972
rect 21361 19941 21373 19944
rect 21407 19941 21419 19975
rect 21361 19935 21419 19941
rect 20456 19876 20760 19904
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 20993 19907 21051 19913
rect 20864 19876 20909 19904
rect 20864 19864 20870 19876
rect 20993 19873 21005 19907
rect 21039 19904 21051 19907
rect 21082 19904 21088 19916
rect 21039 19876 21088 19904
rect 21039 19873 21051 19876
rect 20993 19867 21051 19873
rect 21082 19864 21088 19876
rect 21140 19864 21146 19916
rect 20898 19836 20904 19848
rect 18708 19808 20904 19836
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 20165 19771 20223 19777
rect 18432 19740 20116 19768
rect 17126 19700 17132 19712
rect 16623 19672 16988 19700
rect 17087 19672 17132 19700
rect 16623 19669 16635 19672
rect 16577 19663 16635 19669
rect 17126 19660 17132 19672
rect 17184 19660 17190 19712
rect 17678 19660 17684 19712
rect 17736 19700 17742 19712
rect 18782 19700 18788 19712
rect 17736 19672 18788 19700
rect 17736 19660 17742 19672
rect 18782 19660 18788 19672
rect 18840 19660 18846 19712
rect 18874 19660 18880 19712
rect 18932 19700 18938 19712
rect 19518 19700 19524 19712
rect 18932 19672 19524 19700
rect 18932 19660 18938 19672
rect 19518 19660 19524 19672
rect 19576 19660 19582 19712
rect 20088 19700 20116 19740
rect 20165 19737 20177 19771
rect 20211 19768 20223 19771
rect 20990 19768 20996 19780
rect 20211 19740 20996 19768
rect 20211 19737 20223 19740
rect 20165 19731 20223 19737
rect 20990 19728 20996 19740
rect 21048 19728 21054 19780
rect 21542 19768 21548 19780
rect 21503 19740 21548 19768
rect 21542 19728 21548 19740
rect 21600 19728 21606 19780
rect 20254 19700 20260 19712
rect 20088 19672 20260 19700
rect 20254 19660 20260 19672
rect 20312 19660 20318 19712
rect 20441 19703 20499 19709
rect 20441 19669 20453 19703
rect 20487 19700 20499 19703
rect 21910 19700 21916 19712
rect 20487 19672 21916 19700
rect 20487 19669 20499 19672
rect 20441 19663 20499 19669
rect 21910 19660 21916 19672
rect 21968 19660 21974 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1946 19456 1952 19508
rect 2004 19496 2010 19508
rect 2317 19499 2375 19505
rect 2317 19496 2329 19499
rect 2004 19468 2329 19496
rect 2004 19456 2010 19468
rect 2317 19465 2329 19468
rect 2363 19465 2375 19499
rect 2317 19459 2375 19465
rect 2777 19499 2835 19505
rect 2777 19465 2789 19499
rect 2823 19496 2835 19499
rect 3050 19496 3056 19508
rect 2823 19468 3056 19496
rect 2823 19465 2835 19468
rect 2777 19459 2835 19465
rect 3050 19456 3056 19468
rect 3108 19456 3114 19508
rect 3234 19456 3240 19508
rect 3292 19496 3298 19508
rect 3329 19499 3387 19505
rect 3329 19496 3341 19499
rect 3292 19468 3341 19496
rect 3292 19456 3298 19468
rect 3329 19465 3341 19468
rect 3375 19465 3387 19499
rect 3329 19459 3387 19465
rect 3418 19456 3424 19508
rect 3476 19496 3482 19508
rect 5442 19496 5448 19508
rect 3476 19468 5448 19496
rect 3476 19456 3482 19468
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 7745 19499 7803 19505
rect 7745 19465 7757 19499
rect 7791 19496 7803 19499
rect 9490 19496 9496 19508
rect 7791 19468 9496 19496
rect 7791 19465 7803 19468
rect 7745 19459 7803 19465
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 10594 19496 10600 19508
rect 10555 19468 10600 19496
rect 10594 19456 10600 19468
rect 10652 19456 10658 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19496 11575 19499
rect 11698 19496 11704 19508
rect 11563 19468 11704 19496
rect 11563 19465 11575 19468
rect 11517 19459 11575 19465
rect 11698 19456 11704 19468
rect 11756 19456 11762 19508
rect 12894 19456 12900 19508
rect 12952 19496 12958 19508
rect 15286 19496 15292 19508
rect 12952 19468 15292 19496
rect 12952 19456 12958 19468
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 15470 19456 15476 19508
rect 15528 19496 15534 19508
rect 15749 19499 15807 19505
rect 15749 19496 15761 19499
rect 15528 19468 15761 19496
rect 15528 19456 15534 19468
rect 15749 19465 15761 19468
rect 15795 19465 15807 19499
rect 15749 19459 15807 19465
rect 17126 19456 17132 19508
rect 17184 19496 17190 19508
rect 18782 19496 18788 19508
rect 17184 19468 18460 19496
rect 18743 19468 18788 19496
rect 17184 19456 17190 19468
rect 1578 19388 1584 19440
rect 1636 19428 1642 19440
rect 2041 19431 2099 19437
rect 2041 19428 2053 19431
rect 1636 19400 2053 19428
rect 1636 19388 1642 19400
rect 2041 19397 2053 19400
rect 2087 19397 2099 19431
rect 2041 19391 2099 19397
rect 2682 19388 2688 19440
rect 2740 19428 2746 19440
rect 3145 19431 3203 19437
rect 3145 19428 3157 19431
rect 2740 19400 3157 19428
rect 2740 19388 2746 19400
rect 3145 19397 3157 19400
rect 3191 19397 3203 19431
rect 3145 19391 3203 19397
rect 4062 19388 4068 19440
rect 4120 19428 4126 19440
rect 8110 19428 8116 19440
rect 4120 19400 8116 19428
rect 4120 19388 4126 19400
rect 8110 19388 8116 19400
rect 8168 19388 8174 19440
rect 11333 19431 11391 19437
rect 11333 19397 11345 19431
rect 11379 19428 11391 19431
rect 12066 19428 12072 19440
rect 11379 19400 12072 19428
rect 11379 19397 11391 19400
rect 11333 19391 11391 19397
rect 12066 19388 12072 19400
rect 12124 19388 12130 19440
rect 14553 19431 14611 19437
rect 14553 19397 14565 19431
rect 14599 19428 14611 19431
rect 14642 19428 14648 19440
rect 14599 19400 14648 19428
rect 14599 19397 14611 19400
rect 14553 19391 14611 19397
rect 14642 19388 14648 19400
rect 14700 19428 14706 19440
rect 14700 19400 14780 19428
rect 14700 19388 14706 19400
rect 2130 19320 2136 19372
rect 2188 19360 2194 19372
rect 3234 19360 3240 19372
rect 2188 19332 3240 19360
rect 2188 19320 2194 19332
rect 3234 19320 3240 19332
rect 3292 19320 3298 19372
rect 3694 19320 3700 19372
rect 3752 19360 3758 19372
rect 7742 19360 7748 19372
rect 3752 19332 7748 19360
rect 3752 19320 3758 19332
rect 7742 19320 7748 19332
rect 7800 19320 7806 19372
rect 11238 19360 11244 19372
rect 10704 19332 11244 19360
rect 1394 19292 1400 19304
rect 1355 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19252 1458 19304
rect 1762 19292 1768 19304
rect 1723 19264 1768 19292
rect 1762 19252 1768 19264
rect 1820 19252 1826 19304
rect 2225 19295 2283 19301
rect 2225 19261 2237 19295
rect 2271 19261 2283 19295
rect 2225 19255 2283 19261
rect 1581 19227 1639 19233
rect 1581 19193 1593 19227
rect 1627 19224 1639 19227
rect 2038 19224 2044 19236
rect 1627 19196 2044 19224
rect 1627 19193 1639 19196
rect 1581 19187 1639 19193
rect 2038 19184 2044 19196
rect 2096 19184 2102 19236
rect 2240 19224 2268 19255
rect 2406 19252 2412 19304
rect 2464 19292 2470 19304
rect 2501 19295 2559 19301
rect 2501 19292 2513 19295
rect 2464 19264 2513 19292
rect 2464 19252 2470 19264
rect 2501 19261 2513 19264
rect 2547 19261 2559 19295
rect 2501 19255 2559 19261
rect 2593 19295 2651 19301
rect 2593 19261 2605 19295
rect 2639 19292 2651 19295
rect 2682 19292 2688 19304
rect 2639 19264 2688 19292
rect 2639 19261 2651 19264
rect 2593 19255 2651 19261
rect 2682 19252 2688 19264
rect 2740 19252 2746 19304
rect 2869 19295 2927 19301
rect 2869 19261 2881 19295
rect 2915 19292 2927 19295
rect 3050 19292 3056 19304
rect 2915 19264 3056 19292
rect 2915 19261 2927 19264
rect 2869 19255 2927 19261
rect 3050 19252 3056 19264
rect 3108 19252 3114 19304
rect 3510 19292 3516 19304
rect 3471 19264 3516 19292
rect 3510 19252 3516 19264
rect 3568 19252 3574 19304
rect 3602 19252 3608 19304
rect 3660 19292 3666 19304
rect 3970 19292 3976 19304
rect 3660 19264 3705 19292
rect 3931 19264 3976 19292
rect 3660 19252 3666 19264
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 6273 19295 6331 19301
rect 4632 19264 6224 19292
rect 4632 19224 4660 19264
rect 2240 19196 2544 19224
rect 1946 19156 1952 19168
rect 1907 19128 1952 19156
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 2516 19156 2544 19196
rect 3068 19196 4660 19224
rect 4709 19227 4767 19233
rect 2958 19156 2964 19168
rect 2516 19128 2964 19156
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3068 19165 3096 19196
rect 4709 19193 4721 19227
rect 4755 19224 4767 19227
rect 5902 19224 5908 19236
rect 4755 19196 5908 19224
rect 4755 19193 4767 19196
rect 4709 19187 4767 19193
rect 5902 19184 5908 19196
rect 5960 19184 5966 19236
rect 6196 19224 6224 19264
rect 6273 19261 6285 19295
rect 6319 19292 6331 19295
rect 6454 19292 6460 19304
rect 6319 19264 6460 19292
rect 6319 19261 6331 19264
rect 6273 19255 6331 19261
rect 6454 19252 6460 19264
rect 6512 19252 6518 19304
rect 9122 19292 9128 19304
rect 9083 19264 9128 19292
rect 9122 19252 9128 19264
rect 9180 19292 9186 19304
rect 9217 19295 9275 19301
rect 9217 19292 9229 19295
rect 9180 19264 9229 19292
rect 9180 19252 9186 19264
rect 9217 19261 9229 19264
rect 9263 19261 9275 19295
rect 10704 19292 10732 19332
rect 11238 19320 11244 19332
rect 11296 19360 11302 19372
rect 11698 19360 11704 19372
rect 11296 19332 11704 19360
rect 11296 19320 11302 19332
rect 11698 19320 11704 19332
rect 11756 19320 11762 19372
rect 14752 19369 14780 19400
rect 14918 19388 14924 19440
rect 14976 19388 14982 19440
rect 15381 19431 15439 19437
rect 15381 19397 15393 19431
rect 15427 19428 15439 19431
rect 16114 19428 16120 19440
rect 15427 19400 16120 19428
rect 15427 19397 15439 19400
rect 15381 19391 15439 19397
rect 16114 19388 16120 19400
rect 16172 19388 16178 19440
rect 16945 19431 17003 19437
rect 16945 19397 16957 19431
rect 16991 19397 17003 19431
rect 16945 19391 17003 19397
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19329 14795 19363
rect 14936 19360 14964 19388
rect 16960 19360 16988 19391
rect 18138 19388 18144 19440
rect 18196 19428 18202 19440
rect 18325 19431 18383 19437
rect 18325 19428 18337 19431
rect 18196 19400 18337 19428
rect 18196 19388 18202 19400
rect 18325 19397 18337 19400
rect 18371 19397 18383 19431
rect 18432 19428 18460 19468
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 19610 19496 19616 19508
rect 19352 19468 19616 19496
rect 19352 19428 19380 19468
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 18432 19400 19380 19428
rect 18325 19391 18383 19397
rect 19426 19388 19432 19440
rect 19484 19428 19490 19440
rect 20346 19428 20352 19440
rect 19484 19400 20352 19428
rect 19484 19388 19490 19400
rect 20346 19388 20352 19400
rect 20404 19388 20410 19440
rect 14936 19332 16988 19360
rect 17405 19363 17463 19369
rect 14737 19323 14795 19329
rect 17405 19329 17417 19363
rect 17451 19360 17463 19363
rect 18230 19360 18236 19372
rect 17451 19332 18236 19360
rect 17451 19329 17463 19332
rect 17405 19323 17463 19329
rect 18230 19320 18236 19332
rect 18288 19320 18294 19372
rect 18598 19320 18604 19372
rect 18656 19360 18662 19372
rect 19242 19360 19248 19372
rect 18656 19332 19248 19360
rect 18656 19320 18662 19332
rect 19242 19320 19248 19332
rect 19300 19320 19306 19372
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19360 19763 19363
rect 19794 19360 19800 19372
rect 19751 19332 19800 19360
rect 19751 19329 19763 19332
rect 19705 19323 19763 19329
rect 19794 19320 19800 19332
rect 19852 19360 19858 19372
rect 20441 19363 20499 19369
rect 20441 19360 20453 19363
rect 19852 19332 20453 19360
rect 19852 19320 19858 19332
rect 20441 19329 20453 19332
rect 20487 19329 20499 19363
rect 20441 19323 20499 19329
rect 9217 19255 9275 19261
rect 9416 19264 10732 19292
rect 8880 19227 8938 19233
rect 6196 19196 7880 19224
rect 3053 19159 3111 19165
rect 3053 19125 3065 19159
rect 3099 19125 3111 19159
rect 3053 19119 3111 19125
rect 3694 19116 3700 19168
rect 3752 19156 3758 19168
rect 3789 19159 3847 19165
rect 3789 19156 3801 19159
rect 3752 19128 3801 19156
rect 3752 19116 3758 19128
rect 3789 19125 3801 19128
rect 3835 19125 3847 19159
rect 3789 19119 3847 19125
rect 3970 19116 3976 19168
rect 4028 19156 4034 19168
rect 4985 19159 5043 19165
rect 4985 19156 4997 19159
rect 4028 19128 4997 19156
rect 4028 19116 4034 19128
rect 4985 19125 4997 19128
rect 5031 19125 5043 19159
rect 6086 19156 6092 19168
rect 6047 19128 6092 19156
rect 4985 19119 5043 19125
rect 6086 19116 6092 19128
rect 6144 19116 6150 19168
rect 7852 19156 7880 19196
rect 8880 19193 8892 19227
rect 8926 19224 8938 19227
rect 9416 19224 9444 19264
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 13446 19301 13452 19304
rect 11057 19295 11115 19301
rect 11057 19292 11069 19295
rect 10836 19264 11069 19292
rect 10836 19252 10842 19264
rect 11057 19261 11069 19264
rect 11103 19261 11115 19295
rect 11057 19255 11115 19261
rect 13081 19295 13139 19301
rect 13081 19261 13093 19295
rect 13127 19292 13139 19295
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 13127 19264 13185 19292
rect 13127 19261 13139 19264
rect 13081 19255 13139 19261
rect 13173 19261 13185 19264
rect 13219 19261 13231 19295
rect 13440 19292 13452 19301
rect 13407 19264 13452 19292
rect 13173 19255 13231 19261
rect 13440 19255 13452 19264
rect 9490 19233 9496 19236
rect 8926 19196 9444 19224
rect 8926 19193 8938 19196
rect 8880 19187 8938 19193
rect 9484 19187 9496 19233
rect 9548 19224 9554 19236
rect 9548 19196 9584 19224
rect 10520 19196 12434 19224
rect 9490 19184 9496 19187
rect 9548 19184 9554 19196
rect 10520 19156 10548 19196
rect 7852 19128 10548 19156
rect 10686 19116 10692 19168
rect 10744 19156 10750 19168
rect 11698 19156 11704 19168
rect 10744 19128 10789 19156
rect 11659 19128 11704 19156
rect 10744 19116 10750 19128
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 12406 19156 12434 19196
rect 12802 19184 12808 19236
rect 12860 19233 12866 19236
rect 12860 19224 12872 19233
rect 13096 19224 13124 19255
rect 13446 19252 13452 19255
rect 13504 19252 13510 19304
rect 13906 19292 13912 19304
rect 13556 19264 13912 19292
rect 13556 19224 13584 19264
rect 13906 19252 13912 19264
rect 13964 19252 13970 19304
rect 14182 19252 14188 19304
rect 14240 19292 14246 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14240 19264 14933 19292
rect 14240 19252 14246 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19292 15071 19295
rect 15102 19292 15108 19304
rect 15059 19264 15108 19292
rect 15059 19261 15071 19264
rect 15013 19255 15071 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15212 19264 15945 19292
rect 12860 19196 12905 19224
rect 13096 19196 13584 19224
rect 12860 19187 12872 19196
rect 12860 19184 12866 19187
rect 13814 19184 13820 19236
rect 13872 19224 13878 19236
rect 14826 19224 14832 19236
rect 13872 19196 14832 19224
rect 13872 19184 13878 19196
rect 14826 19184 14832 19196
rect 14884 19184 14890 19236
rect 13722 19156 13728 19168
rect 12406 19128 13728 19156
rect 13722 19116 13728 19128
rect 13780 19116 13786 19168
rect 13906 19116 13912 19168
rect 13964 19156 13970 19168
rect 15212 19156 15240 19264
rect 15933 19261 15945 19264
rect 15979 19261 15991 19295
rect 16298 19292 16304 19304
rect 16259 19264 16304 19292
rect 15933 19255 15991 19261
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 16577 19295 16635 19301
rect 16577 19261 16589 19295
rect 16623 19292 16635 19295
rect 16666 19292 16672 19304
rect 16623 19264 16672 19292
rect 16623 19261 16635 19264
rect 16577 19255 16635 19261
rect 16666 19252 16672 19264
rect 16724 19252 16730 19304
rect 17126 19292 17132 19304
rect 17087 19264 17132 19292
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 18046 19292 18052 19304
rect 18007 19264 18052 19292
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 18517 19295 18575 19301
rect 18517 19292 18529 19295
rect 18196 19264 18529 19292
rect 18196 19252 18202 19264
rect 18517 19261 18529 19264
rect 18563 19261 18575 19295
rect 18966 19292 18972 19304
rect 18927 19264 18972 19292
rect 18517 19255 18575 19261
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 19058 19252 19064 19304
rect 19116 19292 19122 19304
rect 19521 19295 19579 19301
rect 19521 19292 19533 19295
rect 19116 19264 19533 19292
rect 19116 19252 19122 19264
rect 19521 19261 19533 19264
rect 19567 19261 19579 19295
rect 19521 19255 19579 19261
rect 19978 19252 19984 19304
rect 20036 19252 20042 19304
rect 20898 19252 20904 19304
rect 20956 19292 20962 19304
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20956 19264 21005 19292
rect 20956 19252 20962 19264
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 21082 19252 21088 19304
rect 21140 19252 21146 19304
rect 21542 19292 21548 19304
rect 21503 19264 21548 19292
rect 21542 19252 21548 19264
rect 21600 19252 21606 19304
rect 15286 19184 15292 19236
rect 15344 19224 15350 19236
rect 17589 19227 17647 19233
rect 15344 19196 16436 19224
rect 15344 19184 15350 19196
rect 15654 19156 15660 19168
rect 13964 19128 15240 19156
rect 15615 19128 15660 19156
rect 13964 19116 13970 19128
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 16022 19116 16028 19168
rect 16080 19156 16086 19168
rect 16408 19165 16436 19196
rect 17589 19193 17601 19227
rect 17635 19224 17647 19227
rect 17770 19224 17776 19236
rect 17635 19196 17776 19224
rect 17635 19193 17647 19196
rect 17589 19187 17647 19193
rect 17770 19184 17776 19196
rect 17828 19184 17834 19236
rect 19996 19224 20024 19252
rect 18616 19196 20024 19224
rect 20349 19227 20407 19233
rect 16117 19159 16175 19165
rect 16117 19156 16129 19159
rect 16080 19128 16129 19156
rect 16080 19116 16086 19128
rect 16117 19125 16129 19128
rect 16163 19125 16175 19159
rect 16117 19119 16175 19125
rect 16393 19159 16451 19165
rect 16393 19125 16405 19159
rect 16439 19125 16451 19159
rect 16666 19156 16672 19168
rect 16627 19128 16672 19156
rect 16393 19119 16451 19125
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 17494 19156 17500 19168
rect 17455 19128 17500 19156
rect 17494 19116 17500 19128
rect 17552 19116 17558 19168
rect 17678 19116 17684 19168
rect 17736 19156 17742 19168
rect 17957 19159 18015 19165
rect 17957 19156 17969 19159
rect 17736 19128 17969 19156
rect 17736 19116 17742 19128
rect 17957 19125 17969 19128
rect 18003 19125 18015 19159
rect 17957 19119 18015 19125
rect 18233 19159 18291 19165
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18322 19156 18328 19168
rect 18279 19128 18328 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18322 19116 18328 19128
rect 18380 19116 18386 19168
rect 18414 19116 18420 19168
rect 18472 19156 18478 19168
rect 18616 19165 18644 19196
rect 20349 19193 20361 19227
rect 20395 19224 20407 19227
rect 21100 19224 21128 19252
rect 20395 19196 21128 19224
rect 20395 19193 20407 19196
rect 20349 19187 20407 19193
rect 21266 19184 21272 19236
rect 21324 19224 21330 19236
rect 21361 19227 21419 19233
rect 21361 19224 21373 19227
rect 21324 19196 21373 19224
rect 21324 19184 21330 19196
rect 21361 19193 21373 19196
rect 21407 19193 21419 19227
rect 21361 19187 21419 19193
rect 18601 19159 18659 19165
rect 18601 19156 18613 19159
rect 18472 19128 18613 19156
rect 18472 19116 18478 19128
rect 18601 19125 18613 19128
rect 18647 19125 18659 19159
rect 18601 19119 18659 19125
rect 18874 19116 18880 19168
rect 18932 19156 18938 19168
rect 19061 19159 19119 19165
rect 19061 19156 19073 19159
rect 18932 19128 19073 19156
rect 18932 19116 18938 19128
rect 19061 19125 19073 19128
rect 19107 19125 19119 19159
rect 19061 19119 19119 19125
rect 19429 19159 19487 19165
rect 19429 19125 19441 19159
rect 19475 19156 19487 19159
rect 19610 19156 19616 19168
rect 19475 19128 19616 19156
rect 19475 19125 19487 19128
rect 19429 19119 19487 19125
rect 19610 19116 19616 19128
rect 19668 19116 19674 19168
rect 19886 19156 19892 19168
rect 19847 19128 19892 19156
rect 19886 19116 19892 19128
rect 19944 19116 19950 19168
rect 19978 19116 19984 19168
rect 20036 19156 20042 19168
rect 20257 19159 20315 19165
rect 20257 19156 20269 19159
rect 20036 19128 20269 19156
rect 20036 19116 20042 19128
rect 20257 19125 20269 19128
rect 20303 19125 20315 19159
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 20257 19119 20315 19125
rect 20714 19116 20720 19128
rect 20772 19156 20778 19168
rect 20990 19156 20996 19168
rect 20772 19128 20996 19156
rect 20772 19116 20778 19128
rect 20990 19116 20996 19128
rect 21048 19116 21054 19168
rect 21085 19159 21143 19165
rect 21085 19125 21097 19159
rect 21131 19156 21143 19159
rect 22278 19156 22284 19168
rect 21131 19128 22284 19156
rect 21131 19125 21143 19128
rect 21085 19119 21143 19125
rect 22278 19116 22284 19128
rect 22336 19116 22342 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 1949 18955 2007 18961
rect 1949 18921 1961 18955
rect 1995 18921 2007 18955
rect 2498 18952 2504 18964
rect 2459 18924 2504 18952
rect 1949 18915 2007 18921
rect 1964 18884 1992 18915
rect 2498 18912 2504 18924
rect 2556 18912 2562 18964
rect 2777 18955 2835 18961
rect 2777 18921 2789 18955
rect 2823 18952 2835 18955
rect 2866 18952 2872 18964
rect 2823 18924 2872 18952
rect 2823 18921 2835 18924
rect 2777 18915 2835 18921
rect 2866 18912 2872 18924
rect 2924 18912 2930 18964
rect 3142 18912 3148 18964
rect 3200 18952 3206 18964
rect 3421 18955 3479 18961
rect 3421 18952 3433 18955
rect 3200 18924 3433 18952
rect 3200 18912 3206 18924
rect 3421 18921 3433 18924
rect 3467 18952 3479 18955
rect 3602 18952 3608 18964
rect 3467 18924 3608 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 3602 18912 3608 18924
rect 3660 18912 3666 18964
rect 3878 18912 3884 18964
rect 3936 18952 3942 18964
rect 6086 18952 6092 18964
rect 3936 18924 6092 18952
rect 3936 18912 3942 18924
rect 6086 18912 6092 18924
rect 6144 18912 6150 18964
rect 6454 18952 6460 18964
rect 6415 18924 6460 18952
rect 6454 18912 6460 18924
rect 6512 18912 6518 18964
rect 8570 18912 8576 18964
rect 8628 18952 8634 18964
rect 9125 18955 9183 18961
rect 9125 18952 9137 18955
rect 8628 18924 9137 18952
rect 8628 18912 8634 18924
rect 9125 18921 9137 18924
rect 9171 18921 9183 18955
rect 9125 18915 9183 18921
rect 9493 18955 9551 18961
rect 9493 18921 9505 18955
rect 9539 18952 9551 18955
rect 10686 18952 10692 18964
rect 9539 18924 10692 18952
rect 9539 18921 9551 18924
rect 9493 18915 9551 18921
rect 10686 18912 10692 18924
rect 10744 18912 10750 18964
rect 11790 18912 11796 18964
rect 11848 18952 11854 18964
rect 12161 18955 12219 18961
rect 12161 18952 12173 18955
rect 11848 18924 12173 18952
rect 11848 18912 11854 18924
rect 12161 18921 12173 18924
rect 12207 18921 12219 18955
rect 12161 18915 12219 18921
rect 12434 18912 12440 18964
rect 12492 18952 12498 18964
rect 12989 18955 13047 18961
rect 12989 18952 13001 18955
rect 12492 18924 13001 18952
rect 12492 18912 12498 18924
rect 12989 18921 13001 18924
rect 13035 18921 13047 18955
rect 12989 18915 13047 18921
rect 14093 18955 14151 18961
rect 14093 18921 14105 18955
rect 14139 18952 14151 18955
rect 14734 18952 14740 18964
rect 14139 18924 14740 18952
rect 14139 18921 14151 18924
rect 14093 18915 14151 18921
rect 14734 18912 14740 18924
rect 14792 18912 14798 18964
rect 15930 18912 15936 18964
rect 15988 18912 15994 18964
rect 17497 18955 17555 18961
rect 17497 18921 17509 18955
rect 17543 18952 17555 18955
rect 17586 18952 17592 18964
rect 17543 18924 17592 18952
rect 17543 18921 17555 18924
rect 17497 18915 17555 18921
rect 17586 18912 17592 18924
rect 17644 18912 17650 18964
rect 17773 18955 17831 18961
rect 17773 18921 17785 18955
rect 17819 18952 17831 18955
rect 18138 18952 18144 18964
rect 17819 18924 18144 18952
rect 17819 18921 17831 18924
rect 17773 18915 17831 18921
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 3326 18884 3332 18896
rect 1964 18856 3332 18884
rect 3326 18844 3332 18856
rect 3384 18844 3390 18896
rect 3694 18844 3700 18896
rect 3752 18884 3758 18896
rect 5718 18884 5724 18896
rect 3752 18856 5724 18884
rect 3752 18844 3758 18856
rect 5718 18844 5724 18856
rect 5776 18844 5782 18896
rect 5902 18844 5908 18896
rect 5960 18884 5966 18896
rect 8846 18884 8852 18896
rect 5960 18856 8852 18884
rect 5960 18844 5966 18856
rect 8846 18844 8852 18856
rect 8904 18844 8910 18896
rect 9582 18844 9588 18896
rect 9640 18884 9646 18896
rect 10229 18887 10287 18893
rect 10229 18884 10241 18887
rect 9640 18856 10241 18884
rect 9640 18844 9646 18856
rect 10229 18853 10241 18856
rect 10275 18853 10287 18887
rect 10229 18847 10287 18853
rect 10956 18887 11014 18893
rect 10956 18853 10968 18887
rect 11002 18884 11014 18887
rect 11054 18884 11060 18896
rect 11002 18856 11060 18884
rect 11002 18853 11014 18856
rect 10956 18847 11014 18853
rect 11054 18844 11060 18856
rect 11112 18844 11118 18896
rect 14366 18884 14372 18896
rect 11164 18856 14372 18884
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 1578 18816 1584 18828
rect 1539 18788 1584 18816
rect 1578 18776 1584 18788
rect 1636 18776 1642 18828
rect 1762 18816 1768 18828
rect 1723 18788 1768 18816
rect 1762 18776 1768 18788
rect 1820 18776 1826 18828
rect 2041 18819 2099 18825
rect 2041 18785 2053 18819
rect 2087 18816 2099 18819
rect 2130 18816 2136 18828
rect 2087 18788 2136 18816
rect 2087 18785 2099 18788
rect 2041 18779 2099 18785
rect 2130 18776 2136 18788
rect 2188 18776 2194 18828
rect 2314 18816 2320 18828
rect 2275 18788 2320 18816
rect 2314 18776 2320 18788
rect 2372 18776 2378 18828
rect 2593 18819 2651 18825
rect 2593 18785 2605 18819
rect 2639 18785 2651 18819
rect 2593 18779 2651 18785
rect 1670 18708 1676 18760
rect 1728 18748 1734 18760
rect 2608 18748 2636 18779
rect 5350 18776 5356 18828
rect 5408 18816 5414 18828
rect 5997 18819 6055 18825
rect 5997 18816 6009 18819
rect 5408 18788 6009 18816
rect 5408 18776 5414 18788
rect 5997 18785 6009 18788
rect 6043 18785 6055 18819
rect 5997 18779 6055 18785
rect 6641 18819 6699 18825
rect 6641 18785 6653 18819
rect 6687 18816 6699 18819
rect 7006 18816 7012 18828
rect 6687 18788 7012 18816
rect 6687 18785 6699 18788
rect 6641 18779 6699 18785
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 8294 18776 8300 18828
rect 8352 18816 8358 18828
rect 8573 18819 8631 18825
rect 8573 18816 8585 18819
rect 8352 18788 8585 18816
rect 8352 18776 8358 18788
rect 8573 18785 8585 18788
rect 8619 18785 8631 18819
rect 9214 18816 9220 18828
rect 8573 18779 8631 18785
rect 8680 18788 9220 18816
rect 1728 18720 2636 18748
rect 1728 18708 1734 18720
rect 2682 18708 2688 18760
rect 2740 18748 2746 18760
rect 3326 18748 3332 18760
rect 2740 18720 3332 18748
rect 2740 18708 2746 18720
rect 3326 18708 3332 18720
rect 3384 18708 3390 18760
rect 3510 18708 3516 18760
rect 3568 18748 3574 18760
rect 3697 18751 3755 18757
rect 3697 18748 3709 18751
rect 3568 18720 3709 18748
rect 3568 18708 3574 18720
rect 3697 18717 3709 18720
rect 3743 18748 3755 18751
rect 8680 18748 8708 18788
rect 9214 18776 9220 18788
rect 9272 18776 9278 18828
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 9950 18816 9956 18828
rect 9548 18788 9720 18816
rect 9911 18788 9956 18816
rect 9548 18776 9554 18788
rect 3743 18720 8708 18748
rect 8941 18751 8999 18757
rect 3743 18717 3755 18720
rect 3697 18711 3755 18717
rect 8941 18717 8953 18751
rect 8987 18748 8999 18751
rect 9582 18748 9588 18760
rect 8987 18720 9588 18748
rect 8987 18717 8999 18720
rect 8941 18711 8999 18717
rect 9582 18708 9588 18720
rect 9640 18708 9646 18760
rect 9692 18757 9720 18788
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 11164 18816 11192 18856
rect 14366 18844 14372 18856
rect 14424 18844 14430 18896
rect 14642 18893 14648 18896
rect 14636 18884 14648 18893
rect 14603 18856 14648 18884
rect 14636 18847 14648 18856
rect 14642 18844 14648 18847
rect 14700 18844 14706 18896
rect 15948 18884 15976 18912
rect 14752 18856 15976 18884
rect 10060 18788 11192 18816
rect 9677 18751 9735 18757
rect 9677 18717 9689 18751
rect 9723 18717 9735 18751
rect 9677 18711 9735 18717
rect 2222 18680 2228 18692
rect 2183 18652 2228 18680
rect 2222 18640 2228 18652
rect 2280 18640 2286 18692
rect 2958 18640 2964 18692
rect 3016 18680 3022 18692
rect 8386 18680 8392 18692
rect 3016 18652 8392 18680
rect 3016 18640 3022 18652
rect 8386 18640 8392 18652
rect 8444 18640 8450 18692
rect 8757 18683 8815 18689
rect 8757 18649 8769 18683
rect 8803 18680 8815 18683
rect 10060 18680 10088 18788
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 12529 18819 12587 18825
rect 12529 18816 12541 18819
rect 12492 18788 12541 18816
rect 12492 18776 12498 18788
rect 12529 18785 12541 18788
rect 12575 18785 12587 18819
rect 12529 18779 12587 18785
rect 12621 18819 12679 18825
rect 12621 18785 12633 18819
rect 12667 18816 12679 18819
rect 12894 18816 12900 18828
rect 12667 18788 12900 18816
rect 12667 18785 12679 18788
rect 12621 18779 12679 18785
rect 12894 18776 12900 18788
rect 12952 18776 12958 18828
rect 13170 18776 13176 18828
rect 13228 18816 13234 18828
rect 13357 18819 13415 18825
rect 13357 18816 13369 18819
rect 13228 18788 13369 18816
rect 13228 18776 13234 18788
rect 13357 18785 13369 18788
rect 13403 18785 13415 18819
rect 13357 18779 13415 18785
rect 13449 18819 13507 18825
rect 13449 18785 13461 18819
rect 13495 18816 13507 18819
rect 13495 18788 13676 18816
rect 13495 18785 13507 18788
rect 13449 18779 13507 18785
rect 10686 18748 10692 18760
rect 10647 18720 10692 18748
rect 10686 18708 10692 18720
rect 10744 18708 10750 18760
rect 11790 18708 11796 18760
rect 11848 18748 11854 18760
rect 12250 18748 12256 18760
rect 11848 18720 12256 18748
rect 11848 18708 11854 18720
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 12802 18708 12808 18760
rect 12860 18748 12866 18760
rect 13541 18751 13599 18757
rect 12860 18720 12953 18748
rect 12860 18708 12866 18720
rect 13541 18717 13553 18751
rect 13587 18717 13599 18751
rect 13648 18748 13676 18788
rect 13722 18776 13728 18828
rect 13780 18816 13786 18828
rect 14752 18816 14780 18856
rect 16666 18844 16672 18896
rect 16724 18884 16730 18896
rect 18506 18884 18512 18896
rect 16724 18856 18512 18884
rect 16724 18844 16730 18856
rect 18506 18844 18512 18856
rect 18564 18844 18570 18896
rect 18874 18844 18880 18896
rect 18932 18884 18938 18896
rect 19426 18884 19432 18896
rect 18932 18856 19432 18884
rect 18932 18844 18938 18856
rect 19426 18844 19432 18856
rect 19484 18844 19490 18896
rect 19610 18844 19616 18896
rect 19668 18884 19674 18896
rect 19794 18884 19800 18896
rect 19668 18856 19800 18884
rect 19668 18844 19674 18856
rect 19794 18844 19800 18856
rect 19852 18893 19858 18896
rect 19852 18887 19916 18893
rect 19852 18853 19870 18887
rect 19904 18853 19916 18887
rect 19852 18847 19916 18853
rect 19852 18844 19858 18847
rect 13780 18788 14780 18816
rect 13780 18776 13786 18788
rect 15930 18776 15936 18828
rect 15988 18816 15994 18828
rect 16097 18819 16155 18825
rect 16097 18816 16109 18819
rect 15988 18788 16109 18816
rect 15988 18776 15994 18788
rect 16097 18785 16109 18788
rect 16143 18785 16155 18819
rect 16097 18779 16155 18785
rect 16850 18776 16856 18828
rect 16908 18816 16914 18828
rect 17313 18819 17371 18825
rect 17313 18816 17325 18819
rect 16908 18788 17325 18816
rect 16908 18776 16914 18788
rect 17313 18785 17325 18788
rect 17359 18785 17371 18819
rect 17313 18779 17371 18785
rect 17589 18819 17647 18825
rect 17589 18785 17601 18819
rect 17635 18816 17647 18819
rect 17678 18816 17684 18828
rect 17635 18788 17684 18816
rect 17635 18785 17647 18788
rect 17589 18779 17647 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 18230 18825 18236 18828
rect 18224 18816 18236 18825
rect 18191 18788 18236 18816
rect 18224 18779 18236 18788
rect 18230 18776 18236 18779
rect 18288 18776 18294 18828
rect 18782 18776 18788 18828
rect 18840 18816 18846 18828
rect 20806 18816 20812 18828
rect 18840 18788 20812 18816
rect 18840 18776 18846 18788
rect 20806 18776 20812 18788
rect 20864 18776 20870 18828
rect 21358 18816 21364 18828
rect 21319 18788 21364 18816
rect 21358 18776 21364 18788
rect 21416 18776 21422 18828
rect 21542 18816 21548 18828
rect 21503 18788 21548 18816
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 14182 18748 14188 18760
rect 13648 18720 14188 18748
rect 13541 18711 13599 18717
rect 8803 18652 10088 18680
rect 10137 18683 10195 18689
rect 8803 18649 8815 18652
rect 8757 18643 8815 18649
rect 10137 18649 10149 18683
rect 10183 18680 10195 18683
rect 12069 18683 12127 18689
rect 10183 18652 10732 18680
rect 10183 18649 10195 18652
rect 10137 18643 10195 18649
rect 2406 18572 2412 18624
rect 2464 18612 2470 18624
rect 3053 18615 3111 18621
rect 3053 18612 3065 18615
rect 2464 18584 3065 18612
rect 2464 18572 2470 18584
rect 3053 18581 3065 18584
rect 3099 18612 3111 18615
rect 3142 18612 3148 18624
rect 3099 18584 3148 18612
rect 3099 18581 3111 18584
rect 3053 18575 3111 18581
rect 3142 18572 3148 18584
rect 3200 18572 3206 18624
rect 3326 18612 3332 18624
rect 3239 18584 3332 18612
rect 3326 18572 3332 18584
rect 3384 18612 3390 18624
rect 4062 18612 4068 18624
rect 3384 18584 4068 18612
rect 3384 18572 3390 18584
rect 4062 18572 4068 18584
rect 4120 18572 4126 18624
rect 6181 18615 6239 18621
rect 6181 18581 6193 18615
rect 6227 18612 6239 18615
rect 8662 18612 8668 18624
rect 6227 18584 8668 18612
rect 6227 18581 6239 18584
rect 6181 18575 6239 18581
rect 8662 18572 8668 18584
rect 8720 18572 8726 18624
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 9490 18612 9496 18624
rect 9272 18584 9496 18612
rect 9272 18572 9278 18584
rect 9490 18572 9496 18584
rect 9548 18612 9554 18624
rect 10413 18615 10471 18621
rect 10413 18612 10425 18615
rect 9548 18584 10425 18612
rect 9548 18572 9554 18584
rect 10413 18581 10425 18584
rect 10459 18581 10471 18615
rect 10704 18612 10732 18652
rect 12069 18649 12081 18683
rect 12115 18680 12127 18683
rect 12820 18680 12848 18708
rect 13556 18680 13584 18711
rect 14182 18708 14188 18720
rect 14240 18708 14246 18760
rect 14366 18748 14372 18760
rect 14327 18720 14372 18748
rect 14366 18708 14372 18720
rect 14424 18708 14430 18760
rect 15838 18748 15844 18760
rect 15799 18720 15844 18748
rect 15838 18708 15844 18720
rect 15896 18708 15902 18760
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 17957 18751 18015 18757
rect 17957 18748 17969 18751
rect 17000 18720 17969 18748
rect 17000 18708 17006 18720
rect 17957 18717 17969 18720
rect 18003 18717 18015 18751
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 17957 18711 18015 18717
rect 18984 18720 19625 18748
rect 12115 18652 13584 18680
rect 15304 18652 15884 18680
rect 12115 18649 12127 18652
rect 12069 18643 12127 18649
rect 15304 18612 15332 18652
rect 15746 18612 15752 18624
rect 10704 18584 15332 18612
rect 15707 18584 15752 18612
rect 10413 18575 10471 18581
rect 15746 18572 15752 18584
rect 15804 18572 15810 18624
rect 15856 18612 15884 18652
rect 16574 18612 16580 18624
rect 15856 18584 16580 18612
rect 16574 18572 16580 18584
rect 16632 18572 16638 18624
rect 17221 18615 17279 18621
rect 17221 18581 17233 18615
rect 17267 18612 17279 18615
rect 17310 18612 17316 18624
rect 17267 18584 17316 18612
rect 17267 18581 17279 18584
rect 17221 18575 17279 18581
rect 17310 18572 17316 18584
rect 17368 18572 17374 18624
rect 17972 18612 18000 18711
rect 18984 18612 19012 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 17972 18584 19012 18612
rect 19337 18615 19395 18621
rect 19337 18581 19349 18615
rect 19383 18612 19395 18615
rect 19610 18612 19616 18624
rect 19383 18584 19616 18612
rect 19383 18581 19395 18584
rect 19337 18575 19395 18581
rect 19610 18572 19616 18584
rect 19668 18572 19674 18624
rect 19794 18572 19800 18624
rect 19852 18612 19858 18624
rect 20993 18615 21051 18621
rect 20993 18612 21005 18615
rect 19852 18584 21005 18612
rect 19852 18572 19858 18584
rect 20993 18581 21005 18584
rect 21039 18581 21051 18615
rect 20993 18575 21051 18581
rect 21082 18572 21088 18624
rect 21140 18612 21146 18624
rect 21140 18584 21185 18612
rect 21140 18572 21146 18584
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 1486 18408 1492 18420
rect 1447 18380 1492 18408
rect 1486 18368 1492 18380
rect 1544 18368 1550 18420
rect 1578 18368 1584 18420
rect 1636 18408 1642 18420
rect 2133 18411 2191 18417
rect 2133 18408 2145 18411
rect 1636 18380 2145 18408
rect 1636 18368 1642 18380
rect 2133 18377 2145 18380
rect 2179 18377 2191 18411
rect 2133 18371 2191 18377
rect 3142 18368 3148 18420
rect 3200 18368 3206 18420
rect 5350 18408 5356 18420
rect 5311 18380 5356 18408
rect 5350 18368 5356 18380
rect 5408 18368 5414 18420
rect 7650 18368 7656 18420
rect 7708 18408 7714 18420
rect 8294 18408 8300 18420
rect 7708 18380 8217 18408
rect 8255 18380 8300 18408
rect 7708 18368 7714 18380
rect 2038 18300 2044 18352
rect 2096 18340 2102 18352
rect 2409 18343 2467 18349
rect 2409 18340 2421 18343
rect 2096 18312 2421 18340
rect 2096 18300 2102 18312
rect 2409 18309 2421 18312
rect 2455 18309 2467 18343
rect 3160 18340 3188 18368
rect 5626 18340 5632 18352
rect 3160 18312 5632 18340
rect 2409 18303 2467 18309
rect 5626 18300 5632 18312
rect 5684 18300 5690 18352
rect 8189 18340 8217 18380
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 8386 18368 8392 18420
rect 8444 18408 8450 18420
rect 12250 18408 12256 18420
rect 8444 18380 12256 18408
rect 8444 18368 8450 18380
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 12437 18411 12495 18417
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 12483 18380 12664 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 12526 18340 12532 18352
rect 8189 18312 12532 18340
rect 12526 18300 12532 18312
rect 12584 18300 12590 18352
rect 12636 18340 12664 18380
rect 12710 18368 12716 18420
rect 12768 18408 12774 18420
rect 12897 18411 12955 18417
rect 12897 18408 12909 18411
rect 12768 18380 12909 18408
rect 12768 18368 12774 18380
rect 12897 18377 12909 18380
rect 12943 18377 12955 18411
rect 12897 18371 12955 18377
rect 15838 18368 15844 18420
rect 15896 18408 15902 18420
rect 16942 18408 16948 18420
rect 15896 18380 16948 18408
rect 15896 18368 15902 18380
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 18138 18368 18144 18420
rect 18196 18408 18202 18420
rect 18325 18411 18383 18417
rect 18325 18408 18337 18411
rect 18196 18380 18337 18408
rect 18196 18368 18202 18380
rect 18325 18377 18337 18380
rect 18371 18377 18383 18411
rect 18325 18371 18383 18377
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 20073 18411 20131 18417
rect 20073 18408 20085 18411
rect 19392 18380 20085 18408
rect 19392 18368 19398 18380
rect 20073 18377 20085 18380
rect 20119 18377 20131 18411
rect 20073 18371 20131 18377
rect 20533 18411 20591 18417
rect 20533 18377 20545 18411
rect 20579 18408 20591 18411
rect 21358 18408 21364 18420
rect 20579 18380 21364 18408
rect 20579 18377 20591 18380
rect 20533 18371 20591 18377
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 13814 18340 13820 18352
rect 12636 18312 13820 18340
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 14182 18340 14188 18352
rect 13924 18312 14188 18340
rect 1762 18232 1768 18284
rect 1820 18232 1826 18284
rect 2332 18244 2820 18272
rect 1780 18204 1808 18232
rect 2332 18213 2360 18244
rect 2317 18207 2375 18213
rect 1780 18176 2268 18204
rect 1578 18136 1584 18148
rect 1539 18108 1584 18136
rect 1578 18096 1584 18108
rect 1636 18096 1642 18148
rect 1946 18136 1952 18148
rect 1907 18108 1952 18136
rect 1946 18096 1952 18108
rect 2004 18096 2010 18148
rect 2240 18136 2268 18176
rect 2317 18173 2329 18207
rect 2363 18173 2375 18207
rect 2590 18204 2596 18216
rect 2551 18176 2596 18204
rect 2317 18167 2375 18173
rect 2590 18164 2596 18176
rect 2648 18164 2654 18216
rect 2792 18213 2820 18244
rect 7558 18232 7564 18284
rect 7616 18272 7622 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7616 18244 7849 18272
rect 7616 18232 7622 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 7926 18232 7932 18284
rect 7984 18272 7990 18284
rect 10229 18275 10287 18281
rect 10229 18272 10241 18275
rect 7984 18244 10241 18272
rect 7984 18232 7990 18244
rect 10229 18241 10241 18244
rect 10275 18241 10287 18275
rect 10410 18272 10416 18284
rect 10371 18244 10416 18272
rect 10229 18235 10287 18241
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 10594 18272 10600 18284
rect 10555 18244 10600 18272
rect 10594 18232 10600 18244
rect 10652 18232 10658 18284
rect 10778 18232 10784 18284
rect 10836 18272 10842 18284
rect 11149 18275 11207 18281
rect 11149 18272 11161 18275
rect 10836 18244 11161 18272
rect 10836 18232 10842 18244
rect 11149 18241 11161 18244
rect 11195 18241 11207 18275
rect 11149 18235 11207 18241
rect 11606 18232 11612 18284
rect 11664 18272 11670 18284
rect 11793 18275 11851 18281
rect 11793 18272 11805 18275
rect 11664 18244 11805 18272
rect 11664 18232 11670 18244
rect 11793 18241 11805 18244
rect 11839 18241 11851 18275
rect 11793 18235 11851 18241
rect 12713 18275 12771 18281
rect 12713 18241 12725 18275
rect 12759 18272 12771 18275
rect 13078 18272 13084 18284
rect 12759 18244 13084 18272
rect 12759 18241 12771 18244
rect 12713 18235 12771 18241
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18272 13231 18275
rect 13924 18272 13952 18312
rect 14182 18300 14188 18312
rect 14240 18300 14246 18352
rect 18046 18300 18052 18352
rect 18104 18340 18110 18352
rect 18782 18340 18788 18352
rect 18104 18312 18788 18340
rect 18104 18300 18110 18312
rect 18782 18300 18788 18312
rect 18840 18300 18846 18352
rect 19794 18340 19800 18352
rect 19076 18312 19800 18340
rect 13219 18244 13952 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 13998 18232 14004 18284
rect 14056 18272 14062 18284
rect 14366 18272 14372 18284
rect 14056 18244 14372 18272
rect 14056 18232 14062 18244
rect 14366 18232 14372 18244
rect 14424 18272 14430 18284
rect 14553 18275 14611 18281
rect 14553 18272 14565 18275
rect 14424 18244 14565 18272
rect 14424 18232 14430 18244
rect 14553 18241 14565 18244
rect 14599 18241 14611 18275
rect 15746 18272 15752 18284
rect 14553 18235 14611 18241
rect 15580 18244 15752 18272
rect 2777 18207 2835 18213
rect 2777 18173 2789 18207
rect 2823 18204 2835 18207
rect 3142 18204 3148 18216
rect 2823 18176 3148 18204
rect 2823 18173 2835 18176
rect 2777 18167 2835 18173
rect 3142 18164 3148 18176
rect 3200 18164 3206 18216
rect 5166 18204 5172 18216
rect 5127 18176 5172 18204
rect 5166 18164 5172 18176
rect 5224 18164 5230 18216
rect 7282 18204 7288 18216
rect 5920 18176 7288 18204
rect 2961 18139 3019 18145
rect 2961 18136 2973 18139
rect 2240 18108 2973 18136
rect 2961 18105 2973 18108
rect 3007 18136 3019 18139
rect 4982 18136 4988 18148
rect 3007 18108 4988 18136
rect 3007 18105 3019 18108
rect 2961 18099 3019 18105
rect 4982 18096 4988 18108
rect 5040 18096 5046 18148
rect 1854 18068 1860 18080
rect 1815 18040 1860 18068
rect 1854 18028 1860 18040
rect 1912 18028 1918 18080
rect 3145 18071 3203 18077
rect 3145 18037 3157 18071
rect 3191 18068 3203 18071
rect 3234 18068 3240 18080
rect 3191 18040 3240 18068
rect 3191 18037 3203 18040
rect 3145 18031 3203 18037
rect 3234 18028 3240 18040
rect 3292 18068 3298 18080
rect 5920 18068 5948 18176
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 7466 18164 7472 18216
rect 7524 18204 7530 18216
rect 8113 18207 8171 18213
rect 8113 18204 8125 18207
rect 7524 18176 8125 18204
rect 7524 18164 7530 18176
rect 8113 18173 8125 18176
rect 8159 18173 8171 18207
rect 8113 18167 8171 18173
rect 8662 18164 8668 18216
rect 8720 18204 8726 18216
rect 14274 18204 14280 18216
rect 8720 18176 14280 18204
rect 8720 18164 8726 18176
rect 14274 18164 14280 18176
rect 14332 18164 14338 18216
rect 14820 18207 14878 18213
rect 14820 18204 14832 18207
rect 14752 18176 14832 18204
rect 14752 18148 14780 18176
rect 14820 18173 14832 18176
rect 14866 18204 14878 18207
rect 15580 18204 15608 18244
rect 15746 18232 15752 18244
rect 15804 18272 15810 18284
rect 16577 18275 16635 18281
rect 16577 18272 16589 18275
rect 15804 18244 16589 18272
rect 15804 18232 15810 18244
rect 16577 18241 16589 18244
rect 16623 18241 16635 18275
rect 16577 18235 16635 18241
rect 16942 18232 16948 18284
rect 17000 18281 17006 18284
rect 19076 18281 19104 18312
rect 19794 18300 19800 18312
rect 19852 18300 19858 18352
rect 20346 18340 20352 18352
rect 19904 18312 20352 18340
rect 17000 18272 17010 18281
rect 19061 18275 19119 18281
rect 17000 18244 17045 18272
rect 17000 18235 17010 18244
rect 19061 18241 19073 18275
rect 19107 18241 19119 18275
rect 19242 18272 19248 18284
rect 19203 18244 19248 18272
rect 19061 18235 19119 18241
rect 17000 18232 17006 18235
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 19904 18272 19932 18312
rect 20346 18300 20352 18312
rect 20404 18300 20410 18352
rect 21542 18340 21548 18352
rect 21503 18312 21548 18340
rect 21542 18300 21548 18312
rect 21600 18300 21606 18352
rect 19352 18244 19932 18272
rect 14866 18176 15608 18204
rect 14866 18173 14878 18176
rect 14820 18167 14878 18173
rect 15654 18164 15660 18216
rect 15712 18204 15718 18216
rect 16393 18207 16451 18213
rect 16393 18204 16405 18207
rect 15712 18176 16405 18204
rect 15712 18164 15718 18176
rect 16393 18173 16405 18176
rect 16439 18173 16451 18207
rect 18874 18204 18880 18216
rect 16393 18167 16451 18173
rect 16500 18176 18880 18204
rect 7650 18096 7656 18148
rect 7708 18136 7714 18148
rect 7708 18108 7753 18136
rect 7708 18096 7714 18108
rect 8846 18096 8852 18148
rect 8904 18136 8910 18148
rect 9950 18136 9956 18148
rect 8904 18108 9956 18136
rect 8904 18096 8910 18108
rect 9950 18096 9956 18108
rect 10008 18096 10014 18148
rect 11977 18139 12035 18145
rect 11977 18136 11989 18139
rect 11256 18108 11989 18136
rect 7282 18068 7288 18080
rect 3292 18040 5948 18068
rect 7243 18040 7288 18068
rect 3292 18028 3298 18040
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 7745 18071 7803 18077
rect 7745 18037 7757 18071
rect 7791 18068 7803 18071
rect 8294 18068 8300 18080
rect 7791 18040 8300 18068
rect 7791 18037 7803 18040
rect 7745 18031 7803 18037
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 8386 18028 8392 18080
rect 8444 18068 8450 18080
rect 10134 18068 10140 18080
rect 8444 18040 10140 18068
rect 8444 18028 8450 18040
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10229 18071 10287 18077
rect 10229 18037 10241 18071
rect 10275 18068 10287 18071
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 10275 18040 10701 18068
rect 10275 18037 10287 18040
rect 10229 18031 10287 18037
rect 10689 18037 10701 18040
rect 10735 18068 10747 18071
rect 10778 18068 10784 18080
rect 10735 18040 10784 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11057 18071 11115 18077
rect 11057 18037 11069 18071
rect 11103 18068 11115 18071
rect 11256 18068 11284 18108
rect 11977 18105 11989 18108
rect 12023 18105 12035 18139
rect 11977 18099 12035 18105
rect 13814 18096 13820 18148
rect 13872 18136 13878 18148
rect 14093 18139 14151 18145
rect 14093 18136 14105 18139
rect 13872 18108 14105 18136
rect 13872 18096 13878 18108
rect 14093 18105 14105 18108
rect 14139 18105 14151 18139
rect 14093 18099 14151 18105
rect 14182 18096 14188 18148
rect 14240 18136 14246 18148
rect 14642 18136 14648 18148
rect 14240 18108 14648 18136
rect 14240 18096 14246 18108
rect 14642 18096 14648 18108
rect 14700 18096 14706 18148
rect 14734 18096 14740 18148
rect 14792 18096 14798 18148
rect 16500 18136 16528 18176
rect 18874 18164 18880 18176
rect 18932 18164 18938 18216
rect 19352 18204 19380 18244
rect 19886 18204 19892 18216
rect 18984 18176 19380 18204
rect 19444 18176 19892 18204
rect 14844 18108 16528 18136
rect 17212 18139 17270 18145
rect 12066 18068 12072 18080
rect 11103 18040 11284 18068
rect 12027 18040 12072 18068
rect 11103 18037 11115 18040
rect 11057 18031 11115 18037
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 13354 18068 13360 18080
rect 12492 18040 13360 18068
rect 12492 18028 12498 18040
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 13446 18028 13452 18080
rect 13504 18068 13510 18080
rect 14844 18068 14872 18108
rect 17212 18105 17224 18139
rect 17258 18136 17270 18139
rect 17310 18136 17316 18148
rect 17258 18108 17316 18136
rect 17258 18105 17270 18108
rect 17212 18099 17270 18105
rect 17310 18096 17316 18108
rect 17368 18096 17374 18148
rect 18785 18139 18843 18145
rect 18785 18136 18797 18139
rect 17420 18108 18797 18136
rect 13504 18040 14872 18068
rect 13504 18028 13510 18040
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 15933 18071 15991 18077
rect 15933 18068 15945 18071
rect 15896 18040 15945 18068
rect 15896 18028 15902 18040
rect 15933 18037 15945 18040
rect 15979 18037 15991 18071
rect 15933 18031 15991 18037
rect 16025 18071 16083 18077
rect 16025 18037 16037 18071
rect 16071 18068 16083 18071
rect 16114 18068 16120 18080
rect 16071 18040 16120 18068
rect 16071 18037 16083 18040
rect 16025 18031 16083 18037
rect 16114 18028 16120 18040
rect 16172 18028 16178 18080
rect 16482 18068 16488 18080
rect 16443 18040 16488 18068
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 17420 18068 17448 18108
rect 18785 18105 18797 18108
rect 18831 18136 18843 18139
rect 18984 18136 19012 18176
rect 19444 18136 19472 18176
rect 19886 18164 19892 18176
rect 19944 18164 19950 18216
rect 19978 18164 19984 18216
rect 20036 18204 20042 18216
rect 20257 18207 20315 18213
rect 20036 18176 20081 18204
rect 20036 18164 20042 18176
rect 20257 18173 20269 18207
rect 20303 18173 20315 18207
rect 20257 18167 20315 18173
rect 20272 18136 20300 18167
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 20622 18204 20628 18216
rect 20404 18176 20449 18204
rect 20583 18176 20628 18204
rect 20404 18164 20410 18176
rect 20622 18164 20628 18176
rect 20680 18164 20686 18216
rect 18831 18108 19012 18136
rect 19352 18108 19472 18136
rect 19996 18108 20300 18136
rect 18831 18105 18843 18108
rect 18785 18099 18843 18105
rect 16632 18040 17448 18068
rect 16632 18028 16638 18040
rect 18414 18028 18420 18080
rect 18472 18068 18478 18080
rect 19352 18077 19380 18108
rect 19996 18080 20024 18108
rect 20438 18096 20444 18148
rect 20496 18136 20502 18148
rect 20993 18139 21051 18145
rect 20993 18136 21005 18139
rect 20496 18108 21005 18136
rect 20496 18096 20502 18108
rect 20993 18105 21005 18108
rect 21039 18105 21051 18139
rect 21174 18136 21180 18148
rect 21135 18108 21180 18136
rect 20993 18099 21051 18105
rect 21174 18096 21180 18108
rect 21232 18096 21238 18148
rect 21361 18139 21419 18145
rect 21361 18105 21373 18139
rect 21407 18105 21419 18139
rect 21361 18099 21419 18105
rect 19337 18071 19395 18077
rect 18472 18040 18517 18068
rect 18472 18028 18478 18040
rect 19337 18037 19349 18071
rect 19383 18037 19395 18071
rect 19337 18031 19395 18037
rect 19426 18028 19432 18080
rect 19484 18068 19490 18080
rect 19705 18071 19763 18077
rect 19705 18068 19717 18071
rect 19484 18040 19717 18068
rect 19484 18028 19490 18040
rect 19705 18037 19717 18040
rect 19751 18037 19763 18071
rect 19705 18031 19763 18037
rect 19978 18028 19984 18080
rect 20036 18028 20042 18080
rect 20809 18071 20867 18077
rect 20809 18037 20821 18071
rect 20855 18068 20867 18071
rect 21376 18068 21404 18099
rect 20855 18040 21404 18068
rect 20855 18037 20867 18040
rect 20809 18031 20867 18037
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 2317 17867 2375 17873
rect 2317 17833 2329 17867
rect 2363 17864 2375 17867
rect 2590 17864 2596 17876
rect 2363 17836 2596 17864
rect 2363 17833 2375 17836
rect 2317 17827 2375 17833
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 6454 17864 6460 17876
rect 2746 17836 6460 17864
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17728 1639 17731
rect 1854 17728 1860 17740
rect 1627 17700 1860 17728
rect 1627 17697 1639 17700
rect 1581 17691 1639 17697
rect 1854 17688 1860 17700
rect 1912 17688 1918 17740
rect 2133 17731 2191 17737
rect 2133 17697 2145 17731
rect 2179 17728 2191 17731
rect 2746 17728 2774 17836
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 7009 17867 7067 17873
rect 7009 17833 7021 17867
rect 7055 17864 7067 17867
rect 7282 17864 7288 17876
rect 7055 17836 7288 17864
rect 7055 17833 7067 17836
rect 7009 17827 7067 17833
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 7466 17864 7472 17876
rect 7427 17836 7472 17864
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 7742 17824 7748 17876
rect 7800 17864 7806 17876
rect 8021 17867 8079 17873
rect 8021 17864 8033 17867
rect 7800 17836 8033 17864
rect 7800 17824 7806 17836
rect 8021 17833 8033 17836
rect 8067 17864 8079 17867
rect 8389 17867 8447 17873
rect 8389 17864 8401 17867
rect 8067 17836 8401 17864
rect 8067 17833 8079 17836
rect 8021 17827 8079 17833
rect 8389 17833 8401 17836
rect 8435 17864 8447 17867
rect 10962 17864 10968 17876
rect 8435 17836 10968 17864
rect 8435 17833 8447 17836
rect 8389 17827 8447 17833
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 11149 17867 11207 17873
rect 11149 17864 11161 17867
rect 11112 17836 11161 17864
rect 11112 17824 11118 17836
rect 11149 17833 11161 17836
rect 11195 17864 11207 17867
rect 11606 17864 11612 17876
rect 11195 17836 11612 17864
rect 11195 17833 11207 17836
rect 11149 17827 11207 17833
rect 11606 17824 11612 17836
rect 11664 17824 11670 17876
rect 11977 17867 12035 17873
rect 11977 17833 11989 17867
rect 12023 17864 12035 17867
rect 12066 17864 12072 17876
rect 12023 17836 12072 17864
rect 12023 17833 12035 17836
rect 11977 17827 12035 17833
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 14550 17824 14556 17876
rect 14608 17864 14614 17876
rect 14645 17867 14703 17873
rect 14645 17864 14657 17867
rect 14608 17836 14657 17864
rect 14608 17824 14614 17836
rect 14645 17833 14657 17836
rect 14691 17833 14703 17867
rect 14645 17827 14703 17833
rect 15473 17867 15531 17873
rect 15473 17833 15485 17867
rect 15519 17864 15531 17867
rect 15841 17867 15899 17873
rect 15841 17864 15853 17867
rect 15519 17836 15853 17864
rect 15519 17833 15531 17836
rect 15473 17827 15531 17833
rect 15841 17833 15853 17836
rect 15887 17833 15899 17867
rect 15841 17827 15899 17833
rect 15933 17867 15991 17873
rect 15933 17833 15945 17867
rect 15979 17864 15991 17867
rect 16114 17864 16120 17876
rect 15979 17836 16120 17864
rect 15979 17833 15991 17836
rect 15933 17827 15991 17833
rect 16114 17824 16120 17836
rect 16172 17824 16178 17876
rect 16301 17867 16359 17873
rect 16301 17833 16313 17867
rect 16347 17864 16359 17867
rect 16390 17864 16396 17876
rect 16347 17836 16396 17864
rect 16347 17833 16359 17836
rect 16301 17827 16359 17833
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 17494 17824 17500 17876
rect 17552 17864 17558 17876
rect 17681 17867 17739 17873
rect 17681 17864 17693 17867
rect 17552 17836 17693 17864
rect 17552 17824 17558 17836
rect 17681 17833 17693 17836
rect 17727 17833 17739 17867
rect 17681 17827 17739 17833
rect 17770 17824 17776 17876
rect 17828 17864 17834 17876
rect 18141 17867 18199 17873
rect 17828 17836 17873 17864
rect 17828 17824 17834 17836
rect 18141 17833 18153 17867
rect 18187 17864 18199 17867
rect 18414 17864 18420 17876
rect 18187 17836 18420 17864
rect 18187 17833 18199 17836
rect 18141 17827 18199 17833
rect 18414 17824 18420 17836
rect 18472 17824 18478 17876
rect 18966 17824 18972 17876
rect 19024 17864 19030 17876
rect 19245 17867 19303 17873
rect 19245 17864 19257 17867
rect 19024 17836 19257 17864
rect 19024 17824 19030 17836
rect 19245 17833 19257 17836
rect 19291 17833 19303 17867
rect 19245 17827 19303 17833
rect 5350 17756 5356 17808
rect 5408 17805 5414 17808
rect 5408 17799 5472 17805
rect 5408 17765 5426 17799
rect 5460 17765 5472 17799
rect 5408 17759 5472 17765
rect 5408 17756 5414 17759
rect 5534 17756 5540 17808
rect 5592 17796 5598 17808
rect 5592 17768 6868 17796
rect 5592 17756 5598 17768
rect 2179 17700 2774 17728
rect 5169 17731 5227 17737
rect 2179 17697 2191 17700
rect 2133 17691 2191 17697
rect 5169 17697 5181 17731
rect 5215 17728 5227 17731
rect 6178 17728 6184 17740
rect 5215 17700 6184 17728
rect 5215 17697 5227 17700
rect 5169 17691 5227 17697
rect 6178 17688 6184 17700
rect 6236 17688 6242 17740
rect 6840 17728 6868 17768
rect 6914 17756 6920 17808
rect 6972 17796 6978 17808
rect 12894 17796 12900 17808
rect 6972 17768 7788 17796
rect 6972 17756 6978 17768
rect 7760 17740 7788 17768
rect 9646 17768 12900 17796
rect 6840 17700 7052 17728
rect 6914 17660 6920 17672
rect 6875 17632 6920 17660
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 7024 17660 7052 17700
rect 7098 17688 7104 17740
rect 7156 17728 7162 17740
rect 7156 17700 7201 17728
rect 7156 17688 7162 17700
rect 7742 17688 7748 17740
rect 7800 17688 7806 17740
rect 7929 17731 7987 17737
rect 7929 17697 7941 17731
rect 7975 17728 7987 17731
rect 9646 17728 9674 17768
rect 12894 17756 12900 17768
rect 12952 17756 12958 17808
rect 15013 17799 15071 17805
rect 15013 17796 15025 17799
rect 13004 17768 15025 17796
rect 7975 17700 9674 17728
rect 10036 17731 10094 17737
rect 7975 17697 7987 17700
rect 7929 17691 7987 17697
rect 10036 17697 10048 17731
rect 10082 17728 10094 17731
rect 10410 17728 10416 17740
rect 10082 17700 10416 17728
rect 10082 17697 10094 17700
rect 10036 17691 10094 17697
rect 7944 17660 7972 17691
rect 10410 17688 10416 17700
rect 10468 17728 10474 17740
rect 11609 17731 11667 17737
rect 10468 17700 11192 17728
rect 10468 17688 10474 17700
rect 7024 17632 7972 17660
rect 8113 17663 8171 17669
rect 8113 17629 8125 17663
rect 8159 17629 8171 17663
rect 8113 17623 8171 17629
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 4062 17592 4068 17604
rect 3568 17564 4068 17592
rect 3568 17552 3574 17564
rect 4062 17552 4068 17564
rect 4120 17552 4126 17604
rect 8128 17592 8156 17623
rect 9122 17620 9128 17672
rect 9180 17660 9186 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9180 17632 9781 17660
rect 9180 17620 9186 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9769 17623 9827 17629
rect 11164 17660 11192 17700
rect 11609 17697 11621 17731
rect 11655 17728 11667 17731
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 11655 17700 12081 17728
rect 11655 17697 11667 17700
rect 11609 17691 11667 17697
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 12710 17688 12716 17740
rect 12768 17728 12774 17740
rect 13004 17728 13032 17768
rect 15013 17765 15025 17768
rect 15059 17765 15071 17799
rect 15013 17759 15071 17765
rect 16850 17756 16856 17808
rect 16908 17796 16914 17808
rect 18598 17796 18604 17808
rect 16908 17768 18604 17796
rect 16908 17756 16914 17768
rect 18598 17756 18604 17768
rect 18656 17796 18662 17808
rect 19061 17799 19119 17805
rect 19061 17796 19073 17799
rect 18656 17768 19073 17796
rect 18656 17756 18662 17768
rect 19061 17765 19073 17768
rect 19107 17765 19119 17799
rect 19061 17759 19119 17765
rect 19978 17756 19984 17808
rect 20036 17796 20042 17808
rect 21082 17796 21088 17808
rect 20036 17768 21088 17796
rect 20036 17756 20042 17768
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 12768 17700 13032 17728
rect 12768 17688 12774 17700
rect 14274 17688 14280 17740
rect 14332 17728 14338 17740
rect 14461 17731 14519 17737
rect 14461 17728 14473 17731
rect 14332 17700 14473 17728
rect 14332 17688 14338 17700
rect 14461 17697 14473 17700
rect 14507 17697 14519 17731
rect 14461 17691 14519 17697
rect 15105 17731 15163 17737
rect 15105 17697 15117 17731
rect 15151 17728 15163 17731
rect 15378 17728 15384 17740
rect 15151 17700 15384 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 15378 17688 15384 17700
rect 15436 17688 15442 17740
rect 17313 17731 17371 17737
rect 17313 17697 17325 17731
rect 17359 17728 17371 17731
rect 17862 17728 17868 17740
rect 17359 17700 17868 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 17862 17688 17868 17700
rect 17920 17688 17926 17740
rect 18785 17731 18843 17737
rect 18785 17728 18797 17731
rect 18248 17700 18797 17728
rect 11333 17663 11391 17669
rect 11333 17660 11345 17663
rect 11164 17632 11345 17660
rect 8202 17592 8208 17604
rect 6564 17564 8208 17592
rect 6564 17536 6592 17564
rect 8202 17552 8208 17564
rect 8260 17552 8266 17604
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 3878 17484 3884 17536
rect 3936 17524 3942 17536
rect 6086 17524 6092 17536
rect 3936 17496 6092 17524
rect 3936 17484 3942 17496
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 6546 17524 6552 17536
rect 6507 17496 6552 17524
rect 6546 17484 6552 17496
rect 6604 17484 6610 17536
rect 7561 17527 7619 17533
rect 7561 17493 7573 17527
rect 7607 17524 7619 17527
rect 8294 17524 8300 17536
rect 7607 17496 8300 17524
rect 7607 17493 7619 17496
rect 7561 17487 7619 17493
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 9784 17524 9812 17623
rect 10686 17524 10692 17536
rect 9784 17496 10692 17524
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 11164 17524 11192 17632
rect 11333 17629 11345 17632
rect 11379 17629 11391 17663
rect 11333 17623 11391 17629
rect 11517 17663 11575 17669
rect 11517 17629 11529 17663
rect 11563 17660 11575 17663
rect 14090 17660 14096 17672
rect 11563 17632 14096 17660
rect 11563 17629 11575 17632
rect 11517 17623 11575 17629
rect 11238 17552 11244 17604
rect 11296 17592 11302 17604
rect 11532 17592 11560 17623
rect 14090 17620 14096 17632
rect 14148 17660 14154 17672
rect 14148 17632 14688 17660
rect 14148 17620 14154 17632
rect 11296 17564 11560 17592
rect 11296 17552 11302 17564
rect 11606 17552 11612 17604
rect 11664 17592 11670 17604
rect 14366 17592 14372 17604
rect 11664 17564 14372 17592
rect 11664 17552 11670 17564
rect 14366 17552 14372 17564
rect 14424 17552 14430 17604
rect 14660 17592 14688 17632
rect 14734 17620 14740 17672
rect 14792 17660 14798 17672
rect 14829 17663 14887 17669
rect 14829 17660 14841 17663
rect 14792 17632 14841 17660
rect 14792 17620 14798 17632
rect 14829 17629 14841 17632
rect 14875 17629 14887 17663
rect 14829 17623 14887 17629
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17660 15807 17663
rect 15930 17660 15936 17672
rect 15795 17632 15936 17660
rect 15795 17629 15807 17632
rect 15749 17623 15807 17629
rect 15930 17620 15936 17632
rect 15988 17620 15994 17672
rect 17129 17663 17187 17669
rect 17129 17629 17141 17663
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 16574 17592 16580 17604
rect 14660 17564 16580 17592
rect 16574 17552 16580 17564
rect 16632 17552 16638 17604
rect 17144 17592 17172 17623
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 17276 17632 17321 17660
rect 17276 17620 17282 17632
rect 17678 17620 17684 17672
rect 17736 17660 17742 17672
rect 18248 17669 18276 17700
rect 18785 17697 18797 17700
rect 18831 17728 18843 17731
rect 19150 17728 19156 17740
rect 18831 17700 19156 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 19150 17688 19156 17700
rect 19208 17688 19214 17740
rect 19426 17728 19432 17740
rect 19387 17700 19432 17728
rect 19426 17688 19432 17700
rect 19484 17688 19490 17740
rect 20073 17731 20131 17737
rect 20073 17697 20085 17731
rect 20119 17728 20131 17731
rect 20533 17731 20591 17737
rect 20533 17728 20545 17731
rect 20119 17700 20545 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 20533 17697 20545 17700
rect 20579 17697 20591 17731
rect 20533 17691 20591 17697
rect 20809 17731 20867 17737
rect 20809 17697 20821 17731
rect 20855 17697 20867 17731
rect 20809 17691 20867 17697
rect 18233 17663 18291 17669
rect 18233 17660 18245 17663
rect 17736 17632 18245 17660
rect 17736 17620 17742 17632
rect 18233 17629 18245 17632
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17629 18383 17663
rect 20165 17663 20223 17669
rect 20165 17660 20177 17663
rect 18325 17623 18383 17629
rect 18616 17632 20177 17660
rect 17310 17592 17316 17604
rect 17144 17564 17316 17592
rect 17310 17552 17316 17564
rect 17368 17592 17374 17604
rect 18340 17592 18368 17623
rect 17368 17564 18368 17592
rect 17368 17552 17374 17564
rect 16206 17524 16212 17536
rect 11164 17496 16212 17524
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 16482 17524 16488 17536
rect 16395 17496 16488 17524
rect 16482 17484 16488 17496
rect 16540 17524 16546 17536
rect 16850 17524 16856 17536
rect 16540 17496 16856 17524
rect 16540 17484 16546 17496
rect 16850 17484 16856 17496
rect 16908 17484 16914 17536
rect 18138 17484 18144 17536
rect 18196 17524 18202 17536
rect 18616 17533 18644 17632
rect 20165 17629 20177 17632
rect 20211 17629 20223 17663
rect 20346 17660 20352 17672
rect 20307 17632 20352 17660
rect 20165 17623 20223 17629
rect 20180 17592 20208 17623
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20824 17660 20852 17691
rect 20898 17688 20904 17740
rect 20956 17728 20962 17740
rect 21361 17731 21419 17737
rect 21361 17728 21373 17731
rect 20956 17700 21373 17728
rect 20956 17688 20962 17700
rect 21361 17697 21373 17700
rect 21407 17697 21419 17731
rect 21361 17691 21419 17697
rect 21082 17660 21088 17672
rect 20824 17632 21088 17660
rect 21082 17620 21088 17632
rect 21140 17620 21146 17672
rect 20622 17592 20628 17604
rect 20180 17564 20628 17592
rect 20622 17552 20628 17564
rect 20680 17552 20686 17604
rect 21542 17592 21548 17604
rect 21503 17564 21548 17592
rect 21542 17552 21548 17564
rect 21600 17552 21606 17604
rect 18601 17527 18659 17533
rect 18601 17524 18613 17527
rect 18196 17496 18613 17524
rect 18196 17484 18202 17496
rect 18601 17493 18613 17496
rect 18647 17493 18659 17527
rect 18601 17487 18659 17493
rect 19150 17484 19156 17536
rect 19208 17524 19214 17536
rect 19705 17527 19763 17533
rect 19705 17524 19717 17527
rect 19208 17496 19717 17524
rect 19208 17484 19214 17496
rect 19705 17493 19717 17496
rect 19751 17493 19763 17527
rect 20990 17524 20996 17536
rect 20951 17496 20996 17524
rect 19705 17487 19763 17493
rect 20990 17484 20996 17496
rect 21048 17484 21054 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 1765 17323 1823 17329
rect 1765 17289 1777 17323
rect 1811 17320 1823 17323
rect 1946 17320 1952 17332
rect 1811 17292 1952 17320
rect 1811 17289 1823 17292
rect 1765 17283 1823 17289
rect 1946 17280 1952 17292
rect 2004 17280 2010 17332
rect 2409 17323 2467 17329
rect 2409 17289 2421 17323
rect 2455 17320 2467 17323
rect 3878 17320 3884 17332
rect 2455 17292 3884 17320
rect 2455 17289 2467 17292
rect 2409 17283 2467 17289
rect 1578 17212 1584 17264
rect 1636 17252 1642 17264
rect 2041 17255 2099 17261
rect 2041 17252 2053 17255
rect 1636 17224 2053 17252
rect 1636 17212 1642 17224
rect 2041 17221 2053 17224
rect 2087 17221 2099 17255
rect 2041 17215 2099 17221
rect 2424 17184 2452 17283
rect 3878 17280 3884 17292
rect 3936 17280 3942 17332
rect 3988 17292 5120 17320
rect 3988 17252 4016 17292
rect 1964 17156 2452 17184
rect 2746 17224 4016 17252
rect 1964 17125 1992 17156
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17085 2007 17119
rect 1949 17079 2007 17085
rect 2225 17119 2283 17125
rect 2225 17085 2237 17119
rect 2271 17116 2283 17119
rect 2593 17119 2651 17125
rect 2593 17116 2605 17119
rect 2271 17088 2605 17116
rect 2271 17085 2283 17088
rect 2225 17079 2283 17085
rect 2593 17085 2605 17088
rect 2639 17116 2651 17119
rect 2746 17116 2774 17224
rect 2866 17144 2872 17196
rect 2924 17184 2930 17196
rect 3145 17187 3203 17193
rect 3145 17184 3157 17187
rect 2924 17156 3157 17184
rect 2924 17144 2930 17156
rect 3145 17153 3157 17156
rect 3191 17153 3203 17187
rect 5092 17184 5120 17292
rect 5166 17280 5172 17332
rect 5224 17320 5230 17332
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 5224 17292 5457 17320
rect 5224 17280 5230 17292
rect 5445 17289 5457 17292
rect 5491 17289 5503 17323
rect 5445 17283 5503 17289
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 8297 17323 8355 17329
rect 8297 17320 8309 17323
rect 6972 17292 8309 17320
rect 6972 17280 6978 17292
rect 5350 17252 5356 17264
rect 5311 17224 5356 17252
rect 5350 17212 5356 17224
rect 5408 17252 5414 17264
rect 5810 17252 5816 17264
rect 5408 17224 5816 17252
rect 5408 17212 5414 17224
rect 5810 17212 5816 17224
rect 5868 17212 5874 17264
rect 5920 17224 6408 17252
rect 5920 17184 5948 17224
rect 5092 17156 5948 17184
rect 3145 17147 3203 17153
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 6380 17184 6408 17224
rect 6454 17212 6460 17264
rect 6512 17252 6518 17264
rect 6822 17252 6828 17264
rect 6512 17224 6828 17252
rect 6512 17212 6518 17224
rect 6822 17212 6828 17224
rect 6880 17212 6886 17264
rect 8036 17184 8064 17292
rect 8297 17289 8309 17292
rect 8343 17289 8355 17323
rect 8297 17283 8355 17289
rect 8570 17280 8576 17332
rect 8628 17320 8634 17332
rect 8628 17292 9904 17320
rect 8628 17280 8634 17292
rect 9769 17255 9827 17261
rect 9769 17221 9781 17255
rect 9815 17221 9827 17255
rect 9876 17252 9904 17292
rect 10410 17280 10416 17332
rect 10468 17320 10474 17332
rect 10778 17320 10784 17332
rect 10468 17292 10784 17320
rect 10468 17280 10474 17292
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 11149 17323 11207 17329
rect 11149 17289 11161 17323
rect 11195 17320 11207 17323
rect 11238 17320 11244 17332
rect 11195 17292 11244 17320
rect 11195 17289 11207 17292
rect 11149 17283 11207 17289
rect 11238 17280 11244 17292
rect 11296 17280 11302 17332
rect 12989 17323 13047 17329
rect 12989 17289 13001 17323
rect 13035 17320 13047 17323
rect 13906 17320 13912 17332
rect 13035 17292 13912 17320
rect 13035 17289 13047 17292
rect 12989 17283 13047 17289
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 14366 17280 14372 17332
rect 14424 17320 14430 17332
rect 15378 17320 15384 17332
rect 14424 17292 15384 17320
rect 14424 17280 14430 17292
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 16298 17280 16304 17332
rect 16356 17320 16362 17332
rect 16393 17323 16451 17329
rect 16393 17320 16405 17323
rect 16356 17292 16405 17320
rect 16356 17280 16362 17292
rect 16393 17289 16405 17292
rect 16439 17289 16451 17323
rect 16393 17283 16451 17289
rect 17126 17280 17132 17332
rect 17184 17320 17190 17332
rect 17405 17323 17463 17329
rect 17405 17320 17417 17323
rect 17184 17292 17417 17320
rect 17184 17280 17190 17292
rect 17405 17289 17417 17292
rect 17451 17289 17463 17323
rect 17405 17283 17463 17289
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 18693 17323 18751 17329
rect 18693 17320 18705 17323
rect 17644 17292 18705 17320
rect 17644 17280 17650 17292
rect 18693 17289 18705 17292
rect 18739 17320 18751 17323
rect 19058 17320 19064 17332
rect 18739 17292 19064 17320
rect 18739 17289 18751 17292
rect 18693 17283 18751 17289
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 19337 17323 19395 17329
rect 19337 17289 19349 17323
rect 19383 17320 19395 17323
rect 20438 17320 20444 17332
rect 19383 17292 20444 17320
rect 19383 17289 19395 17292
rect 19337 17283 19395 17289
rect 20438 17280 20444 17292
rect 20496 17280 20502 17332
rect 17218 17252 17224 17264
rect 9876 17224 13400 17252
rect 9769 17215 9827 17221
rect 9784 17184 9812 17215
rect 10505 17187 10563 17193
rect 10505 17184 10517 17187
rect 6052 17156 6097 17184
rect 6380 17156 7052 17184
rect 8036 17156 8524 17184
rect 9784 17156 10517 17184
rect 6052 17144 6058 17156
rect 2639 17088 2774 17116
rect 3421 17119 3479 17125
rect 2639 17085 2651 17088
rect 2593 17079 2651 17085
rect 3421 17085 3433 17119
rect 3467 17116 3479 17119
rect 3786 17116 3792 17128
rect 3467 17088 3792 17116
rect 3467 17085 3479 17088
rect 3421 17079 3479 17085
rect 3786 17076 3792 17088
rect 3844 17076 3850 17128
rect 3878 17076 3884 17128
rect 3936 17116 3942 17128
rect 3973 17119 4031 17125
rect 3973 17116 3985 17119
rect 3936 17088 3985 17116
rect 3936 17076 3942 17088
rect 3973 17085 3985 17088
rect 4019 17085 4031 17119
rect 3973 17079 4031 17085
rect 4172 17088 6132 17116
rect 1394 17048 1400 17060
rect 1355 17020 1400 17048
rect 1394 17008 1400 17020
rect 1452 17008 1458 17060
rect 1578 17048 1584 17060
rect 1539 17020 1584 17048
rect 1578 17008 1584 17020
rect 1636 17008 1642 17060
rect 2958 17008 2964 17060
rect 3016 17048 3022 17060
rect 4172 17048 4200 17088
rect 3016 17020 4200 17048
rect 4240 17051 4298 17057
rect 3016 17008 3022 17020
rect 4240 17017 4252 17051
rect 4286 17048 4298 17051
rect 4338 17048 4344 17060
rect 4286 17020 4344 17048
rect 4286 17017 4298 17020
rect 4240 17011 4298 17017
rect 4338 17008 4344 17020
rect 4396 17008 4402 17060
rect 5810 17048 5816 17060
rect 5771 17020 5816 17048
rect 5810 17008 5816 17020
rect 5868 17008 5874 17060
rect 3326 16980 3332 16992
rect 3287 16952 3332 16980
rect 3326 16940 3332 16952
rect 3384 16940 3390 16992
rect 3789 16983 3847 16989
rect 3789 16949 3801 16983
rect 3835 16980 3847 16983
rect 4154 16980 4160 16992
rect 3835 16952 4160 16980
rect 3835 16949 3847 16952
rect 3789 16943 3847 16949
rect 4154 16940 4160 16952
rect 4212 16940 4218 16992
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 5905 16983 5963 16989
rect 5905 16980 5917 16983
rect 5592 16952 5917 16980
rect 5592 16940 5598 16952
rect 5905 16949 5917 16952
rect 5951 16949 5963 16983
rect 6104 16980 6132 17088
rect 6178 17076 6184 17128
rect 6236 17116 6242 17128
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 6236 17088 6929 17116
rect 6236 17076 6242 17088
rect 6917 17085 6929 17088
rect 6963 17085 6975 17119
rect 7024 17116 7052 17156
rect 8294 17116 8300 17128
rect 7024 17088 8300 17116
rect 6917 17079 6975 17085
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 8389 17119 8447 17125
rect 8389 17085 8401 17119
rect 8435 17085 8447 17119
rect 8496 17116 8524 17156
rect 10505 17153 10517 17156
rect 10551 17184 10563 17187
rect 10778 17184 10784 17196
rect 10551 17156 10784 17184
rect 10551 17153 10563 17156
rect 10505 17147 10563 17153
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 13262 17184 13268 17196
rect 13223 17156 13268 17184
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 13372 17193 13400 17224
rect 14016 17224 17224 17252
rect 13357 17187 13415 17193
rect 13357 17153 13369 17187
rect 13403 17184 13415 17187
rect 13538 17184 13544 17196
rect 13403 17156 13544 17184
rect 13403 17153 13415 17156
rect 13357 17147 13415 17153
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 8645 17119 8703 17125
rect 8645 17116 8657 17119
rect 8496 17088 8657 17116
rect 8389 17079 8447 17085
rect 8645 17085 8657 17088
rect 8691 17085 8703 17119
rect 8645 17079 8703 17085
rect 7184 17051 7242 17057
rect 7184 17017 7196 17051
rect 7230 17048 7242 17051
rect 7558 17048 7564 17060
rect 7230 17020 7564 17048
rect 7230 17017 7242 17020
rect 7184 17011 7242 17017
rect 7558 17008 7564 17020
rect 7616 17008 7622 17060
rect 8404 17048 8432 17079
rect 9398 17076 9404 17128
rect 9456 17116 9462 17128
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 9456 17088 10333 17116
rect 9456 17076 9462 17088
rect 10321 17085 10333 17088
rect 10367 17085 10379 17119
rect 10321 17079 10379 17085
rect 11606 17076 11612 17128
rect 11664 17116 11670 17128
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 11664 17088 12817 17116
rect 11664 17076 11670 17088
rect 12805 17085 12817 17088
rect 12851 17085 12863 17119
rect 13449 17119 13507 17125
rect 13449 17116 13461 17119
rect 12805 17079 12863 17085
rect 12912 17088 13461 17116
rect 9122 17048 9128 17060
rect 8404 17020 9128 17048
rect 9122 17008 9128 17020
rect 9180 17008 9186 17060
rect 9582 17008 9588 17060
rect 9640 17048 9646 17060
rect 10229 17051 10287 17057
rect 10229 17048 10241 17051
rect 9640 17020 10241 17048
rect 9640 17008 9646 17020
rect 10229 17017 10241 17020
rect 10275 17048 10287 17051
rect 12710 17048 12716 17060
rect 10275 17020 12716 17048
rect 10275 17017 10287 17020
rect 10229 17011 10287 17017
rect 12710 17008 12716 17020
rect 12768 17008 12774 17060
rect 9766 16980 9772 16992
rect 6104 16952 9772 16980
rect 5905 16943 5963 16949
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 9858 16940 9864 16992
rect 9916 16980 9922 16992
rect 9916 16952 9961 16980
rect 9916 16940 9922 16952
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 12912 16980 12940 17088
rect 13449 17085 13461 17088
rect 13495 17116 13507 17119
rect 14016 17116 14044 17224
rect 17218 17212 17224 17224
rect 17276 17212 17282 17264
rect 17862 17252 17868 17264
rect 17823 17224 17868 17252
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 18046 17252 18052 17264
rect 18007 17224 18052 17252
rect 18046 17212 18052 17224
rect 18104 17212 18110 17264
rect 18325 17255 18383 17261
rect 18325 17221 18337 17255
rect 18371 17252 18383 17255
rect 18598 17252 18604 17264
rect 18371 17224 18604 17252
rect 18371 17221 18383 17224
rect 18325 17215 18383 17221
rect 18598 17212 18604 17224
rect 18656 17212 18662 17264
rect 19429 17255 19487 17261
rect 19429 17221 19441 17255
rect 19475 17221 19487 17255
rect 19429 17215 19487 17221
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17184 15163 17187
rect 15286 17184 15292 17196
rect 15151 17156 15292 17184
rect 15151 17153 15163 17156
rect 15105 17147 15163 17153
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 16206 17144 16212 17196
rect 16264 17184 16270 17196
rect 19444 17184 19472 17215
rect 16264 17156 19472 17184
rect 16264 17144 16270 17156
rect 13495 17088 14044 17116
rect 14093 17119 14151 17125
rect 13495 17085 13507 17088
rect 13449 17079 13507 17085
rect 14093 17085 14105 17119
rect 14139 17116 14151 17119
rect 16482 17116 16488 17128
rect 14139 17088 16488 17116
rect 14139 17085 14151 17088
rect 14093 17079 14151 17085
rect 16482 17076 16488 17088
rect 16540 17076 16546 17128
rect 16574 17076 16580 17128
rect 16632 17116 16638 17128
rect 17589 17119 17647 17125
rect 16632 17088 16677 17116
rect 16632 17076 16638 17088
rect 17589 17085 17601 17119
rect 17635 17116 17647 17119
rect 18690 17116 18696 17128
rect 17635 17088 18696 17116
rect 17635 17085 17647 17088
rect 17589 17079 17647 17085
rect 18690 17076 18696 17088
rect 18748 17076 18754 17128
rect 18966 17116 18972 17128
rect 18927 17088 18972 17116
rect 18966 17076 18972 17088
rect 19024 17116 19030 17128
rect 19153 17119 19211 17125
rect 19153 17116 19165 17119
rect 19024 17088 19165 17116
rect 19024 17076 19030 17088
rect 19153 17085 19165 17088
rect 19199 17085 19211 17119
rect 19153 17079 19211 17085
rect 20809 17119 20867 17125
rect 20809 17085 20821 17119
rect 20855 17085 20867 17119
rect 20990 17116 20996 17128
rect 20951 17088 20996 17116
rect 20809 17079 20867 17085
rect 15013 17051 15071 17057
rect 15013 17048 15025 17051
rect 14384 17020 15025 17048
rect 14384 16992 14412 17020
rect 15013 17017 15025 17020
rect 15059 17017 15071 17051
rect 15013 17011 15071 17017
rect 17126 17008 17132 17060
rect 17184 17048 17190 17060
rect 17184 17020 17816 17048
rect 17184 17008 17190 17020
rect 10192 16952 12940 16980
rect 10192 16940 10198 16952
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 13817 16983 13875 16989
rect 13817 16980 13829 16983
rect 13780 16952 13829 16980
rect 13780 16940 13786 16952
rect 13817 16949 13829 16952
rect 13863 16949 13875 16983
rect 13817 16943 13875 16949
rect 13906 16940 13912 16992
rect 13964 16980 13970 16992
rect 14366 16980 14372 16992
rect 13964 16952 14009 16980
rect 14327 16952 14372 16980
rect 13964 16940 13970 16952
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 14550 16980 14556 16992
rect 14511 16952 14556 16980
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 14734 16940 14740 16992
rect 14792 16980 14798 16992
rect 14921 16983 14979 16989
rect 14921 16980 14933 16983
rect 14792 16952 14933 16980
rect 14792 16940 14798 16952
rect 14921 16949 14933 16952
rect 14967 16949 14979 16983
rect 14921 16943 14979 16949
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 15657 16983 15715 16989
rect 15657 16980 15669 16983
rect 15436 16952 15669 16980
rect 15436 16940 15442 16952
rect 15657 16949 15669 16952
rect 15703 16980 15715 16983
rect 17034 16980 17040 16992
rect 15703 16952 17040 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 17218 16940 17224 16992
rect 17276 16980 17282 16992
rect 17678 16980 17684 16992
rect 17276 16952 17684 16980
rect 17276 16940 17282 16952
rect 17678 16940 17684 16952
rect 17736 16940 17742 16992
rect 17788 16980 17816 17020
rect 18138 17008 18144 17060
rect 18196 17048 18202 17060
rect 18785 17051 18843 17057
rect 18785 17048 18797 17051
rect 18196 17020 18797 17048
rect 18196 17008 18202 17020
rect 18785 17017 18797 17020
rect 18831 17017 18843 17051
rect 18785 17011 18843 17017
rect 19610 17008 19616 17060
rect 19668 17048 19674 17060
rect 20542 17051 20600 17057
rect 20542 17048 20554 17051
rect 19668 17020 20554 17048
rect 19668 17008 19674 17020
rect 20542 17017 20554 17020
rect 20588 17017 20600 17051
rect 20542 17011 20600 17017
rect 18417 16983 18475 16989
rect 18417 16980 18429 16983
rect 17788 16952 18429 16980
rect 18417 16949 18429 16952
rect 18463 16980 18475 16983
rect 19518 16980 19524 16992
rect 18463 16952 19524 16980
rect 18463 16949 18475 16952
rect 18417 16943 18475 16949
rect 19518 16940 19524 16952
rect 19576 16980 19582 16992
rect 19886 16980 19892 16992
rect 19576 16952 19892 16980
rect 19576 16940 19582 16952
rect 19886 16940 19892 16952
rect 19944 16940 19950 16992
rect 20824 16980 20852 17079
rect 20990 17076 20996 17088
rect 21048 17076 21054 17128
rect 21174 17048 21180 17060
rect 21135 17020 21180 17048
rect 21174 17008 21180 17020
rect 21232 17008 21238 17060
rect 21358 17048 21364 17060
rect 21319 17020 21364 17048
rect 21358 17008 21364 17020
rect 21416 17008 21422 17060
rect 20990 16980 20996 16992
rect 20824 16952 20996 16980
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 21450 16980 21456 16992
rect 21411 16952 21456 16980
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 2958 16736 2964 16788
rect 3016 16776 3022 16788
rect 3237 16779 3295 16785
rect 3237 16776 3249 16779
rect 3016 16748 3249 16776
rect 3016 16736 3022 16748
rect 3237 16745 3249 16748
rect 3283 16745 3295 16779
rect 3237 16739 3295 16745
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 3605 16779 3663 16785
rect 3605 16776 3617 16779
rect 3384 16748 3617 16776
rect 3384 16736 3390 16748
rect 3605 16745 3617 16748
rect 3651 16745 3663 16779
rect 3605 16739 3663 16745
rect 5718 16736 5724 16788
rect 5776 16776 5782 16788
rect 5813 16779 5871 16785
rect 5813 16776 5825 16779
rect 5776 16748 5825 16776
rect 5776 16736 5782 16748
rect 5813 16745 5825 16748
rect 5859 16776 5871 16779
rect 9582 16776 9588 16788
rect 5859 16748 7512 16776
rect 5859 16745 5871 16748
rect 5813 16739 5871 16745
rect 6448 16711 6506 16717
rect 3160 16680 6408 16708
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16640 1639 16643
rect 1946 16640 1952 16652
rect 1627 16612 1952 16640
rect 1627 16609 1639 16612
rect 1581 16603 1639 16609
rect 1946 16600 1952 16612
rect 2004 16600 2010 16652
rect 2682 16640 2688 16652
rect 2595 16612 2688 16640
rect 2682 16600 2688 16612
rect 2740 16640 2746 16652
rect 3160 16649 3188 16680
rect 3145 16643 3203 16649
rect 3145 16640 3157 16643
rect 2740 16612 3157 16640
rect 2740 16600 2746 16612
rect 3145 16609 3157 16612
rect 3191 16609 3203 16643
rect 3145 16603 3203 16609
rect 3970 16600 3976 16652
rect 4028 16640 4034 16652
rect 4148 16643 4206 16649
rect 4148 16640 4160 16643
rect 4028 16612 4160 16640
rect 4028 16600 4034 16612
rect 4148 16609 4160 16612
rect 4194 16640 4206 16643
rect 5721 16643 5779 16649
rect 4194 16612 4936 16640
rect 4194 16609 4206 16612
rect 4148 16603 4206 16609
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16541 3111 16575
rect 3878 16572 3884 16584
rect 3839 16544 3884 16572
rect 3053 16535 3111 16541
rect 3068 16504 3096 16535
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 3694 16504 3700 16516
rect 3068 16476 3700 16504
rect 3694 16464 3700 16476
rect 3752 16464 3758 16516
rect 4908 16504 4936 16612
rect 5721 16609 5733 16643
rect 5767 16640 5779 16643
rect 6270 16640 6276 16652
rect 5767 16612 6276 16640
rect 5767 16609 5779 16612
rect 5721 16603 5779 16609
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 6380 16640 6408 16680
rect 6448 16677 6460 16711
rect 6494 16708 6506 16711
rect 6546 16708 6552 16720
rect 6494 16680 6552 16708
rect 6494 16677 6506 16680
rect 6448 16671 6506 16677
rect 6546 16668 6552 16680
rect 6604 16668 6610 16720
rect 7484 16708 7512 16748
rect 7668 16748 9588 16776
rect 7668 16708 7696 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 10413 16779 10471 16785
rect 10413 16776 10425 16779
rect 9824 16748 10425 16776
rect 9824 16736 9830 16748
rect 10413 16745 10425 16748
rect 10459 16776 10471 16779
rect 10594 16776 10600 16788
rect 10459 16748 10600 16776
rect 10459 16745 10471 16748
rect 10413 16739 10471 16745
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 11606 16776 11612 16788
rect 11567 16748 11612 16776
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 12894 16776 12900 16788
rect 12855 16748 12900 16776
rect 12894 16736 12900 16748
rect 12952 16736 12958 16788
rect 13265 16779 13323 16785
rect 13265 16745 13277 16779
rect 13311 16745 13323 16779
rect 13722 16776 13728 16788
rect 13683 16748 13728 16776
rect 13265 16739 13323 16745
rect 7484 16680 7696 16708
rect 7760 16680 10272 16708
rect 7760 16640 7788 16680
rect 6380 16612 7788 16640
rect 7834 16600 7840 16652
rect 7892 16640 7898 16652
rect 8021 16643 8079 16649
rect 8021 16640 8033 16643
rect 7892 16612 8033 16640
rect 7892 16600 7898 16612
rect 8021 16609 8033 16612
rect 8067 16640 8079 16643
rect 9214 16640 9220 16652
rect 8067 16612 9076 16640
rect 9175 16612 9220 16640
rect 8067 16609 8079 16612
rect 8021 16603 8079 16609
rect 5994 16572 6000 16584
rect 5955 16544 6000 16572
rect 5994 16532 6000 16544
rect 6052 16532 6058 16584
rect 6178 16572 6184 16584
rect 6139 16544 6184 16572
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 8110 16572 8116 16584
rect 8071 16544 8116 16572
rect 8110 16532 8116 16544
rect 8168 16532 8174 16584
rect 8202 16532 8208 16584
rect 8260 16572 8266 16584
rect 9048 16572 9076 16612
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 10134 16640 10140 16652
rect 9324 16612 10140 16640
rect 9324 16572 9352 16612
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 8260 16544 8305 16572
rect 9048 16544 9352 16572
rect 9953 16575 10011 16581
rect 8260 16532 8266 16544
rect 9953 16541 9965 16575
rect 9999 16572 10011 16575
rect 10244 16572 10272 16680
rect 10962 16668 10968 16720
rect 11020 16708 11026 16720
rect 12345 16711 12403 16717
rect 12345 16708 12357 16711
rect 11020 16680 12357 16708
rect 11020 16668 11026 16680
rect 12345 16677 12357 16680
rect 12391 16708 12403 16711
rect 12805 16711 12863 16717
rect 12805 16708 12817 16711
rect 12391 16680 12817 16708
rect 12391 16677 12403 16680
rect 12345 16671 12403 16677
rect 12805 16677 12817 16680
rect 12851 16708 12863 16711
rect 13280 16708 13308 16739
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 14093 16779 14151 16785
rect 14093 16745 14105 16779
rect 14139 16776 14151 16779
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 14139 16748 16313 16776
rect 14139 16745 14151 16748
rect 14093 16739 14151 16745
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 16301 16739 16359 16745
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 16853 16779 16911 16785
rect 16853 16776 16865 16779
rect 16632 16748 16865 16776
rect 16632 16736 16638 16748
rect 16853 16745 16865 16748
rect 16899 16745 16911 16779
rect 16853 16739 16911 16745
rect 17034 16736 17040 16788
rect 17092 16776 17098 16788
rect 18690 16776 18696 16788
rect 17092 16748 18184 16776
rect 18651 16748 18696 16776
rect 17092 16736 17098 16748
rect 13633 16711 13691 16717
rect 13633 16708 13645 16711
rect 12851 16680 13216 16708
rect 13280 16680 13645 16708
rect 12851 16677 12863 16680
rect 12805 16671 12863 16677
rect 11238 16640 11244 16652
rect 11199 16612 11244 16640
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 13078 16640 13084 16652
rect 12728 16612 13084 16640
rect 10505 16575 10563 16581
rect 10505 16572 10517 16575
rect 9999 16544 10517 16572
rect 9999 16541 10011 16544
rect 9953 16535 10011 16541
rect 10505 16541 10517 16544
rect 10551 16572 10563 16575
rect 10594 16572 10600 16584
rect 10551 16544 10600 16572
rect 10551 16541 10563 16544
rect 10505 16535 10563 16541
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 10689 16575 10747 16581
rect 10689 16541 10701 16575
rect 10735 16572 10747 16575
rect 10778 16572 10784 16584
rect 10735 16544 10784 16572
rect 10735 16541 10747 16544
rect 10689 16535 10747 16541
rect 10778 16532 10784 16544
rect 10836 16532 10842 16584
rect 11054 16572 11060 16584
rect 11015 16544 11060 16572
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 12728 16581 12756 16612
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 13188 16640 13216 16680
rect 13633 16677 13645 16680
rect 13679 16677 13691 16711
rect 17126 16708 17132 16720
rect 13633 16671 13691 16677
rect 13740 16680 17132 16708
rect 13740 16640 13768 16680
rect 17126 16668 17132 16680
rect 17184 16668 17190 16720
rect 17221 16711 17279 16717
rect 17221 16677 17233 16711
rect 17267 16708 17279 16711
rect 18046 16708 18052 16720
rect 17267 16680 18052 16708
rect 17267 16677 17279 16680
rect 17221 16671 17279 16677
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 14625 16643 14683 16649
rect 14625 16640 14637 16643
rect 13188 16612 13768 16640
rect 13832 16612 14637 16640
rect 13832 16584 13860 16612
rect 14625 16609 14637 16612
rect 14671 16609 14683 16643
rect 14625 16603 14683 16609
rect 15378 16600 15384 16652
rect 15436 16640 15442 16652
rect 16209 16643 16267 16649
rect 16209 16640 16221 16643
rect 15436 16612 16221 16640
rect 15436 16600 15442 16612
rect 16209 16609 16221 16612
rect 16255 16609 16267 16643
rect 17310 16640 17316 16652
rect 17271 16612 17316 16640
rect 16209 16603 16267 16609
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 18156 16640 18184 16748
rect 18690 16736 18696 16748
rect 18748 16736 18754 16788
rect 19061 16779 19119 16785
rect 19061 16745 19073 16779
rect 19107 16776 19119 16779
rect 19150 16776 19156 16788
rect 19107 16748 19156 16776
rect 19107 16745 19119 16748
rect 19061 16739 19119 16745
rect 19150 16736 19156 16748
rect 19208 16736 19214 16788
rect 19610 16776 19616 16788
rect 19571 16748 19616 16776
rect 19610 16736 19616 16748
rect 19668 16736 19674 16788
rect 20714 16736 20720 16788
rect 20772 16736 20778 16788
rect 21082 16776 21088 16788
rect 21043 16748 21088 16776
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 18601 16711 18659 16717
rect 18601 16677 18613 16711
rect 18647 16708 18659 16711
rect 18874 16708 18880 16720
rect 18647 16680 18880 16708
rect 18647 16677 18659 16680
rect 18601 16671 18659 16677
rect 18874 16668 18880 16680
rect 18932 16668 18938 16720
rect 20732 16708 20760 16736
rect 19168 16680 20760 16708
rect 19168 16649 19196 16680
rect 19153 16643 19211 16649
rect 18156 16612 19104 16640
rect 11149 16575 11207 16581
rect 11149 16541 11161 16575
rect 11195 16541 11207 16575
rect 11149 16535 11207 16541
rect 12713 16575 12771 16581
rect 12713 16541 12725 16575
rect 12759 16541 12771 16575
rect 12713 16535 12771 16541
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16572 13599 16575
rect 13814 16572 13820 16584
rect 13587 16544 13820 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 6012 16504 6040 16532
rect 7558 16504 7564 16516
rect 4908 16476 6040 16504
rect 7519 16476 7564 16504
rect 7558 16464 7564 16476
rect 7616 16464 7622 16516
rect 7650 16464 7656 16516
rect 7708 16504 7714 16516
rect 7708 16476 7753 16504
rect 7708 16464 7714 16476
rect 7834 16464 7840 16516
rect 7892 16504 7898 16516
rect 8386 16504 8392 16516
rect 7892 16476 8392 16504
rect 7892 16464 7898 16476
rect 8386 16464 8392 16476
rect 8444 16464 8450 16516
rect 10226 16464 10232 16516
rect 10284 16504 10290 16516
rect 11164 16504 11192 16535
rect 13814 16532 13820 16544
rect 13872 16532 13878 16584
rect 13906 16532 13912 16584
rect 13964 16572 13970 16584
rect 14369 16575 14427 16581
rect 14369 16572 14381 16575
rect 13964 16544 14381 16572
rect 13964 16532 13970 16544
rect 14369 16541 14381 16544
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 15930 16532 15936 16584
rect 15988 16572 15994 16584
rect 16393 16575 16451 16581
rect 16393 16572 16405 16575
rect 15988 16544 16405 16572
rect 15988 16532 15994 16544
rect 16393 16541 16405 16544
rect 16439 16541 16451 16575
rect 17494 16572 17500 16584
rect 17455 16544 17500 16572
rect 16393 16535 16451 16541
rect 17494 16532 17500 16544
rect 17552 16532 17558 16584
rect 15841 16507 15899 16513
rect 15841 16504 15853 16507
rect 10284 16476 11192 16504
rect 15304 16476 15853 16504
rect 10284 16464 10290 16476
rect 2038 16436 2044 16448
rect 1999 16408 2044 16436
rect 2038 16396 2044 16408
rect 2096 16396 2102 16448
rect 5258 16436 5264 16448
rect 5219 16408 5264 16436
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 5350 16396 5356 16448
rect 5408 16436 5414 16448
rect 5408 16408 5453 16436
rect 5408 16396 5414 16408
rect 8110 16396 8116 16448
rect 8168 16436 8174 16448
rect 8478 16436 8484 16448
rect 8168 16408 8484 16436
rect 8168 16396 8174 16408
rect 8478 16396 8484 16408
rect 8536 16396 8542 16448
rect 9122 16396 9128 16448
rect 9180 16436 9186 16448
rect 9401 16439 9459 16445
rect 9401 16436 9413 16439
rect 9180 16408 9413 16436
rect 9180 16396 9186 16408
rect 9401 16405 9413 16408
rect 9447 16405 9459 16439
rect 9401 16399 9459 16405
rect 9950 16396 9956 16448
rect 10008 16436 10014 16448
rect 10045 16439 10103 16445
rect 10045 16436 10057 16439
rect 10008 16408 10057 16436
rect 10008 16396 10014 16408
rect 10045 16405 10057 16408
rect 10091 16405 10103 16439
rect 10045 16399 10103 16405
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 15304 16436 15332 16476
rect 15841 16473 15853 16476
rect 15887 16473 15899 16507
rect 19076 16504 19104 16612
rect 19153 16609 19165 16643
rect 19199 16609 19211 16643
rect 19153 16603 19211 16609
rect 20346 16600 20352 16652
rect 20404 16640 20410 16652
rect 20726 16643 20784 16649
rect 20726 16640 20738 16643
rect 20404 16612 20738 16640
rect 20404 16600 20410 16612
rect 20726 16609 20738 16612
rect 20772 16609 20784 16643
rect 20726 16603 20784 16609
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 21361 16643 21419 16649
rect 21361 16640 21373 16643
rect 20956 16612 21373 16640
rect 20956 16600 20962 16612
rect 21361 16609 21373 16612
rect 21407 16609 21419 16643
rect 21542 16640 21548 16652
rect 21503 16612 21548 16640
rect 21361 16603 21419 16609
rect 21542 16600 21548 16612
rect 21600 16600 21606 16652
rect 19245 16575 19303 16581
rect 19245 16541 19257 16575
rect 19291 16572 19303 16575
rect 19610 16572 19616 16584
rect 19291 16544 19616 16572
rect 19291 16541 19303 16544
rect 19245 16535 19303 16541
rect 19610 16532 19616 16544
rect 19668 16532 19674 16584
rect 20990 16572 20996 16584
rect 20951 16544 20996 16572
rect 20990 16532 20996 16544
rect 21048 16532 21054 16584
rect 19076 16476 19380 16504
rect 15841 16467 15899 16473
rect 15746 16436 15752 16448
rect 14332 16408 15332 16436
rect 15707 16408 15752 16436
rect 14332 16396 14338 16408
rect 15746 16396 15752 16408
rect 15804 16396 15810 16448
rect 17402 16396 17408 16448
rect 17460 16436 17466 16448
rect 17773 16439 17831 16445
rect 17773 16436 17785 16439
rect 17460 16408 17785 16436
rect 17460 16396 17466 16408
rect 17773 16405 17785 16408
rect 17819 16405 17831 16439
rect 19352 16436 19380 16476
rect 21726 16436 21732 16448
rect 19352 16408 21732 16436
rect 17773 16399 17831 16405
rect 21726 16396 21732 16408
rect 21784 16396 21790 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 1765 16235 1823 16241
rect 1765 16232 1777 16235
rect 1636 16204 1777 16232
rect 1636 16192 1642 16204
rect 1765 16201 1777 16204
rect 1811 16201 1823 16235
rect 1765 16195 1823 16201
rect 2409 16235 2467 16241
rect 2409 16201 2421 16235
rect 2455 16232 2467 16235
rect 2866 16232 2872 16244
rect 2455 16204 2872 16232
rect 2455 16201 2467 16204
rect 2409 16195 2467 16201
rect 2866 16192 2872 16204
rect 2924 16232 2930 16244
rect 3970 16232 3976 16244
rect 2924 16204 3976 16232
rect 2924 16192 2930 16204
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 5810 16232 5816 16244
rect 4908 16204 5672 16232
rect 5771 16204 5816 16232
rect 2038 16124 2044 16176
rect 2096 16164 2102 16176
rect 2096 16136 2774 16164
rect 2096 16124 2102 16136
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 2038 16028 2044 16040
rect 1995 16000 2044 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 2038 15988 2044 16000
rect 2096 15988 2102 16040
rect 2225 16031 2283 16037
rect 2225 15997 2237 16031
rect 2271 16028 2283 16031
rect 2314 16028 2320 16040
rect 2271 16000 2320 16028
rect 2271 15997 2283 16000
rect 2225 15991 2283 15997
rect 2314 15988 2320 16000
rect 2372 15988 2378 16040
rect 2746 16028 2774 16136
rect 3786 16124 3792 16176
rect 3844 16164 3850 16176
rect 4908 16164 4936 16204
rect 3844 16136 4936 16164
rect 4985 16167 5043 16173
rect 3844 16124 3850 16136
rect 4985 16133 4997 16167
rect 5031 16164 5043 16167
rect 5534 16164 5540 16176
rect 5031 16136 5540 16164
rect 5031 16133 5043 16136
rect 4985 16127 5043 16133
rect 5534 16124 5540 16136
rect 5592 16124 5598 16176
rect 5644 16164 5672 16204
rect 5810 16192 5816 16204
rect 5868 16192 5874 16244
rect 6825 16235 6883 16241
rect 6825 16201 6837 16235
rect 6871 16232 6883 16235
rect 7098 16232 7104 16244
rect 6871 16204 7104 16232
rect 6871 16201 6883 16204
rect 6825 16195 6883 16201
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 9953 16235 10011 16241
rect 9953 16201 9965 16235
rect 9999 16232 10011 16235
rect 10226 16232 10232 16244
rect 9999 16204 10232 16232
rect 9999 16201 10011 16204
rect 9953 16195 10011 16201
rect 10226 16192 10232 16204
rect 10284 16192 10290 16244
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11425 16235 11483 16241
rect 11425 16232 11437 16235
rect 11112 16204 11437 16232
rect 11112 16192 11118 16204
rect 11425 16201 11437 16204
rect 11471 16201 11483 16235
rect 11425 16195 11483 16201
rect 8846 16164 8852 16176
rect 5644 16136 8852 16164
rect 8846 16124 8852 16136
rect 8904 16124 8910 16176
rect 9122 16124 9128 16176
rect 9180 16164 9186 16176
rect 9180 16136 10088 16164
rect 9180 16124 9186 16136
rect 3804 16096 3832 16124
rect 4338 16096 4344 16108
rect 3712 16068 3832 16096
rect 4299 16068 4344 16096
rect 3712 16028 3740 16068
rect 4338 16056 4344 16068
rect 4396 16096 4402 16108
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 4396 16068 5181 16096
rect 4396 16056 4402 16068
rect 5169 16065 5181 16068
rect 5215 16096 5227 16099
rect 5258 16096 5264 16108
rect 5215 16068 5264 16096
rect 5215 16065 5227 16068
rect 5169 16059 5227 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16096 7527 16099
rect 7558 16096 7564 16108
rect 7515 16068 7564 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 8202 16096 8208 16108
rect 8163 16068 8208 16096
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 9401 16099 9459 16105
rect 9401 16065 9413 16099
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 9493 16099 9551 16105
rect 9493 16065 9505 16099
rect 9539 16096 9551 16099
rect 9950 16096 9956 16108
rect 9539 16068 9956 16096
rect 9539 16065 9551 16068
rect 9493 16059 9551 16065
rect 2746 16000 3740 16028
rect 3789 16031 3847 16037
rect 3789 15997 3801 16031
rect 3835 16028 3847 16031
rect 3878 16028 3884 16040
rect 3835 16000 3884 16028
rect 3835 15997 3847 16000
rect 3789 15991 3847 15997
rect 3878 15988 3884 16000
rect 3936 16028 3942 16040
rect 4062 16028 4068 16040
rect 3936 16000 4068 16028
rect 3936 15988 3942 16000
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 4154 15988 4160 16040
rect 4212 16028 4218 16040
rect 4525 16031 4583 16037
rect 4525 16028 4537 16031
rect 4212 16000 4537 16028
rect 4212 15988 4218 16000
rect 4525 15997 4537 16000
rect 4571 15997 4583 16031
rect 4525 15991 4583 15997
rect 4617 16031 4675 16037
rect 4617 15997 4629 16031
rect 4663 16028 4675 16031
rect 5350 16028 5356 16040
rect 4663 16000 5356 16028
rect 4663 15997 4675 16000
rect 4617 15991 4675 15997
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 8386 16028 8392 16040
rect 7116 16000 8392 16028
rect 1578 15960 1584 15972
rect 1539 15932 1584 15960
rect 1578 15920 1584 15932
rect 1636 15920 1642 15972
rect 3544 15963 3602 15969
rect 3544 15929 3556 15963
rect 3590 15960 3602 15963
rect 3694 15960 3700 15972
rect 3590 15932 3700 15960
rect 3590 15929 3602 15932
rect 3544 15923 3602 15929
rect 3694 15920 3700 15932
rect 3752 15920 3758 15972
rect 3970 15920 3976 15972
rect 4028 15960 4034 15972
rect 7116 15960 7144 16000
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 9416 16028 9444 16059
rect 9950 16056 9956 16068
rect 10008 16056 10014 16108
rect 10060 16105 10088 16136
rect 10045 16099 10103 16105
rect 10045 16065 10057 16099
rect 10091 16065 10103 16099
rect 10045 16059 10103 16065
rect 9585 16031 9643 16037
rect 9416 16000 9536 16028
rect 4028 15932 7144 15960
rect 7193 15963 7251 15969
rect 4028 15920 4034 15932
rect 7193 15929 7205 15963
rect 7239 15960 7251 15963
rect 8021 15963 8079 15969
rect 7239 15932 7696 15960
rect 7239 15929 7251 15932
rect 7193 15923 7251 15929
rect 1854 15852 1860 15904
rect 1912 15892 1918 15904
rect 2041 15895 2099 15901
rect 2041 15892 2053 15895
rect 1912 15864 2053 15892
rect 1912 15852 1918 15864
rect 2041 15861 2053 15864
rect 2087 15861 2099 15895
rect 5350 15892 5356 15904
rect 5311 15864 5356 15892
rect 2041 15855 2099 15861
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 5442 15852 5448 15904
rect 5500 15892 5506 15904
rect 6270 15892 6276 15904
rect 5500 15864 5545 15892
rect 6231 15864 6276 15892
rect 5500 15852 5506 15864
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 7282 15892 7288 15904
rect 7243 15864 7288 15892
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 7668 15901 7696 15932
rect 8021 15929 8033 15963
rect 8067 15960 8079 15963
rect 8754 15960 8760 15972
rect 8067 15932 8760 15960
rect 8067 15929 8079 15932
rect 8021 15923 8079 15929
rect 8754 15920 8760 15932
rect 8812 15920 8818 15972
rect 9508 15960 9536 16000
rect 9585 15997 9597 16031
rect 9631 16028 9643 16031
rect 9858 16028 9864 16040
rect 9631 16000 9864 16028
rect 9631 15997 9643 16000
rect 9585 15991 9643 15997
rect 9858 15988 9864 16000
rect 9916 15988 9922 16040
rect 10312 15963 10370 15969
rect 10312 15960 10324 15963
rect 9508 15932 10324 15960
rect 10312 15929 10324 15932
rect 10358 15960 10370 15963
rect 10594 15960 10600 15972
rect 10358 15932 10600 15960
rect 10358 15929 10370 15932
rect 10312 15923 10370 15929
rect 10594 15920 10600 15932
rect 10652 15920 10658 15972
rect 11440 15960 11468 16195
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 14553 16235 14611 16241
rect 14553 16232 14565 16235
rect 13872 16204 14565 16232
rect 13872 16192 13878 16204
rect 14553 16201 14565 16204
rect 14599 16201 14611 16235
rect 14553 16195 14611 16201
rect 16114 16192 16120 16244
rect 16172 16232 16178 16244
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 16172 16204 16773 16232
rect 16172 16192 16178 16204
rect 16761 16201 16773 16204
rect 16807 16232 16819 16235
rect 16942 16232 16948 16244
rect 16807 16204 16948 16232
rect 16807 16201 16819 16204
rect 16761 16195 16819 16201
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 16301 16167 16359 16173
rect 16301 16133 16313 16167
rect 16347 16133 16359 16167
rect 16960 16164 16988 16192
rect 16960 16136 17816 16164
rect 16301 16127 16359 16133
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 14829 16099 14887 16105
rect 14829 16096 14841 16099
rect 14792 16068 14841 16096
rect 14792 16056 14798 16068
rect 14829 16065 14841 16068
rect 14875 16065 14887 16099
rect 16316 16096 16344 16127
rect 16390 16096 16396 16108
rect 16303 16068 16396 16096
rect 14829 16059 14887 16065
rect 16390 16056 16396 16068
rect 16448 16096 16454 16108
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 16448 16068 17049 16096
rect 16448 16056 16454 16068
rect 17037 16065 17049 16068
rect 17083 16065 17095 16099
rect 17037 16059 17095 16065
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16096 17279 16099
rect 17586 16096 17592 16108
rect 17267 16068 17592 16096
rect 17267 16065 17279 16068
rect 17221 16059 17279 16065
rect 11701 16031 11759 16037
rect 11701 15997 11713 16031
rect 11747 16028 11759 16031
rect 13173 16031 13231 16037
rect 13173 16028 13185 16031
rect 11747 16000 13185 16028
rect 11747 15997 11759 16000
rect 11701 15991 11759 15997
rect 13173 15997 13185 16000
rect 13219 16028 13231 16031
rect 13906 16028 13912 16040
rect 13219 16000 13912 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 13906 15988 13912 16000
rect 13964 16028 13970 16040
rect 14921 16031 14979 16037
rect 14921 16028 14933 16031
rect 13964 16000 14933 16028
rect 13964 15988 13970 16000
rect 14921 15997 14933 16000
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 15188 16031 15246 16037
rect 15188 15997 15200 16031
rect 15234 16028 15246 16031
rect 15746 16028 15752 16040
rect 15234 16000 15752 16028
rect 15234 15997 15246 16000
rect 15188 15991 15246 15997
rect 15746 15988 15752 16000
rect 15804 15988 15810 16040
rect 16482 15988 16488 16040
rect 16540 16028 16546 16040
rect 16577 16031 16635 16037
rect 16577 16028 16589 16031
rect 16540 16000 16589 16028
rect 16540 15988 16546 16000
rect 16577 15997 16589 16000
rect 16623 15997 16635 16031
rect 16577 15991 16635 15997
rect 11946 15963 12004 15969
rect 11946 15960 11958 15963
rect 11440 15932 11958 15960
rect 11946 15929 11958 15932
rect 11992 15929 12004 15963
rect 13262 15960 13268 15972
rect 11946 15923 12004 15929
rect 13096 15932 13268 15960
rect 7653 15895 7711 15901
rect 7653 15861 7665 15895
rect 7699 15861 7711 15895
rect 7653 15855 7711 15861
rect 8113 15895 8171 15901
rect 8113 15861 8125 15895
rect 8159 15892 8171 15895
rect 8202 15892 8208 15904
rect 8159 15864 8208 15892
rect 8159 15861 8171 15864
rect 8113 15855 8171 15861
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 13096 15901 13124 15932
rect 13262 15920 13268 15932
rect 13320 15960 13326 15972
rect 13440 15963 13498 15969
rect 13440 15960 13452 15963
rect 13320 15932 13452 15960
rect 13320 15920 13326 15932
rect 13440 15929 13452 15932
rect 13486 15960 13498 15963
rect 15286 15960 15292 15972
rect 13486 15932 15292 15960
rect 13486 15929 13498 15932
rect 13440 15923 13498 15929
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 15470 15920 15476 15972
rect 15528 15960 15534 15972
rect 16393 15963 16451 15969
rect 16393 15960 16405 15963
rect 15528 15932 16405 15960
rect 15528 15920 15534 15932
rect 16393 15929 16405 15932
rect 16439 15960 16451 15963
rect 17236 15960 17264 16059
rect 17586 16056 17592 16068
rect 17644 16056 17650 16108
rect 17788 16105 17816 16136
rect 20346 16124 20352 16176
rect 20404 16164 20410 16176
rect 20625 16167 20683 16173
rect 20625 16164 20637 16167
rect 20404 16136 20637 16164
rect 20404 16124 20410 16136
rect 20625 16133 20637 16136
rect 20671 16164 20683 16167
rect 20671 16136 21312 16164
rect 20671 16133 20683 16136
rect 20625 16127 20683 16133
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16065 17831 16099
rect 17773 16059 17831 16065
rect 17788 16028 17816 16059
rect 20990 16056 20996 16108
rect 21048 16056 21054 16108
rect 21284 16105 21312 16136
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 19245 16031 19303 16037
rect 19245 16028 19257 16031
rect 17788 16000 19257 16028
rect 19245 15997 19257 16000
rect 19291 16028 19303 16031
rect 19334 16028 19340 16040
rect 19291 16000 19340 16028
rect 19291 15997 19303 16000
rect 19245 15991 19303 15997
rect 19334 15988 19340 16000
rect 19392 16028 19398 16040
rect 21008 16028 21036 16056
rect 19392 16000 21036 16028
rect 19392 15988 19398 16000
rect 16439 15932 17264 15960
rect 16439 15929 16451 15932
rect 16393 15923 16451 15929
rect 17494 15920 17500 15972
rect 17552 15960 17558 15972
rect 18018 15963 18076 15969
rect 18018 15960 18030 15963
rect 17552 15932 18030 15960
rect 17552 15920 17558 15932
rect 18018 15929 18030 15932
rect 18064 15929 18076 15963
rect 19490 15963 19548 15969
rect 19490 15960 19502 15963
rect 18018 15923 18076 15929
rect 19168 15932 19502 15960
rect 13081 15895 13139 15901
rect 13081 15861 13093 15895
rect 13127 15861 13139 15895
rect 13081 15855 13139 15861
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 17313 15895 17371 15901
rect 17313 15892 17325 15895
rect 15712 15864 17325 15892
rect 15712 15852 15718 15864
rect 17313 15861 17325 15864
rect 17359 15892 17371 15895
rect 17402 15892 17408 15904
rect 17359 15864 17408 15892
rect 17359 15861 17371 15864
rect 17313 15855 17371 15861
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 17586 15852 17592 15904
rect 17644 15892 17650 15904
rect 19168 15901 19196 15932
rect 19490 15929 19502 15932
rect 19536 15960 19548 15963
rect 19702 15960 19708 15972
rect 19536 15932 19708 15960
rect 19536 15929 19548 15932
rect 19490 15923 19548 15929
rect 19702 15920 19708 15932
rect 19760 15920 19766 15972
rect 20346 15920 20352 15972
rect 20404 15960 20410 15972
rect 21177 15963 21235 15969
rect 21177 15960 21189 15963
rect 20404 15932 21189 15960
rect 20404 15920 20410 15932
rect 21177 15929 21189 15932
rect 21223 15929 21235 15963
rect 21177 15923 21235 15929
rect 17681 15895 17739 15901
rect 17681 15892 17693 15895
rect 17644 15864 17693 15892
rect 17644 15852 17650 15864
rect 17681 15861 17693 15864
rect 17727 15861 17739 15895
rect 17681 15855 17739 15861
rect 19153 15895 19211 15901
rect 19153 15861 19165 15895
rect 19199 15861 19211 15895
rect 21082 15892 21088 15904
rect 21043 15864 21088 15892
rect 19153 15855 19211 15861
rect 21082 15852 21088 15864
rect 21140 15852 21146 15904
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1578 15648 1584 15700
rect 1636 15688 1642 15700
rect 1765 15691 1823 15697
rect 1765 15688 1777 15691
rect 1636 15660 1777 15688
rect 1636 15648 1642 15660
rect 1765 15657 1777 15660
rect 1811 15657 1823 15691
rect 1765 15651 1823 15657
rect 1946 15648 1952 15700
rect 2004 15688 2010 15700
rect 2041 15691 2099 15697
rect 2041 15688 2053 15691
rect 2004 15660 2053 15688
rect 2004 15648 2010 15660
rect 2041 15657 2053 15660
rect 2087 15657 2099 15691
rect 2314 15688 2320 15700
rect 2275 15660 2320 15688
rect 2041 15651 2099 15657
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 2685 15691 2743 15697
rect 2685 15657 2697 15691
rect 2731 15688 2743 15691
rect 3970 15688 3976 15700
rect 2731 15660 3976 15688
rect 2731 15657 2743 15660
rect 2685 15651 2743 15657
rect 2700 15620 2728 15651
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 4338 15648 4344 15700
rect 4396 15688 4402 15700
rect 4709 15691 4767 15697
rect 4709 15688 4721 15691
rect 4396 15660 4721 15688
rect 4396 15648 4402 15660
rect 4709 15657 4721 15660
rect 4755 15657 4767 15691
rect 4709 15651 4767 15657
rect 5169 15691 5227 15697
rect 5169 15657 5181 15691
rect 5215 15688 5227 15691
rect 5442 15688 5448 15700
rect 5215 15660 5448 15688
rect 5215 15657 5227 15660
rect 5169 15651 5227 15657
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 7282 15648 7288 15700
rect 7340 15688 7346 15700
rect 7929 15691 7987 15697
rect 7929 15688 7941 15691
rect 7340 15660 7941 15688
rect 7340 15648 7346 15660
rect 7929 15657 7941 15660
rect 7975 15657 7987 15691
rect 7929 15651 7987 15657
rect 8297 15691 8355 15697
rect 8297 15657 8309 15691
rect 8343 15688 8355 15691
rect 8386 15688 8392 15700
rect 8343 15660 8392 15688
rect 8343 15657 8355 15660
rect 8297 15651 8355 15657
rect 8386 15648 8392 15660
rect 8444 15648 8450 15700
rect 8754 15688 8760 15700
rect 8715 15660 8760 15688
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 8846 15648 8852 15700
rect 8904 15688 8910 15700
rect 11425 15691 11483 15697
rect 8904 15660 11376 15688
rect 8904 15648 8910 15660
rect 1964 15592 2728 15620
rect 4249 15623 4307 15629
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 1964 15561 1992 15592
rect 4249 15589 4261 15623
rect 4295 15620 4307 15623
rect 5537 15623 5595 15629
rect 5537 15620 5549 15623
rect 4295 15592 5549 15620
rect 4295 15589 4307 15592
rect 4249 15583 4307 15589
rect 5537 15589 5549 15592
rect 5583 15589 5595 15623
rect 5537 15583 5595 15589
rect 7561 15623 7619 15629
rect 7561 15589 7573 15623
rect 7607 15620 7619 15623
rect 8202 15620 8208 15632
rect 7607 15592 8208 15620
rect 7607 15589 7619 15592
rect 7561 15583 7619 15589
rect 8202 15580 8208 15592
rect 8260 15620 8266 15632
rect 11348 15620 11376 15660
rect 11425 15657 11437 15691
rect 11471 15688 11483 15691
rect 11885 15691 11943 15697
rect 11885 15688 11897 15691
rect 11471 15660 11897 15688
rect 11471 15657 11483 15660
rect 11425 15651 11483 15657
rect 11885 15657 11897 15660
rect 11931 15657 11943 15691
rect 11885 15651 11943 15657
rect 13725 15691 13783 15697
rect 13725 15657 13737 15691
rect 13771 15688 13783 15691
rect 14737 15691 14795 15697
rect 14737 15688 14749 15691
rect 13771 15660 14749 15688
rect 13771 15657 13783 15660
rect 13725 15651 13783 15657
rect 14737 15657 14749 15660
rect 14783 15657 14795 15691
rect 14737 15651 14795 15657
rect 15580 15660 17448 15688
rect 13538 15620 13544 15632
rect 8260 15592 11284 15620
rect 11348 15592 13544 15620
rect 8260 15580 8266 15592
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15521 1639 15555
rect 1581 15515 1639 15521
rect 1949 15555 2007 15561
rect 1949 15521 1961 15555
rect 1995 15521 2007 15555
rect 1949 15515 2007 15521
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15521 2283 15555
rect 2225 15515 2283 15521
rect 2501 15555 2559 15561
rect 2501 15521 2513 15555
rect 2547 15552 2559 15555
rect 6181 15555 6239 15561
rect 2547 15524 4384 15552
rect 2547 15521 2559 15524
rect 2501 15515 2559 15521
rect 1596 15484 1624 15515
rect 2130 15484 2136 15496
rect 1596 15456 2136 15484
rect 2130 15444 2136 15456
rect 2188 15444 2194 15496
rect 2240 15484 2268 15515
rect 2240 15456 2774 15484
rect 2746 15348 2774 15456
rect 4356 15425 4384 15524
rect 6181 15521 6193 15555
rect 6227 15552 6239 15555
rect 9484 15555 9542 15561
rect 6227 15524 8248 15552
rect 6227 15521 6239 15524
rect 6181 15515 6239 15521
rect 8220 15496 8248 15524
rect 9484 15521 9496 15555
rect 9530 15552 9542 15555
rect 11054 15552 11060 15564
rect 9530 15524 10824 15552
rect 11015 15524 11060 15552
rect 9530 15521 9542 15524
rect 9484 15515 9542 15521
rect 10796 15496 10824 15524
rect 11054 15512 11060 15524
rect 11112 15512 11118 15564
rect 11256 15552 11284 15592
rect 13538 15580 13544 15592
rect 13596 15580 13602 15632
rect 13817 15623 13875 15629
rect 13817 15589 13829 15623
rect 13863 15620 13875 15623
rect 14550 15620 14556 15632
rect 13863 15592 14556 15620
rect 13863 15589 13875 15592
rect 13817 15583 13875 15589
rect 14550 15580 14556 15592
rect 14608 15580 14614 15632
rect 15580 15629 15608 15660
rect 16390 15629 16396 15632
rect 15197 15623 15255 15629
rect 15197 15620 15209 15623
rect 14936 15592 15209 15620
rect 11256 15524 13492 15552
rect 4798 15484 4804 15496
rect 4759 15456 4804 15484
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15484 5043 15487
rect 5534 15484 5540 15496
rect 5031 15456 5540 15484
rect 5031 15453 5043 15456
rect 4985 15447 5043 15453
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 5626 15444 5632 15496
rect 5684 15484 5690 15496
rect 5813 15487 5871 15493
rect 5684 15456 5729 15484
rect 5684 15444 5690 15456
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 5994 15484 6000 15496
rect 5859 15456 6000 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 8202 15444 8208 15496
rect 8260 15444 8266 15496
rect 8386 15484 8392 15496
rect 8347 15456 8392 15484
rect 8386 15444 8392 15456
rect 8444 15444 8450 15496
rect 8481 15487 8539 15493
rect 8481 15453 8493 15487
rect 8527 15453 8539 15487
rect 8481 15447 8539 15453
rect 4341 15419 4399 15425
rect 4341 15385 4353 15419
rect 4387 15385 4399 15419
rect 7282 15416 7288 15428
rect 4341 15379 4399 15385
rect 4448 15388 7288 15416
rect 2869 15351 2927 15357
rect 2869 15348 2881 15351
rect 2746 15320 2881 15348
rect 2869 15317 2881 15320
rect 2915 15348 2927 15351
rect 4448 15348 4476 15388
rect 7282 15376 7288 15388
rect 7340 15376 7346 15428
rect 8294 15376 8300 15428
rect 8352 15416 8358 15428
rect 8496 15416 8524 15447
rect 9122 15444 9128 15496
rect 9180 15484 9186 15496
rect 9217 15487 9275 15493
rect 9217 15484 9229 15487
rect 9180 15456 9229 15484
rect 9180 15444 9186 15456
rect 9217 15453 9229 15456
rect 9263 15453 9275 15487
rect 10778 15484 10784 15496
rect 10739 15456 10784 15484
rect 9217 15447 9275 15453
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 10962 15484 10968 15496
rect 10923 15456 10968 15484
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11974 15484 11980 15496
rect 11935 15456 11980 15484
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 8352 15388 8524 15416
rect 8352 15376 8358 15388
rect 11238 15376 11244 15428
rect 11296 15416 11302 15428
rect 11517 15419 11575 15425
rect 11517 15416 11529 15419
rect 11296 15388 11529 15416
rect 11296 15376 11302 15388
rect 11517 15385 11529 15388
rect 11563 15385 11575 15419
rect 11517 15379 11575 15385
rect 2915 15320 4476 15348
rect 2915 15317 2927 15320
rect 2869 15311 2927 15317
rect 5902 15308 5908 15360
rect 5960 15348 5966 15360
rect 5997 15351 6055 15357
rect 5997 15348 6009 15351
rect 5960 15320 6009 15348
rect 5960 15308 5966 15320
rect 5997 15317 6009 15320
rect 6043 15348 6055 15351
rect 6178 15348 6184 15360
rect 6043 15320 6184 15348
rect 6043 15317 6055 15320
rect 5997 15311 6055 15317
rect 6178 15308 6184 15320
rect 6236 15308 6242 15360
rect 8478 15308 8484 15360
rect 8536 15348 8542 15360
rect 8846 15348 8852 15360
rect 8536 15320 8852 15348
rect 8536 15308 8542 15320
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 10594 15348 10600 15360
rect 10507 15320 10600 15348
rect 10594 15308 10600 15320
rect 10652 15348 10658 15360
rect 12084 15348 12112 15447
rect 10652 15320 12112 15348
rect 13464 15348 13492 15524
rect 13633 15487 13691 15493
rect 13633 15453 13645 15487
rect 13679 15484 13691 15487
rect 13814 15484 13820 15496
rect 13679 15456 13820 15484
rect 13679 15453 13691 15456
rect 13633 15447 13691 15453
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 14936 15484 14964 15592
rect 15197 15589 15209 15592
rect 15243 15620 15255 15623
rect 15565 15623 15623 15629
rect 15565 15620 15577 15623
rect 15243 15592 15577 15620
rect 15243 15589 15255 15592
rect 15197 15583 15255 15589
rect 15565 15589 15577 15592
rect 15611 15589 15623 15623
rect 16384 15620 16396 15629
rect 16351 15592 16396 15620
rect 15565 15583 15623 15589
rect 16384 15583 16396 15592
rect 16390 15580 16396 15583
rect 16448 15580 16454 15632
rect 17420 15620 17448 15660
rect 17494 15648 17500 15700
rect 17552 15688 17558 15700
rect 17589 15691 17647 15697
rect 17589 15688 17601 15691
rect 17552 15660 17601 15688
rect 17552 15648 17558 15660
rect 17589 15657 17601 15660
rect 17635 15657 17647 15691
rect 19610 15688 19616 15700
rect 17589 15651 17647 15657
rect 17696 15660 19616 15688
rect 17696 15620 17724 15660
rect 19610 15648 19616 15660
rect 19668 15648 19674 15700
rect 19886 15688 19892 15700
rect 19847 15660 19892 15688
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20346 15688 20352 15700
rect 20307 15660 20352 15688
rect 20346 15648 20352 15660
rect 20404 15648 20410 15700
rect 20717 15691 20775 15697
rect 20717 15657 20729 15691
rect 20763 15688 20775 15691
rect 20898 15688 20904 15700
rect 20763 15660 20904 15688
rect 20763 15657 20775 15660
rect 20717 15651 20775 15657
rect 20898 15648 20904 15660
rect 20956 15648 20962 15700
rect 20993 15691 21051 15697
rect 20993 15657 21005 15691
rect 21039 15657 21051 15691
rect 20993 15651 21051 15657
rect 21008 15620 21036 15651
rect 21361 15623 21419 15629
rect 21361 15620 21373 15623
rect 17420 15592 17724 15620
rect 17880 15592 20944 15620
rect 21008 15592 21373 15620
rect 15105 15555 15163 15561
rect 15105 15521 15117 15555
rect 15151 15552 15163 15555
rect 17880 15552 17908 15592
rect 18702 15555 18760 15561
rect 18702 15552 18714 15555
rect 15151 15524 17908 15552
rect 17972 15524 18714 15552
rect 15151 15521 15163 15524
rect 15105 15515 15163 15521
rect 15286 15484 15292 15496
rect 14108 15456 14964 15484
rect 15247 15456 15292 15484
rect 13538 15376 13544 15428
rect 13596 15416 13602 15428
rect 14108 15416 14136 15456
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 16114 15484 16120 15496
rect 16075 15456 16120 15484
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 17972 15428 18000 15524
rect 18702 15521 18714 15524
rect 18748 15521 18760 15555
rect 18702 15515 18760 15521
rect 18969 15555 19027 15561
rect 18969 15521 18981 15555
rect 19015 15552 19027 15555
rect 19334 15552 19340 15564
rect 19015 15524 19340 15552
rect 19015 15521 19027 15524
rect 18969 15515 19027 15521
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 19426 15512 19432 15564
rect 19484 15552 19490 15564
rect 19981 15555 20039 15561
rect 19981 15552 19993 15555
rect 19484 15524 19993 15552
rect 19484 15512 19490 15524
rect 19981 15521 19993 15524
rect 20027 15552 20039 15555
rect 20346 15552 20352 15564
rect 20027 15524 20352 15552
rect 20027 15521 20039 15524
rect 19981 15515 20039 15521
rect 20346 15512 20352 15524
rect 20404 15512 20410 15564
rect 20533 15555 20591 15561
rect 20533 15521 20545 15555
rect 20579 15521 20591 15555
rect 20533 15515 20591 15521
rect 19058 15444 19064 15496
rect 19116 15484 19122 15496
rect 19702 15484 19708 15496
rect 19116 15456 19161 15484
rect 19663 15456 19708 15484
rect 19116 15444 19122 15456
rect 19702 15444 19708 15456
rect 19760 15444 19766 15496
rect 13596 15388 14136 15416
rect 14185 15419 14243 15425
rect 13596 15376 13602 15388
rect 14185 15385 14197 15419
rect 14231 15416 14243 15419
rect 15378 15416 15384 15428
rect 14231 15388 15384 15416
rect 14231 15385 14243 15388
rect 14185 15379 14243 15385
rect 15378 15376 15384 15388
rect 15436 15376 15442 15428
rect 17497 15419 17555 15425
rect 17497 15385 17509 15419
rect 17543 15416 17555 15419
rect 17954 15416 17960 15428
rect 17543 15388 17960 15416
rect 17543 15385 17555 15388
rect 17497 15379 17555 15385
rect 17954 15376 17960 15388
rect 18012 15376 18018 15428
rect 20548 15416 20576 15515
rect 20622 15512 20628 15564
rect 20680 15552 20686 15564
rect 20809 15555 20867 15561
rect 20809 15552 20821 15555
rect 20680 15524 20821 15552
rect 20680 15512 20686 15524
rect 20809 15521 20821 15524
rect 20855 15521 20867 15555
rect 20809 15515 20867 15521
rect 20916 15484 20944 15592
rect 21361 15589 21373 15592
rect 21407 15589 21419 15623
rect 21361 15583 21419 15589
rect 21542 15552 21548 15564
rect 21503 15524 21548 15552
rect 21542 15512 21548 15524
rect 21600 15512 21606 15564
rect 21450 15484 21456 15496
rect 20916 15456 21456 15484
rect 21450 15444 21456 15456
rect 21508 15444 21514 15496
rect 21085 15419 21143 15425
rect 21085 15416 21097 15419
rect 19306 15388 21097 15416
rect 14458 15348 14464 15360
rect 13464 15320 14464 15348
rect 10652 15308 10658 15320
rect 14458 15308 14464 15320
rect 14516 15348 14522 15360
rect 19306 15348 19334 15388
rect 21085 15385 21097 15388
rect 21131 15385 21143 15419
rect 21085 15379 21143 15385
rect 19426 15348 19432 15360
rect 14516 15320 19334 15348
rect 19387 15320 19432 15348
rect 14516 15308 14522 15320
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 19610 15308 19616 15360
rect 19668 15348 19674 15360
rect 21818 15348 21824 15360
rect 19668 15320 21824 15348
rect 19668 15308 19674 15320
rect 21818 15308 21824 15320
rect 21876 15308 21882 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 1486 15144 1492 15156
rect 1447 15116 1492 15144
rect 1486 15104 1492 15116
rect 1544 15104 1550 15156
rect 3697 15147 3755 15153
rect 3697 15113 3709 15147
rect 3743 15144 3755 15147
rect 5350 15144 5356 15156
rect 3743 15116 5356 15144
rect 3743 15113 3755 15116
rect 3697 15107 3755 15113
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 5534 15104 5540 15156
rect 5592 15144 5598 15156
rect 5629 15147 5687 15153
rect 5629 15144 5641 15147
rect 5592 15116 5641 15144
rect 5592 15104 5598 15116
rect 5629 15113 5641 15116
rect 5675 15113 5687 15147
rect 5629 15107 5687 15113
rect 6914 15104 6920 15156
rect 6972 15144 6978 15156
rect 7469 15147 7527 15153
rect 7469 15144 7481 15147
rect 6972 15116 7481 15144
rect 6972 15104 6978 15116
rect 7469 15113 7481 15116
rect 7515 15113 7527 15147
rect 8294 15144 8300 15156
rect 8207 15116 8300 15144
rect 7469 15107 7527 15113
rect 8294 15104 8300 15116
rect 8352 15144 8358 15156
rect 9214 15144 9220 15156
rect 8352 15116 9220 15144
rect 8352 15104 8358 15116
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 11517 15147 11575 15153
rect 11517 15113 11529 15147
rect 11563 15144 11575 15147
rect 11974 15144 11980 15156
rect 11563 15116 11980 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 11974 15104 11980 15116
rect 12032 15104 12038 15156
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 15654 15144 15660 15156
rect 12308 15116 15660 15144
rect 12308 15104 12314 15116
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 15749 15147 15807 15153
rect 15749 15113 15761 15147
rect 15795 15144 15807 15147
rect 16482 15144 16488 15156
rect 15795 15116 16488 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 17129 15147 17187 15153
rect 17129 15113 17141 15147
rect 17175 15144 17187 15147
rect 17310 15144 17316 15156
rect 17175 15116 17316 15144
rect 17175 15113 17187 15116
rect 17129 15107 17187 15113
rect 17310 15104 17316 15116
rect 17368 15104 17374 15156
rect 17957 15147 18015 15153
rect 17957 15113 17969 15147
rect 18003 15144 18015 15147
rect 18046 15144 18052 15156
rect 18003 15116 18052 15144
rect 18003 15113 18015 15116
rect 17957 15107 18015 15113
rect 18046 15104 18052 15116
rect 18104 15104 18110 15156
rect 19337 15147 19395 15153
rect 19337 15113 19349 15147
rect 19383 15144 19395 15147
rect 19886 15144 19892 15156
rect 19383 15116 19892 15144
rect 19383 15113 19395 15116
rect 19337 15107 19395 15113
rect 19886 15104 19892 15116
rect 19944 15104 19950 15156
rect 20533 15147 20591 15153
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 21358 15144 21364 15156
rect 20579 15116 21364 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 21358 15104 21364 15116
rect 21416 15104 21422 15156
rect 9950 15076 9956 15088
rect 6012 15048 9956 15076
rect 2866 14968 2872 15020
rect 2924 15008 2930 15020
rect 3053 15011 3111 15017
rect 3053 15008 3065 15011
rect 2924 14980 3065 15008
rect 2924 14968 2930 14980
rect 3053 14977 3065 14980
rect 3099 14977 3111 15011
rect 3053 14971 3111 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 1995 14912 2176 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2148 14881 2176 14912
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4249 14943 4307 14949
rect 4249 14940 4261 14943
rect 4120 14912 4261 14940
rect 4120 14900 4126 14912
rect 4249 14909 4261 14912
rect 4295 14940 4307 14943
rect 5902 14940 5908 14952
rect 4295 14912 5908 14940
rect 4295 14909 4307 14912
rect 4249 14903 4307 14909
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 1581 14875 1639 14881
rect 1581 14841 1593 14875
rect 1627 14872 1639 14875
rect 2133 14875 2191 14881
rect 1627 14844 1808 14872
rect 1627 14841 1639 14844
rect 1581 14835 1639 14841
rect 1780 14813 1808 14844
rect 2133 14841 2145 14875
rect 2179 14872 2191 14875
rect 3237 14875 3295 14881
rect 3237 14872 3249 14875
rect 2179 14844 3249 14872
rect 2179 14841 2191 14844
rect 2133 14835 2191 14841
rect 3237 14841 3249 14844
rect 3283 14872 3295 14875
rect 3283 14844 3832 14872
rect 3283 14841 3295 14844
rect 3237 14835 3295 14841
rect 1765 14807 1823 14813
rect 1765 14773 1777 14807
rect 1811 14773 1823 14807
rect 1765 14767 1823 14773
rect 3326 14764 3332 14816
rect 3384 14804 3390 14816
rect 3804 14813 3832 14844
rect 3878 14832 3884 14884
rect 3936 14872 3942 14884
rect 4494 14875 4552 14881
rect 4494 14872 4506 14875
rect 3936 14844 4506 14872
rect 3936 14832 3942 14844
rect 4494 14841 4506 14844
rect 4540 14841 4552 14875
rect 6012 14872 6040 15048
rect 9950 15036 9956 15048
rect 10008 15036 10014 15088
rect 10689 15079 10747 15085
rect 10689 15045 10701 15079
rect 10735 15076 10747 15079
rect 15378 15076 15384 15088
rect 10735 15048 15384 15076
rect 10735 15045 10747 15048
rect 10689 15039 10747 15045
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 15473 15079 15531 15085
rect 15473 15045 15485 15079
rect 15519 15076 15531 15079
rect 19981 15079 20039 15085
rect 15519 15048 19840 15076
rect 15519 15045 15531 15048
rect 15473 15039 15531 15045
rect 6822 14968 6828 15020
rect 6880 15008 6886 15020
rect 7009 15011 7067 15017
rect 7009 15008 7021 15011
rect 6880 14980 7021 15008
rect 6880 14968 6886 14980
rect 7009 14977 7021 14980
rect 7055 14977 7067 15011
rect 7009 14971 7067 14977
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 15008 8079 15011
rect 8294 15008 8300 15020
rect 8067 14980 8300 15008
rect 8067 14977 8079 14980
rect 8021 14971 8079 14977
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 8846 14968 8852 15020
rect 8904 15008 8910 15020
rect 8941 15011 8999 15017
rect 8941 15008 8953 15011
rect 8904 14980 8953 15008
rect 8904 14968 8910 14980
rect 8941 14977 8953 14980
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 10778 14968 10784 15020
rect 10836 15008 10842 15020
rect 10873 15011 10931 15017
rect 10873 15008 10885 15011
rect 10836 14980 10885 15008
rect 10836 14968 10842 14980
rect 10873 14977 10885 14980
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11112 14980 11713 15008
rect 11112 14968 11118 14980
rect 11701 14977 11713 14980
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12345 15011 12403 15017
rect 12032 14980 12296 15008
rect 12032 14968 12038 14980
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14940 6975 14943
rect 7190 14940 7196 14952
rect 6963 14912 7196 14940
rect 6963 14909 6975 14912
rect 6917 14903 6975 14909
rect 7190 14900 7196 14912
rect 7248 14940 7254 14952
rect 8202 14940 8208 14952
rect 7248 14912 8208 14940
rect 7248 14900 7254 14912
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8489 14943 8547 14949
rect 8489 14909 8501 14943
rect 8535 14940 8547 14943
rect 8662 14940 8668 14952
rect 8535 14912 8668 14940
rect 8535 14909 8547 14912
rect 8489 14903 8547 14909
rect 8662 14900 8668 14912
rect 8720 14900 8726 14952
rect 9766 14900 9772 14952
rect 9824 14940 9830 14952
rect 11149 14943 11207 14949
rect 9824 14912 10824 14940
rect 9824 14900 9830 14912
rect 4494 14835 4552 14841
rect 5000 14844 6040 14872
rect 6288 14844 8340 14872
rect 3789 14807 3847 14813
rect 3384 14776 3429 14804
rect 3384 14764 3390 14776
rect 3789 14773 3801 14807
rect 3835 14804 3847 14807
rect 5000 14804 5028 14844
rect 3835 14776 5028 14804
rect 3835 14773 3847 14776
rect 3789 14767 3847 14773
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 5813 14807 5871 14813
rect 5813 14804 5825 14807
rect 5684 14776 5825 14804
rect 5684 14764 5690 14776
rect 5813 14773 5825 14776
rect 5859 14804 5871 14807
rect 5994 14804 6000 14816
rect 5859 14776 6000 14804
rect 5859 14773 5871 14776
rect 5813 14767 5871 14773
rect 5994 14764 6000 14776
rect 6052 14804 6058 14816
rect 6288 14804 6316 14844
rect 6454 14804 6460 14816
rect 6052 14776 6316 14804
rect 6415 14776 6460 14804
rect 6052 14764 6058 14776
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 6825 14807 6883 14813
rect 6825 14773 6837 14807
rect 6871 14804 6883 14807
rect 7650 14804 7656 14816
rect 6871 14776 7656 14804
rect 6871 14773 6883 14776
rect 6825 14767 6883 14773
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 7742 14764 7748 14816
rect 7800 14804 7806 14816
rect 7837 14807 7895 14813
rect 7837 14804 7849 14807
rect 7800 14776 7849 14804
rect 7800 14764 7806 14776
rect 7837 14773 7849 14776
rect 7883 14773 7895 14807
rect 7837 14767 7895 14773
rect 7929 14807 7987 14813
rect 7929 14773 7941 14807
rect 7975 14804 7987 14807
rect 8202 14804 8208 14816
rect 7975 14776 8208 14804
rect 7975 14773 7987 14776
rect 7929 14767 7987 14773
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 8312 14804 8340 14844
rect 8386 14832 8392 14884
rect 8444 14872 8450 14884
rect 8849 14875 8907 14881
rect 8849 14872 8861 14875
rect 8444 14844 8861 14872
rect 8444 14832 8450 14844
rect 8849 14841 8861 14844
rect 8895 14872 8907 14875
rect 9398 14872 9404 14884
rect 8895 14844 9404 14872
rect 8895 14841 8907 14844
rect 8849 14835 8907 14841
rect 9398 14832 9404 14844
rect 9456 14832 9462 14884
rect 10689 14875 10747 14881
rect 10689 14872 10701 14875
rect 9646 14844 10701 14872
rect 9646 14804 9674 14844
rect 10689 14841 10701 14844
rect 10735 14841 10747 14875
rect 10796 14872 10824 14912
rect 11149 14909 11161 14943
rect 11195 14940 11207 14943
rect 12158 14940 12164 14952
rect 11195 14912 12164 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 12158 14900 12164 14912
rect 12216 14900 12222 14952
rect 12268 14940 12296 14980
rect 12345 14977 12357 15011
rect 12391 15008 12403 15011
rect 12802 15008 12808 15020
rect 12391 14980 12808 15008
rect 12391 14977 12403 14980
rect 12345 14971 12403 14977
rect 12802 14968 12808 14980
rect 12860 14968 12866 15020
rect 13173 15011 13231 15017
rect 13173 14977 13185 15011
rect 13219 15008 13231 15011
rect 13998 15008 14004 15020
rect 13219 14980 14004 15008
rect 13219 14977 13231 14980
rect 13173 14971 13231 14977
rect 13998 14968 14004 14980
rect 14056 14968 14062 15020
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 15008 14979 15011
rect 15746 15008 15752 15020
rect 14967 14980 15752 15008
rect 14967 14977 14979 14980
rect 14921 14971 14979 14977
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 17586 15008 17592 15020
rect 17547 14980 17592 15008
rect 17586 14968 17592 14980
rect 17644 14968 17650 15020
rect 17773 15011 17831 15017
rect 17773 14977 17785 15011
rect 17819 15008 17831 15011
rect 17954 15008 17960 15020
rect 17819 14980 17960 15008
rect 17819 14977 17831 14980
rect 17773 14971 17831 14977
rect 17954 14968 17960 14980
rect 18012 15008 18018 15020
rect 18509 15011 18567 15017
rect 18509 15008 18521 15011
rect 18012 14980 18521 15008
rect 18012 14968 18018 14980
rect 18509 14977 18521 14980
rect 18555 14977 18567 15011
rect 18509 14971 18567 14977
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12268 14912 12449 14940
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 14550 14900 14556 14952
rect 14608 14940 14614 14952
rect 15565 14943 15623 14949
rect 15565 14940 15577 14943
rect 14608 14912 15577 14940
rect 14608 14900 14614 14912
rect 15565 14909 15577 14912
rect 15611 14909 15623 14943
rect 15565 14903 15623 14909
rect 18325 14943 18383 14949
rect 18325 14909 18337 14943
rect 18371 14940 18383 14943
rect 19058 14940 19064 14952
rect 18371 14912 19064 14940
rect 18371 14909 18383 14912
rect 18325 14903 18383 14909
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 19613 14943 19671 14949
rect 19613 14940 19625 14943
rect 19168 14912 19625 14940
rect 10870 14872 10876 14884
rect 10783 14844 10876 14872
rect 10689 14835 10747 14841
rect 10870 14832 10876 14844
rect 10928 14872 10934 14884
rect 12529 14875 12587 14881
rect 12529 14872 12541 14875
rect 10928 14844 12541 14872
rect 10928 14832 10934 14844
rect 12529 14841 12541 14844
rect 12575 14841 12587 14875
rect 12529 14835 12587 14841
rect 14734 14832 14740 14884
rect 14792 14872 14798 14884
rect 15105 14875 15163 14881
rect 15105 14872 15117 14875
rect 14792 14844 15117 14872
rect 14792 14832 14798 14844
rect 15105 14841 15117 14844
rect 15151 14841 15163 14875
rect 15105 14835 15163 14841
rect 15378 14832 15384 14884
rect 15436 14872 15442 14884
rect 19168 14872 19196 14912
rect 19613 14909 19625 14912
rect 19659 14940 19671 14943
rect 19702 14940 19708 14952
rect 19659 14912 19708 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 19702 14900 19708 14912
rect 19760 14900 19766 14952
rect 19812 14949 19840 15048
rect 19981 15045 19993 15079
rect 20027 15045 20039 15079
rect 19981 15039 20039 15045
rect 20257 15079 20315 15085
rect 20257 15045 20269 15079
rect 20303 15076 20315 15079
rect 20806 15076 20812 15088
rect 20303 15048 20812 15076
rect 20303 15045 20315 15048
rect 20257 15039 20315 15045
rect 19797 14943 19855 14949
rect 19797 14909 19809 14943
rect 19843 14909 19855 14943
rect 19996 14940 20024 15039
rect 20806 15036 20812 15048
rect 20864 15036 20870 15088
rect 21174 15076 21180 15088
rect 21135 15048 21180 15076
rect 21174 15036 21180 15048
rect 21232 15036 21238 15088
rect 20073 14943 20131 14949
rect 20073 14940 20085 14943
rect 19996 14912 20085 14940
rect 19797 14903 19855 14909
rect 20073 14909 20085 14912
rect 20119 14909 20131 14943
rect 20073 14903 20131 14909
rect 20349 14943 20407 14949
rect 20349 14909 20361 14943
rect 20395 14909 20407 14943
rect 20349 14903 20407 14909
rect 20625 14943 20683 14949
rect 20625 14909 20637 14943
rect 20671 14909 20683 14943
rect 20625 14903 20683 14909
rect 20364 14872 20392 14903
rect 15436 14844 19196 14872
rect 19444 14844 20392 14872
rect 15436 14832 15442 14844
rect 10594 14804 10600 14816
rect 8312 14776 9674 14804
rect 10555 14776 10600 14804
rect 10594 14764 10600 14776
rect 10652 14804 10658 14816
rect 10962 14804 10968 14816
rect 10652 14776 10968 14804
rect 10652 14764 10658 14776
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11057 14807 11115 14813
rect 11057 14773 11069 14807
rect 11103 14804 11115 14807
rect 11698 14804 11704 14816
rect 11103 14776 11704 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 11698 14764 11704 14776
rect 11756 14804 11762 14816
rect 11977 14807 12035 14813
rect 11977 14804 11989 14807
rect 11756 14776 11989 14804
rect 11756 14764 11762 14776
rect 11977 14773 11989 14776
rect 12023 14773 12035 14807
rect 11977 14767 12035 14773
rect 12897 14807 12955 14813
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 13265 14807 13323 14813
rect 13265 14804 13277 14807
rect 12943 14776 13277 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 13265 14773 13277 14776
rect 13311 14773 13323 14807
rect 13265 14767 13323 14773
rect 13357 14807 13415 14813
rect 13357 14773 13369 14807
rect 13403 14804 13415 14807
rect 13538 14804 13544 14816
rect 13403 14776 13544 14804
rect 13403 14773 13415 14776
rect 13357 14767 13415 14773
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 13725 14807 13783 14813
rect 13725 14773 13737 14807
rect 13771 14804 13783 14807
rect 15013 14807 15071 14813
rect 15013 14804 15025 14807
rect 13771 14776 15025 14804
rect 13771 14773 13783 14776
rect 13725 14767 13783 14773
rect 15013 14773 15025 14776
rect 15059 14773 15071 14807
rect 15013 14767 15071 14773
rect 15654 14764 15660 14816
rect 15712 14804 15718 14816
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15712 14776 15853 14804
rect 15712 14764 15718 14776
rect 15841 14773 15853 14776
rect 15887 14804 15899 14807
rect 16298 14804 16304 14816
rect 15887 14776 16304 14804
rect 15887 14773 15899 14776
rect 15841 14767 15899 14773
rect 16298 14764 16304 14776
rect 16356 14804 16362 14816
rect 17218 14804 17224 14816
rect 16356 14776 17224 14804
rect 16356 14764 16362 14776
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 17494 14804 17500 14816
rect 17455 14776 17500 14804
rect 17494 14764 17500 14776
rect 17552 14764 17558 14816
rect 18138 14764 18144 14816
rect 18196 14804 18202 14816
rect 18417 14807 18475 14813
rect 18417 14804 18429 14807
rect 18196 14776 18429 14804
rect 18196 14764 18202 14776
rect 18417 14773 18429 14776
rect 18463 14804 18475 14807
rect 18966 14804 18972 14816
rect 18463 14776 18972 14804
rect 18463 14773 18475 14776
rect 18417 14767 18475 14773
rect 18966 14764 18972 14776
rect 19024 14764 19030 14816
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 19444 14813 19472 14844
rect 19429 14807 19487 14813
rect 19429 14804 19441 14807
rect 19392 14776 19441 14804
rect 19392 14764 19398 14776
rect 19429 14773 19441 14776
rect 19475 14773 19487 14807
rect 19429 14767 19487 14773
rect 19702 14764 19708 14816
rect 19760 14804 19766 14816
rect 19886 14804 19892 14816
rect 19760 14776 19892 14804
rect 19760 14764 19766 14776
rect 19886 14764 19892 14776
rect 19944 14804 19950 14816
rect 20640 14804 20668 14903
rect 20993 14875 21051 14881
rect 20993 14841 21005 14875
rect 21039 14841 21051 14875
rect 21358 14872 21364 14884
rect 21319 14844 21364 14872
rect 20993 14835 21051 14841
rect 19944 14776 20668 14804
rect 20809 14807 20867 14813
rect 19944 14764 19950 14776
rect 20809 14773 20821 14807
rect 20855 14804 20867 14807
rect 21008 14804 21036 14835
rect 21358 14832 21364 14844
rect 21416 14832 21422 14884
rect 21542 14872 21548 14884
rect 21503 14844 21548 14872
rect 21542 14832 21548 14844
rect 21600 14832 21606 14884
rect 20855 14776 21036 14804
rect 20855 14773 20867 14776
rect 20809 14767 20867 14773
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 2130 14600 2136 14612
rect 2091 14572 2136 14600
rect 2130 14560 2136 14572
rect 2188 14560 2194 14612
rect 3602 14560 3608 14612
rect 3660 14600 3666 14612
rect 14274 14600 14280 14612
rect 3660 14572 14280 14600
rect 3660 14560 3666 14572
rect 14274 14560 14280 14572
rect 14332 14600 14338 14612
rect 15746 14600 15752 14612
rect 14332 14572 15608 14600
rect 15707 14572 15752 14600
rect 14332 14560 14338 14572
rect 5534 14492 5540 14544
rect 5592 14532 5598 14544
rect 5782 14535 5840 14541
rect 5782 14532 5794 14535
rect 5592 14504 5794 14532
rect 5592 14492 5598 14504
rect 5782 14501 5794 14504
rect 5828 14501 5840 14535
rect 5782 14495 5840 14501
rect 6546 14492 6552 14544
rect 6604 14532 6610 14544
rect 6730 14532 6736 14544
rect 6604 14504 6736 14532
rect 6604 14492 6610 14504
rect 6730 14492 6736 14504
rect 6788 14492 6794 14544
rect 7466 14492 7472 14544
rect 7524 14532 7530 14544
rect 9401 14535 9459 14541
rect 9401 14532 9413 14535
rect 7524 14504 9413 14532
rect 7524 14492 7530 14504
rect 9401 14501 9413 14504
rect 9447 14501 9459 14535
rect 9401 14495 9459 14501
rect 9493 14535 9551 14541
rect 9493 14501 9505 14535
rect 9539 14532 9551 14535
rect 9766 14532 9772 14544
rect 9539 14504 9772 14532
rect 9539 14501 9551 14504
rect 9493 14495 9551 14501
rect 1578 14464 1584 14476
rect 1539 14436 1584 14464
rect 1578 14424 1584 14436
rect 1636 14424 1642 14476
rect 2041 14467 2099 14473
rect 2041 14433 2053 14467
rect 2087 14464 2099 14467
rect 2130 14464 2136 14476
rect 2087 14436 2136 14464
rect 2087 14433 2099 14436
rect 2041 14427 2099 14433
rect 2130 14424 2136 14436
rect 2188 14424 2194 14476
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14464 2375 14467
rect 2590 14464 2596 14476
rect 2363 14436 2452 14464
rect 2551 14436 2596 14464
rect 2363 14433 2375 14436
rect 2317 14427 2375 14433
rect 2424 14337 2452 14436
rect 2590 14424 2596 14436
rect 2648 14424 2654 14476
rect 4982 14464 4988 14476
rect 5040 14473 5046 14476
rect 5040 14467 5063 14473
rect 4915 14436 4988 14464
rect 4982 14424 4988 14436
rect 5051 14464 5063 14467
rect 6822 14464 6828 14476
rect 5051 14436 6828 14464
rect 5051 14433 5063 14436
rect 5040 14427 5063 14433
rect 5040 14424 5046 14427
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 6914 14424 6920 14476
rect 6972 14464 6978 14476
rect 7552 14467 7610 14473
rect 7552 14464 7564 14467
rect 6972 14436 7564 14464
rect 6972 14424 6978 14436
rect 7552 14433 7564 14436
rect 7598 14464 7610 14467
rect 9416 14464 9444 14495
rect 9766 14492 9772 14504
rect 9824 14532 9830 14544
rect 11146 14532 11152 14544
rect 9824 14504 11152 14532
rect 9824 14492 9830 14504
rect 11146 14492 11152 14504
rect 11204 14492 11210 14544
rect 12802 14492 12808 14544
rect 12860 14541 12866 14544
rect 12860 14535 12924 14541
rect 12860 14501 12878 14535
rect 12912 14532 12924 14535
rect 12912 14504 13952 14532
rect 12912 14501 12924 14504
rect 12860 14495 12924 14501
rect 12860 14492 12866 14495
rect 10962 14464 10968 14476
rect 7598 14436 9260 14464
rect 9416 14436 10968 14464
rect 7598 14433 7610 14436
rect 7552 14427 7610 14433
rect 9232 14408 9260 14436
rect 10962 14424 10968 14436
rect 11020 14424 11026 14476
rect 12621 14467 12679 14473
rect 12621 14433 12633 14467
rect 12667 14464 12679 14467
rect 13924 14464 13952 14504
rect 13998 14492 14004 14544
rect 14056 14532 14062 14544
rect 14614 14535 14672 14541
rect 14614 14532 14626 14535
rect 14056 14504 14626 14532
rect 14056 14492 14062 14504
rect 14614 14501 14626 14504
rect 14660 14532 14672 14535
rect 15470 14532 15476 14544
rect 14660 14504 15476 14532
rect 14660 14501 14672 14504
rect 14614 14495 14672 14501
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 15580 14532 15608 14572
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 16298 14600 16304 14612
rect 16259 14572 16304 14600
rect 16298 14560 16304 14572
rect 16356 14560 16362 14612
rect 16666 14560 16672 14612
rect 16724 14600 16730 14612
rect 19334 14600 19340 14612
rect 16724 14572 19340 14600
rect 16724 14560 16730 14572
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 19429 14603 19487 14609
rect 19429 14569 19441 14603
rect 19475 14600 19487 14603
rect 20622 14600 20628 14612
rect 19475 14572 20628 14600
rect 19475 14569 19487 14572
rect 19429 14563 19487 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 20809 14603 20867 14609
rect 20809 14569 20821 14603
rect 20855 14600 20867 14603
rect 21266 14600 21272 14612
rect 20855 14572 21272 14600
rect 20855 14569 20867 14572
rect 20809 14563 20867 14569
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 15580 14504 17448 14532
rect 16209 14467 16267 14473
rect 12667 14436 13768 14464
rect 13924 14436 16160 14464
rect 12667 14433 12679 14436
rect 12621 14427 12679 14433
rect 5261 14399 5319 14405
rect 5261 14365 5273 14399
rect 5307 14396 5319 14399
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 5307 14368 5549 14396
rect 5307 14365 5319 14368
rect 5261 14359 5319 14365
rect 5537 14365 5549 14368
rect 5583 14365 5595 14399
rect 7285 14399 7343 14405
rect 7285 14396 7297 14399
rect 5537 14359 5595 14365
rect 6564 14368 7297 14396
rect 2409 14331 2467 14337
rect 2409 14297 2421 14331
rect 2455 14297 2467 14331
rect 2409 14291 2467 14297
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 3878 14260 3884 14272
rect 3839 14232 3884 14260
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 5552 14260 5580 14359
rect 5902 14260 5908 14272
rect 5552 14232 5908 14260
rect 5902 14220 5908 14232
rect 5960 14260 5966 14272
rect 6564 14260 6592 14368
rect 7285 14365 7297 14368
rect 7331 14365 7343 14399
rect 7285 14359 7343 14365
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 8662 14396 8668 14408
rect 8536 14368 8668 14396
rect 8536 14356 8542 14368
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 9214 14396 9220 14408
rect 9175 14368 9220 14396
rect 9214 14356 9220 14368
rect 9272 14356 9278 14408
rect 13740 14396 13768 14436
rect 13906 14396 13912 14408
rect 13740 14368 13912 14396
rect 13906 14356 13912 14368
rect 13964 14396 13970 14408
rect 14369 14399 14427 14405
rect 14369 14396 14381 14399
rect 13964 14368 14381 14396
rect 13964 14356 13970 14368
rect 14369 14365 14381 14368
rect 14415 14365 14427 14399
rect 16132 14396 16160 14436
rect 16209 14433 16221 14467
rect 16255 14464 16267 14467
rect 16574 14464 16580 14476
rect 16255 14436 16580 14464
rect 16255 14433 16267 14436
rect 16209 14427 16267 14433
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 17420 14464 17448 14504
rect 17494 14492 17500 14544
rect 17552 14532 17558 14544
rect 19702 14532 19708 14544
rect 17552 14504 19708 14532
rect 17552 14492 17558 14504
rect 19702 14492 19708 14504
rect 19760 14492 19766 14544
rect 19978 14532 19984 14544
rect 19904 14504 19984 14532
rect 19245 14467 19303 14473
rect 17420 14436 19104 14464
rect 16298 14396 16304 14408
rect 16132 14368 16304 14396
rect 14369 14359 14427 14365
rect 16298 14356 16304 14368
rect 16356 14396 16362 14408
rect 16393 14399 16451 14405
rect 16393 14396 16405 14399
rect 16356 14368 16405 14396
rect 16356 14356 16362 14368
rect 16393 14365 16405 14368
rect 16439 14365 16451 14399
rect 19076 14396 19104 14436
rect 19245 14433 19257 14467
rect 19291 14464 19303 14467
rect 19426 14464 19432 14476
rect 19291 14436 19432 14464
rect 19291 14433 19303 14436
rect 19245 14427 19303 14433
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 19904 14464 19932 14504
rect 19978 14492 19984 14504
rect 20036 14492 20042 14544
rect 20070 14464 20076 14476
rect 19536 14436 19932 14464
rect 20031 14436 20076 14464
rect 19536 14396 19564 14436
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 20162 14424 20168 14476
rect 20220 14464 20226 14476
rect 20625 14467 20683 14473
rect 20625 14464 20637 14467
rect 20220 14436 20637 14464
rect 20220 14424 20226 14436
rect 20625 14433 20637 14436
rect 20671 14433 20683 14467
rect 20990 14464 20996 14476
rect 20951 14436 20996 14464
rect 20625 14427 20683 14433
rect 20990 14424 20996 14436
rect 21048 14424 21054 14476
rect 21266 14424 21272 14476
rect 21324 14464 21330 14476
rect 21361 14467 21419 14473
rect 21361 14464 21373 14467
rect 21324 14436 21373 14464
rect 21324 14424 21330 14436
rect 21361 14433 21373 14436
rect 21407 14433 21419 14467
rect 21361 14427 21419 14433
rect 19076 14368 19564 14396
rect 16393 14359 16451 14365
rect 19610 14356 19616 14408
rect 19668 14396 19674 14408
rect 19797 14399 19855 14405
rect 19797 14396 19809 14399
rect 19668 14368 19809 14396
rect 19668 14356 19674 14368
rect 19797 14365 19809 14368
rect 19843 14365 19855 14399
rect 19978 14396 19984 14408
rect 19939 14368 19984 14396
rect 19797 14359 19855 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 6914 14328 6920 14340
rect 6875 14300 6920 14328
rect 6914 14288 6920 14300
rect 6972 14288 6978 14340
rect 9674 14328 9680 14340
rect 8220 14300 9680 14328
rect 5960 14232 6592 14260
rect 5960 14220 5966 14232
rect 7098 14220 7104 14272
rect 7156 14260 7162 14272
rect 8220 14260 8248 14300
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 13998 14328 14004 14340
rect 9784 14300 10088 14328
rect 13959 14300 14004 14328
rect 7156 14232 8248 14260
rect 8665 14263 8723 14269
rect 7156 14220 7162 14232
rect 8665 14229 8677 14263
rect 8711 14260 8723 14263
rect 8846 14260 8852 14272
rect 8711 14232 8852 14260
rect 8711 14229 8723 14232
rect 8665 14223 8723 14229
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 9490 14220 9496 14272
rect 9548 14260 9554 14272
rect 9784 14260 9812 14300
rect 9548 14232 9812 14260
rect 9548 14220 9554 14232
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 10060 14269 10088 14300
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 16666 14328 16672 14340
rect 15304 14300 16672 14328
rect 10045 14263 10103 14269
rect 9916 14232 9961 14260
rect 9916 14220 9922 14232
rect 10045 14229 10057 14263
rect 10091 14260 10103 14263
rect 15304 14260 15332 14300
rect 16666 14288 16672 14300
rect 16724 14288 16730 14340
rect 17402 14288 17408 14340
rect 17460 14328 17466 14340
rect 18690 14328 18696 14340
rect 17460 14300 18696 14328
rect 17460 14288 17466 14300
rect 18690 14288 18696 14300
rect 18748 14288 18754 14340
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 20622 14328 20628 14340
rect 19484 14300 20628 14328
rect 19484 14288 19490 14300
rect 20622 14288 20628 14300
rect 20680 14288 20686 14340
rect 21174 14328 21180 14340
rect 21135 14300 21180 14328
rect 21174 14288 21180 14300
rect 21232 14288 21238 14340
rect 21542 14328 21548 14340
rect 21503 14300 21548 14328
rect 21542 14288 21548 14300
rect 21600 14288 21606 14340
rect 15838 14260 15844 14272
rect 10091 14232 15332 14260
rect 15799 14232 15844 14260
rect 10091 14229 10103 14232
rect 10045 14223 10103 14229
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 16482 14220 16488 14272
rect 16540 14260 16546 14272
rect 17773 14263 17831 14269
rect 17773 14260 17785 14263
rect 16540 14232 17785 14260
rect 16540 14220 16546 14232
rect 17773 14229 17785 14232
rect 17819 14260 17831 14263
rect 18138 14260 18144 14272
rect 17819 14232 18144 14260
rect 17819 14229 17831 14232
rect 17773 14223 17831 14229
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 20441 14263 20499 14269
rect 20441 14229 20453 14263
rect 20487 14260 20499 14263
rect 20714 14260 20720 14272
rect 20487 14232 20720 14260
rect 20487 14229 20499 14232
rect 20441 14223 20499 14229
rect 20714 14220 20720 14232
rect 20772 14220 20778 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 2130 14056 2136 14068
rect 2091 14028 2136 14056
rect 2130 14016 2136 14028
rect 2188 14016 2194 14068
rect 2332 14028 2636 14056
rect 1673 13991 1731 13997
rect 1673 13957 1685 13991
rect 1719 13988 1731 13991
rect 2332 13988 2360 14028
rect 1719 13960 2360 13988
rect 2409 13991 2467 13997
rect 1719 13957 1731 13960
rect 1673 13951 1731 13957
rect 2409 13957 2421 13991
rect 2455 13988 2467 13991
rect 2455 13960 2544 13988
rect 2455 13957 2467 13960
rect 2409 13951 2467 13957
rect 1394 13812 1400 13864
rect 1452 13852 1458 13864
rect 1489 13855 1547 13861
rect 1489 13852 1501 13855
rect 1452 13824 1501 13852
rect 1452 13812 1458 13824
rect 1489 13821 1501 13824
rect 1535 13821 1547 13855
rect 1762 13852 1768 13864
rect 1723 13824 1768 13852
rect 1489 13815 1547 13821
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 1949 13855 2007 13861
rect 1949 13821 1961 13855
rect 1995 13852 2007 13855
rect 2038 13852 2044 13864
rect 1995 13824 2044 13852
rect 1995 13821 2007 13824
rect 1949 13815 2007 13821
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 2516 13852 2544 13960
rect 2608 13920 2636 14028
rect 2682 14016 2688 14068
rect 2740 14056 2746 14068
rect 2869 14059 2927 14065
rect 2869 14056 2881 14059
rect 2740 14028 2881 14056
rect 2740 14016 2746 14028
rect 2869 14025 2881 14028
rect 2915 14025 2927 14059
rect 2869 14019 2927 14025
rect 4249 14059 4307 14065
rect 4249 14025 4261 14059
rect 4295 14056 4307 14059
rect 4338 14056 4344 14068
rect 4295 14028 4344 14056
rect 4295 14025 4307 14028
rect 4249 14019 4307 14025
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 4798 14016 4804 14068
rect 4856 14056 4862 14068
rect 5169 14059 5227 14065
rect 5169 14056 5181 14059
rect 4856 14028 5181 14056
rect 4856 14016 4862 14028
rect 5169 14025 5181 14028
rect 5215 14025 5227 14059
rect 5169 14019 5227 14025
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 9953 14059 10011 14065
rect 9953 14056 9965 14059
rect 8260 14028 9965 14056
rect 8260 14016 8266 14028
rect 9953 14025 9965 14028
rect 9999 14025 10011 14059
rect 11790 14056 11796 14068
rect 9953 14019 10011 14025
rect 10888 14028 11796 14056
rect 3878 13988 3884 14000
rect 3712 13960 3884 13988
rect 3602 13920 3608 13932
rect 2608 13892 3608 13920
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 3712 13929 3740 13960
rect 3878 13948 3884 13960
rect 3936 13988 3942 14000
rect 6454 13988 6460 14000
rect 3936 13960 5028 13988
rect 3936 13948 3942 13960
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13889 3755 13923
rect 3697 13883 3755 13889
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 2363 13824 2544 13852
rect 2593 13855 2651 13861
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2593 13821 2605 13855
rect 2639 13852 2651 13855
rect 3418 13852 3424 13864
rect 2639 13824 3424 13852
rect 2639 13821 2651 13824
rect 2593 13815 2651 13821
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 3789 13855 3847 13861
rect 3789 13821 3801 13855
rect 3835 13852 3847 13855
rect 4614 13852 4620 13864
rect 3835 13824 4620 13852
rect 3835 13821 3847 13824
rect 3789 13815 3847 13821
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 4798 13852 4804 13864
rect 4759 13824 4804 13852
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 1854 13744 1860 13796
rect 1912 13784 1918 13796
rect 2130 13784 2136 13796
rect 1912 13756 2136 13784
rect 1912 13744 1918 13756
rect 2130 13744 2136 13756
rect 2188 13744 2194 13796
rect 3881 13787 3939 13793
rect 3881 13753 3893 13787
rect 3927 13784 3939 13787
rect 4908 13784 4936 13883
rect 5000 13852 5028 13960
rect 5644 13960 6460 13988
rect 5644 13929 5672 13960
rect 6454 13948 6460 13960
rect 6512 13948 6518 14000
rect 7098 13988 7104 14000
rect 6932 13960 7104 13988
rect 6932 13929 6960 13960
rect 7098 13948 7104 13960
rect 7156 13948 7162 14000
rect 7469 13991 7527 13997
rect 7469 13957 7481 13991
rect 7515 13988 7527 13991
rect 7515 13960 7880 13988
rect 7515 13957 7527 13960
rect 7469 13951 7527 13957
rect 5629 13923 5687 13929
rect 5629 13889 5641 13923
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 6917 13923 6975 13929
rect 6917 13889 6929 13923
rect 6963 13889 6975 13923
rect 6917 13883 6975 13889
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13889 7067 13923
rect 7009 13883 7067 13889
rect 5736 13852 5764 13883
rect 5000 13824 5764 13852
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6144 13824 6776 13852
rect 6144 13812 6150 13824
rect 4982 13784 4988 13796
rect 3927 13756 4384 13784
rect 4908 13756 4988 13784
rect 3927 13753 3939 13756
rect 3881 13747 3939 13753
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 4356 13725 4384 13756
rect 4982 13744 4988 13756
rect 5040 13784 5046 13796
rect 5166 13784 5172 13796
rect 5040 13756 5172 13784
rect 5040 13744 5046 13756
rect 5166 13744 5172 13756
rect 5224 13744 5230 13796
rect 5537 13787 5595 13793
rect 5537 13753 5549 13787
rect 5583 13784 5595 13787
rect 6748 13784 6776 13824
rect 6822 13812 6828 13864
rect 6880 13852 6886 13864
rect 7024 13852 7052 13883
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 6880 13824 7052 13852
rect 7116 13824 7297 13852
rect 6880 13812 6886 13824
rect 7116 13784 7144 13824
rect 7285 13821 7297 13824
rect 7331 13852 7343 13855
rect 7852 13852 7880 13960
rect 8846 13948 8852 14000
rect 8904 13988 8910 14000
rect 8904 13960 10548 13988
rect 8904 13948 8910 13960
rect 8864 13920 8892 13948
rect 9214 13920 9220 13932
rect 8772 13892 8892 13920
rect 9175 13892 9220 13920
rect 8294 13852 8300 13864
rect 7331 13824 7788 13852
rect 7852 13824 8300 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 5583 13756 6500 13784
rect 5583 13753 5595 13756
rect 5537 13747 5595 13753
rect 2685 13719 2743 13725
rect 2685 13716 2697 13719
rect 1820 13688 2697 13716
rect 1820 13676 1826 13688
rect 2685 13685 2697 13688
rect 2731 13685 2743 13719
rect 2685 13679 2743 13685
rect 4341 13719 4399 13725
rect 4341 13685 4353 13719
rect 4387 13685 4399 13719
rect 4706 13716 4712 13728
rect 4667 13688 4712 13716
rect 4341 13679 4399 13685
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 6472 13725 6500 13756
rect 6748 13756 7144 13784
rect 7760 13784 7788 13824
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 8570 13852 8576 13864
rect 8628 13861 8634 13864
rect 8628 13855 8651 13861
rect 8503 13824 8576 13852
rect 8570 13812 8576 13824
rect 8639 13852 8651 13855
rect 8772 13852 8800 13892
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 9401 13923 9459 13929
rect 9401 13889 9413 13923
rect 9447 13920 9459 13923
rect 9447 13892 9812 13920
rect 9447 13889 9459 13892
rect 9401 13883 9459 13889
rect 8639 13824 8800 13852
rect 8849 13855 8907 13861
rect 8639 13821 8651 13824
rect 8628 13815 8651 13821
rect 8849 13821 8861 13855
rect 8895 13852 8907 13855
rect 9122 13852 9128 13864
rect 8895 13824 9128 13852
rect 8895 13821 8907 13824
rect 8849 13815 8907 13821
rect 8628 13812 8634 13815
rect 9122 13812 9128 13824
rect 9180 13852 9186 13864
rect 9582 13852 9588 13864
rect 9180 13824 9588 13852
rect 9180 13812 9186 13824
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 9784 13852 9812 13892
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 10520 13929 10548 13960
rect 10413 13923 10471 13929
rect 10413 13920 10425 13923
rect 9916 13892 10425 13920
rect 9916 13880 9922 13892
rect 10413 13889 10425 13892
rect 10459 13889 10471 13923
rect 10413 13883 10471 13889
rect 10505 13923 10563 13929
rect 10505 13889 10517 13923
rect 10551 13889 10563 13923
rect 10888 13920 10916 14028
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 13538 14056 13544 14068
rect 13499 14028 13544 14056
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 14734 14016 14740 14068
rect 14792 14056 14798 14068
rect 14921 14059 14979 14065
rect 14921 14056 14933 14059
rect 14792 14028 14933 14056
rect 14792 14016 14798 14028
rect 14921 14025 14933 14028
rect 14967 14025 14979 14059
rect 18417 14059 18475 14065
rect 18417 14056 18429 14059
rect 14921 14019 14979 14025
rect 15304 14028 18429 14056
rect 11517 13991 11575 13997
rect 11517 13957 11529 13991
rect 11563 13988 11575 13991
rect 12713 13991 12771 13997
rect 11563 13960 12296 13988
rect 11563 13957 11575 13960
rect 11517 13951 11575 13957
rect 10505 13883 10563 13889
rect 10796 13892 10916 13920
rect 10965 13923 11023 13929
rect 10796 13852 10824 13892
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 11054 13920 11060 13932
rect 11011 13892 11060 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 11054 13880 11060 13892
rect 11112 13880 11118 13932
rect 12268 13929 12296 13960
rect 12713 13957 12725 13991
rect 12759 13988 12771 13991
rect 15304 13988 15332 14028
rect 18417 14025 18429 14028
rect 18463 14025 18475 14059
rect 18417 14019 18475 14025
rect 18509 14059 18567 14065
rect 18509 14025 18521 14059
rect 18555 14056 18567 14059
rect 18555 14028 21404 14056
rect 18555 14025 18567 14028
rect 18509 14019 18567 14025
rect 15749 13991 15807 13997
rect 15749 13988 15761 13991
rect 12759 13960 15332 13988
rect 15396 13960 15761 13988
rect 12759 13957 12771 13960
rect 12713 13951 12771 13957
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13889 12311 13923
rect 12253 13883 12311 13889
rect 11146 13852 11152 13864
rect 9784 13824 10824 13852
rect 11107 13824 11152 13852
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 12176 13852 12204 13883
rect 12802 13880 12808 13932
rect 12860 13920 12866 13932
rect 12897 13923 12955 13929
rect 12897 13920 12909 13923
rect 12860 13892 12909 13920
rect 12860 13880 12866 13892
rect 12897 13889 12909 13892
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 12986 13880 12992 13932
rect 13044 13920 13050 13932
rect 13538 13920 13544 13932
rect 13044 13892 13544 13920
rect 13044 13880 13050 13892
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 15396 13929 15424 13960
rect 15749 13957 15761 13960
rect 15795 13957 15807 13991
rect 16945 13991 17003 13997
rect 16945 13988 16957 13991
rect 15749 13951 15807 13957
rect 16316 13960 16957 13988
rect 16316 13932 16344 13960
rect 16945 13957 16957 13960
rect 16991 13957 17003 13991
rect 18524 13988 18552 14019
rect 16945 13951 17003 13957
rect 18340 13960 18552 13988
rect 20717 13991 20775 13997
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13889 15439 13923
rect 15562 13920 15568 13932
rect 15523 13892 15568 13920
rect 15381 13883 15439 13889
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 16298 13920 16304 13932
rect 16259 13892 16304 13920
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 18340 13920 18368 13960
rect 20717 13957 20729 13991
rect 20763 13988 20775 13991
rect 20763 13960 21312 13988
rect 20763 13957 20775 13960
rect 20717 13951 20775 13957
rect 20073 13923 20131 13929
rect 20073 13920 20085 13923
rect 18248 13892 18368 13920
rect 19812 13892 20085 13920
rect 12176 13824 12434 13852
rect 12250 13784 12256 13796
rect 7760 13756 12256 13784
rect 6457 13719 6515 13725
rect 6457 13685 6469 13719
rect 6503 13685 6515 13719
rect 6748 13716 6776 13756
rect 12250 13744 12256 13756
rect 12308 13744 12314 13796
rect 12406 13784 12434 13824
rect 12618 13812 12624 13864
rect 12676 13852 12682 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12676 13824 13093 13852
rect 12676 13812 12682 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 15194 13852 15200 13864
rect 14875 13824 15200 13852
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15838 13852 15844 13864
rect 15335 13824 15844 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 16114 13812 16120 13864
rect 16172 13852 16178 13864
rect 16209 13855 16267 13861
rect 16209 13852 16221 13855
rect 16172 13824 16221 13852
rect 16172 13812 16178 13824
rect 16209 13821 16221 13824
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 18069 13855 18127 13861
rect 18069 13821 18081 13855
rect 18115 13852 18127 13855
rect 18248 13852 18276 13892
rect 18115 13824 18276 13852
rect 18325 13855 18383 13861
rect 18115 13821 18127 13824
rect 18069 13815 18127 13821
rect 18325 13821 18337 13855
rect 18371 13821 18383 13855
rect 18325 13815 18383 13821
rect 18417 13855 18475 13861
rect 18417 13821 18429 13855
rect 18463 13852 18475 13855
rect 19334 13852 19340 13864
rect 18463 13824 19340 13852
rect 18463 13821 18475 13824
rect 18417 13815 18475 13821
rect 12986 13784 12992 13796
rect 12406 13756 12992 13784
rect 12986 13744 12992 13756
rect 13044 13744 13050 13796
rect 15654 13784 15660 13796
rect 13096 13756 15660 13784
rect 13096 13728 13124 13756
rect 15654 13744 15660 13756
rect 15712 13744 15718 13796
rect 16574 13784 16580 13796
rect 16535 13756 16580 13784
rect 16574 13744 16580 13756
rect 16632 13744 16638 13796
rect 17586 13744 17592 13796
rect 17644 13784 17650 13796
rect 18340 13784 18368 13815
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19610 13812 19616 13864
rect 19668 13861 19674 13864
rect 19668 13852 19680 13861
rect 19812 13852 19840 13892
rect 20073 13889 20085 13892
rect 20119 13889 20131 13923
rect 20073 13883 20131 13889
rect 20346 13880 20352 13932
rect 20404 13920 20410 13932
rect 21174 13920 21180 13932
rect 20404 13892 21180 13920
rect 20404 13880 20410 13892
rect 21174 13880 21180 13892
rect 21232 13880 21238 13932
rect 21284 13929 21312 13960
rect 21376 13929 21404 14028
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 21361 13923 21419 13929
rect 21361 13889 21373 13923
rect 21407 13889 21419 13923
rect 21361 13883 21419 13889
rect 19668 13824 19840 13852
rect 19889 13855 19947 13861
rect 19668 13815 19680 13824
rect 19889 13821 19901 13855
rect 19935 13821 19947 13855
rect 19889 13815 19947 13821
rect 20257 13855 20315 13861
rect 20257 13821 20269 13855
rect 20303 13852 20315 13855
rect 20438 13852 20444 13864
rect 20303 13824 20444 13852
rect 20303 13821 20315 13824
rect 20257 13815 20315 13821
rect 19668 13812 19674 13815
rect 17644 13756 19104 13784
rect 17644 13744 17650 13756
rect 19076 13728 19104 13756
rect 6825 13719 6883 13725
rect 6825 13716 6837 13719
rect 6748 13688 6837 13716
rect 6457 13679 6515 13685
rect 6825 13685 6837 13688
rect 6871 13685 6883 13719
rect 6825 13679 6883 13685
rect 8662 13676 8668 13728
rect 8720 13716 8726 13728
rect 9490 13716 9496 13728
rect 8720 13688 9496 13716
rect 8720 13676 8726 13688
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 9861 13719 9919 13725
rect 9861 13685 9873 13719
rect 9907 13716 9919 13719
rect 10321 13719 10379 13725
rect 10321 13716 10333 13719
rect 9907 13688 10333 13716
rect 9907 13685 9919 13688
rect 9861 13679 9919 13685
rect 10321 13685 10333 13688
rect 10367 13685 10379 13719
rect 10321 13679 10379 13685
rect 10962 13676 10968 13728
rect 11020 13716 11026 13728
rect 11057 13719 11115 13725
rect 11057 13716 11069 13719
rect 11020 13688 11069 13716
rect 11020 13676 11026 13688
rect 11057 13685 11069 13688
rect 11103 13685 11115 13719
rect 11057 13679 11115 13685
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 12345 13719 12403 13725
rect 12345 13716 12357 13719
rect 11848 13688 12357 13716
rect 11848 13676 11854 13688
rect 12345 13685 12357 13688
rect 12391 13685 12403 13719
rect 12345 13679 12403 13685
rect 13078 13676 13084 13728
rect 13136 13676 13142 13728
rect 13173 13719 13231 13725
rect 13173 13685 13185 13719
rect 13219 13716 13231 13719
rect 13446 13716 13452 13728
rect 13219 13688 13452 13716
rect 13219 13685 13231 13688
rect 13173 13679 13231 13685
rect 13446 13676 13452 13688
rect 13504 13716 13510 13728
rect 13633 13719 13691 13725
rect 13633 13716 13645 13719
rect 13504 13688 13645 13716
rect 13504 13676 13510 13688
rect 13633 13685 13645 13688
rect 13679 13685 13691 13719
rect 13633 13679 13691 13685
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 16117 13719 16175 13725
rect 16117 13716 16129 13719
rect 15252 13688 16129 13716
rect 15252 13676 15258 13688
rect 16117 13685 16129 13688
rect 16163 13716 16175 13719
rect 16482 13716 16488 13728
rect 16163 13688 16488 13716
rect 16163 13685 16175 13688
rect 16117 13679 16175 13685
rect 16482 13676 16488 13688
rect 16540 13676 16546 13728
rect 19058 13676 19064 13728
rect 19116 13716 19122 13728
rect 19904 13716 19932 13815
rect 20438 13812 20444 13824
rect 20496 13812 20502 13864
rect 20714 13744 20720 13796
rect 20772 13784 20778 13796
rect 21177 13787 21235 13793
rect 21177 13784 21189 13787
rect 20772 13756 21189 13784
rect 20772 13744 20778 13756
rect 21177 13753 21189 13756
rect 21223 13753 21235 13787
rect 21177 13747 21235 13753
rect 19116 13688 19932 13716
rect 19116 13676 19122 13688
rect 20346 13676 20352 13728
rect 20404 13716 20410 13728
rect 20404 13688 20449 13716
rect 20404 13676 20410 13688
rect 20622 13676 20628 13728
rect 20680 13716 20686 13728
rect 20809 13719 20867 13725
rect 20809 13716 20821 13719
rect 20680 13688 20821 13716
rect 20680 13676 20686 13688
rect 20809 13685 20821 13688
rect 20855 13685 20867 13719
rect 20809 13679 20867 13685
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 4614 13512 4620 13524
rect 4575 13484 4620 13512
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 4706 13472 4712 13524
rect 4764 13512 4770 13524
rect 5445 13515 5503 13521
rect 5445 13512 5457 13515
rect 4764 13484 5457 13512
rect 4764 13472 4770 13484
rect 5445 13481 5457 13484
rect 5491 13481 5503 13515
rect 5445 13475 5503 13481
rect 7193 13515 7251 13521
rect 7193 13481 7205 13515
rect 7239 13512 7251 13515
rect 7558 13512 7564 13524
rect 7239 13484 7564 13512
rect 7239 13481 7251 13484
rect 7193 13475 7251 13481
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 7742 13512 7748 13524
rect 7703 13484 7748 13512
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 8757 13515 8815 13521
rect 8757 13512 8769 13515
rect 8536 13484 8769 13512
rect 8536 13472 8542 13484
rect 8757 13481 8769 13484
rect 8803 13481 8815 13515
rect 14185 13515 14243 13521
rect 8757 13475 8815 13481
rect 8956 13484 12434 13512
rect 1486 13444 1492 13456
rect 1399 13416 1492 13444
rect 1486 13404 1492 13416
rect 1544 13444 1550 13456
rect 2133 13447 2191 13453
rect 2133 13444 2145 13447
rect 1544 13416 2145 13444
rect 1544 13404 1550 13416
rect 2133 13413 2145 13416
rect 2179 13413 2191 13447
rect 2133 13407 2191 13413
rect 2240 13416 8708 13444
rect 1762 13336 1768 13388
rect 1820 13376 1826 13388
rect 1857 13379 1915 13385
rect 1857 13376 1869 13379
rect 1820 13348 1869 13376
rect 1820 13336 1826 13348
rect 1857 13345 1869 13348
rect 1903 13345 1915 13379
rect 1857 13339 1915 13345
rect 2041 13379 2099 13385
rect 2041 13345 2053 13379
rect 2087 13376 2099 13379
rect 2240 13376 2268 13416
rect 2087 13348 2268 13376
rect 2584 13379 2642 13385
rect 2087 13345 2099 13348
rect 2041 13339 2099 13345
rect 2584 13345 2596 13379
rect 2630 13376 2642 13379
rect 2958 13376 2964 13388
rect 2630 13348 2964 13376
rect 2630 13345 2642 13348
rect 2584 13339 2642 13345
rect 2958 13336 2964 13348
rect 3016 13336 3022 13388
rect 4982 13376 4988 13388
rect 4943 13348 4988 13376
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5074 13336 5080 13388
rect 5132 13376 5138 13388
rect 5132 13348 5764 13376
rect 5132 13336 5138 13348
rect 2314 13308 2320 13320
rect 2275 13280 2320 13308
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 5166 13308 5172 13320
rect 5127 13280 5172 13308
rect 5166 13268 5172 13280
rect 5224 13268 5230 13320
rect 5736 13308 5764 13348
rect 5810 13336 5816 13388
rect 5868 13376 5874 13388
rect 7285 13379 7343 13385
rect 7285 13376 7297 13379
rect 5868 13348 7297 13376
rect 5868 13336 5874 13348
rect 7285 13345 7297 13348
rect 7331 13345 7343 13379
rect 7285 13339 7343 13345
rect 7558 13336 7564 13388
rect 7616 13376 7622 13388
rect 8113 13379 8171 13385
rect 8113 13376 8125 13379
rect 7616 13348 8125 13376
rect 7616 13336 7622 13348
rect 8113 13345 8125 13348
rect 8159 13345 8171 13379
rect 8113 13339 8171 13345
rect 5736 13280 5856 13308
rect 1673 13243 1731 13249
rect 1673 13209 1685 13243
rect 1719 13240 1731 13243
rect 3697 13243 3755 13249
rect 1719 13212 2268 13240
rect 1719 13209 1731 13212
rect 1673 13203 1731 13209
rect 2240 13172 2268 13212
rect 3697 13209 3709 13243
rect 3743 13240 3755 13243
rect 5184 13240 5212 13268
rect 3743 13212 5212 13240
rect 3743 13209 3755 13212
rect 3697 13203 3755 13209
rect 3602 13172 3608 13184
rect 2240 13144 3608 13172
rect 3602 13132 3608 13144
rect 3660 13132 3666 13184
rect 5828 13181 5856 13280
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6972 13280 7021 13308
rect 6972 13268 6978 13280
rect 7009 13277 7021 13280
rect 7055 13277 7067 13311
rect 8205 13311 8263 13317
rect 8205 13308 8217 13311
rect 7009 13271 7067 13277
rect 7668 13280 8217 13308
rect 7668 13249 7696 13280
rect 8205 13277 8217 13280
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 8570 13308 8576 13320
rect 8435 13280 8576 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 8680 13308 8708 13416
rect 8956 13385 8984 13484
rect 9852 13447 9910 13453
rect 9852 13413 9864 13447
rect 9898 13444 9910 13447
rect 12406 13444 12434 13484
rect 14185 13481 14197 13515
rect 14231 13512 14243 13515
rect 18969 13515 19027 13521
rect 14231 13484 18920 13512
rect 14231 13481 14243 13484
rect 14185 13475 14243 13481
rect 13081 13447 13139 13453
rect 13081 13444 13093 13447
rect 9898 13416 12296 13444
rect 12406 13416 13093 13444
rect 9898 13413 9910 13416
rect 9852 13407 9910 13413
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 9048 13348 10640 13376
rect 9048 13308 9076 13348
rect 9582 13308 9588 13320
rect 8680 13280 9076 13308
rect 9543 13280 9588 13308
rect 9582 13268 9588 13280
rect 9640 13268 9646 13320
rect 10612 13308 10640 13348
rect 10778 13336 10784 13388
rect 10836 13376 10842 13388
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 10836 13348 11345 13376
rect 10836 13336 10842 13348
rect 11333 13345 11345 13348
rect 11379 13345 11391 13379
rect 12268 13376 12296 13416
rect 13081 13413 13093 13416
rect 13127 13444 13139 13447
rect 15470 13444 15476 13456
rect 13127 13416 14412 13444
rect 13127 13413 13139 13416
rect 13081 13407 13139 13413
rect 13354 13376 13360 13388
rect 12268 13348 13360 13376
rect 11333 13339 11391 13345
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 14384 13385 14412 13416
rect 14568 13416 15476 13444
rect 13817 13379 13875 13385
rect 13817 13345 13829 13379
rect 13863 13345 13875 13379
rect 13817 13339 13875 13345
rect 14369 13379 14427 13385
rect 14369 13345 14381 13379
rect 14415 13345 14427 13379
rect 14369 13339 14427 13345
rect 13078 13308 13084 13320
rect 10612 13280 13084 13308
rect 13078 13268 13084 13280
rect 13136 13268 13142 13320
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13277 13599 13311
rect 13541 13271 13599 13277
rect 7653 13243 7711 13249
rect 7653 13209 7665 13243
rect 7699 13209 7711 13243
rect 13556 13240 13584 13271
rect 13630 13268 13636 13320
rect 13688 13308 13694 13320
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13688 13280 13737 13308
rect 13688 13268 13694 13280
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 13832 13308 13860 13339
rect 14568 13308 14596 13416
rect 15470 13404 15476 13416
rect 15528 13404 15534 13456
rect 15746 13404 15752 13456
rect 15804 13444 15810 13456
rect 15850 13447 15908 13453
rect 15850 13444 15862 13447
rect 15804 13416 15862 13444
rect 15804 13404 15810 13416
rect 15850 13413 15862 13416
rect 15896 13413 15908 13447
rect 18892 13444 18920 13484
rect 18969 13481 18981 13515
rect 19015 13512 19027 13515
rect 19610 13512 19616 13524
rect 19015 13484 19616 13512
rect 19015 13481 19027 13484
rect 18969 13475 19027 13481
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 19797 13515 19855 13521
rect 19797 13481 19809 13515
rect 19843 13481 19855 13515
rect 19797 13475 19855 13481
rect 19812 13444 19840 13475
rect 20070 13472 20076 13524
rect 20128 13512 20134 13524
rect 20165 13515 20223 13521
rect 20165 13512 20177 13515
rect 20128 13484 20177 13512
rect 20128 13472 20134 13484
rect 20165 13481 20177 13484
rect 20211 13481 20223 13515
rect 20622 13512 20628 13524
rect 20583 13484 20628 13512
rect 20165 13475 20223 13481
rect 20622 13472 20628 13484
rect 20680 13472 20686 13524
rect 21177 13515 21235 13521
rect 21177 13481 21189 13515
rect 21223 13512 21235 13515
rect 21358 13512 21364 13524
rect 21223 13484 21364 13512
rect 21223 13481 21235 13484
rect 21177 13475 21235 13481
rect 21358 13472 21364 13484
rect 21416 13472 21422 13524
rect 18892 13416 19748 13444
rect 19812 13416 21036 13444
rect 15850 13407 15908 13413
rect 17845 13379 17903 13385
rect 17845 13376 17857 13379
rect 13832 13280 14596 13308
rect 14660 13348 17857 13376
rect 13725 13271 13783 13277
rect 14090 13240 14096 13252
rect 7653 13203 7711 13209
rect 7760 13212 8708 13240
rect 13556 13212 14096 13240
rect 5813 13175 5871 13181
rect 5813 13141 5825 13175
rect 5859 13172 5871 13175
rect 7760 13172 7788 13212
rect 5859 13144 7788 13172
rect 5859 13141 5871 13144
rect 5813 13135 5871 13141
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 8573 13175 8631 13181
rect 8573 13172 8585 13175
rect 7892 13144 8585 13172
rect 7892 13132 7898 13144
rect 8573 13141 8585 13144
rect 8619 13141 8631 13175
rect 8680 13172 8708 13212
rect 14090 13200 14096 13212
rect 14148 13200 14154 13252
rect 14550 13240 14556 13252
rect 14511 13212 14556 13240
rect 14550 13200 14556 13212
rect 14608 13200 14614 13252
rect 10870 13172 10876 13184
rect 8680 13144 10876 13172
rect 8573 13135 8631 13141
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 10965 13175 11023 13181
rect 10965 13141 10977 13175
rect 11011 13172 11023 13175
rect 11054 13172 11060 13184
rect 11011 13144 11060 13172
rect 11011 13141 11023 13144
rect 10965 13135 11023 13141
rect 11054 13132 11060 13144
rect 11112 13172 11118 13184
rect 11790 13172 11796 13184
rect 11112 13144 11796 13172
rect 11112 13132 11118 13144
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 14660 13172 14688 13348
rect 17845 13345 17857 13348
rect 17891 13376 17903 13379
rect 17891 13348 18644 13376
rect 17891 13345 17903 13348
rect 17845 13339 17903 13345
rect 16117 13311 16175 13317
rect 16117 13277 16129 13311
rect 16163 13308 16175 13311
rect 17586 13308 17592 13320
rect 16163 13280 17592 13308
rect 16163 13277 16175 13280
rect 16117 13271 16175 13277
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 18616 13308 18644 13348
rect 18966 13336 18972 13388
rect 19024 13376 19030 13388
rect 19613 13379 19671 13385
rect 19613 13376 19625 13379
rect 19024 13348 19625 13376
rect 19024 13336 19030 13348
rect 19613 13345 19625 13348
rect 19659 13345 19671 13379
rect 19720 13376 19748 13416
rect 19889 13379 19947 13385
rect 19889 13376 19901 13379
rect 19720 13348 19901 13376
rect 19613 13339 19671 13345
rect 19889 13345 19901 13348
rect 19935 13345 19947 13379
rect 19889 13339 19947 13345
rect 20533 13379 20591 13385
rect 20533 13345 20545 13379
rect 20579 13376 20591 13379
rect 20898 13376 20904 13388
rect 20579 13348 20904 13376
rect 20579 13345 20591 13348
rect 20533 13339 20591 13345
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 21008 13385 21036 13416
rect 20993 13379 21051 13385
rect 20993 13345 21005 13379
rect 21039 13345 21051 13379
rect 21542 13376 21548 13388
rect 21503 13348 21548 13376
rect 20993 13339 21051 13345
rect 21542 13336 21548 13348
rect 21600 13336 21606 13388
rect 20438 13308 20444 13320
rect 18616 13280 20444 13308
rect 20438 13268 20444 13280
rect 20496 13308 20502 13320
rect 20717 13311 20775 13317
rect 20717 13308 20729 13311
rect 20496 13280 20729 13308
rect 20496 13268 20502 13280
rect 20717 13277 20729 13280
rect 20763 13277 20775 13311
rect 20717 13271 20775 13277
rect 19610 13240 19616 13252
rect 19306 13212 19616 13240
rect 13044 13144 14688 13172
rect 14737 13175 14795 13181
rect 13044 13132 13050 13144
rect 14737 13141 14749 13175
rect 14783 13172 14795 13175
rect 14918 13172 14924 13184
rect 14783 13144 14924 13172
rect 14783 13141 14795 13144
rect 14737 13135 14795 13141
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 16850 13132 16856 13184
rect 16908 13172 16914 13184
rect 19153 13175 19211 13181
rect 19153 13172 19165 13175
rect 16908 13144 19165 13172
rect 16908 13132 16914 13144
rect 19153 13141 19165 13144
rect 19199 13172 19211 13175
rect 19306 13172 19334 13212
rect 19610 13200 19616 13212
rect 19668 13200 19674 13252
rect 20073 13243 20131 13249
rect 20073 13209 20085 13243
rect 20119 13240 20131 13243
rect 20162 13240 20168 13252
rect 20119 13212 20168 13240
rect 20119 13209 20131 13212
rect 20073 13203 20131 13209
rect 20162 13200 20168 13212
rect 20220 13200 20226 13252
rect 21082 13200 21088 13252
rect 21140 13240 21146 13252
rect 21361 13243 21419 13249
rect 21361 13240 21373 13243
rect 21140 13212 21373 13240
rect 21140 13200 21146 13212
rect 21361 13209 21373 13212
rect 21407 13209 21419 13243
rect 21361 13203 21419 13209
rect 19199 13144 19334 13172
rect 19429 13175 19487 13181
rect 19199 13141 19211 13144
rect 19153 13135 19211 13141
rect 19429 13141 19441 13175
rect 19475 13172 19487 13175
rect 21542 13172 21548 13184
rect 19475 13144 21548 13172
rect 19475 13141 19487 13144
rect 19429 13135 19487 13141
rect 21542 13132 21548 13144
rect 21600 13132 21606 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 2130 12968 2136 12980
rect 1627 12940 2136 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 2130 12928 2136 12940
rect 2188 12928 2194 12980
rect 2409 12971 2467 12977
rect 2409 12937 2421 12971
rect 2455 12968 2467 12971
rect 2590 12968 2596 12980
rect 2455 12940 2596 12968
rect 2455 12937 2467 12940
rect 2409 12931 2467 12937
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 3510 12968 3516 12980
rect 2832 12940 3516 12968
rect 2832 12928 2838 12940
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 3786 12968 3792 12980
rect 3747 12940 3792 12968
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 7558 12968 7564 12980
rect 7519 12940 7564 12968
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 12986 12928 12992 12980
rect 13044 12968 13050 12980
rect 13081 12971 13139 12977
rect 13081 12968 13093 12971
rect 13044 12940 13093 12968
rect 13044 12928 13050 12940
rect 13081 12937 13093 12940
rect 13127 12937 13139 12971
rect 13630 12968 13636 12980
rect 13591 12940 13636 12968
rect 13081 12931 13139 12937
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 14366 12928 14372 12980
rect 14424 12968 14430 12980
rect 14734 12968 14740 12980
rect 14424 12940 14740 12968
rect 14424 12928 14430 12940
rect 14734 12928 14740 12940
rect 14792 12968 14798 12980
rect 19610 12968 19616 12980
rect 14792 12940 19616 12968
rect 14792 12928 14798 12940
rect 19610 12928 19616 12940
rect 19668 12928 19674 12980
rect 19978 12928 19984 12980
rect 20036 12968 20042 12980
rect 20165 12971 20223 12977
rect 20165 12968 20177 12971
rect 20036 12940 20177 12968
rect 20036 12928 20042 12940
rect 20165 12937 20177 12940
rect 20211 12937 20223 12971
rect 20165 12931 20223 12937
rect 20530 12928 20536 12980
rect 20588 12968 20594 12980
rect 21361 12971 21419 12977
rect 21361 12968 21373 12971
rect 20588 12940 21373 12968
rect 20588 12928 20594 12940
rect 21361 12937 21373 12940
rect 21407 12937 21419 12971
rect 21361 12931 21419 12937
rect 1394 12860 1400 12912
rect 1452 12900 1458 12912
rect 3329 12903 3387 12909
rect 3329 12900 3341 12903
rect 1452 12872 3341 12900
rect 1452 12860 1458 12872
rect 3329 12869 3341 12872
rect 3375 12869 3387 12903
rect 3329 12863 3387 12869
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12832 1915 12835
rect 1946 12832 1952 12844
rect 1903 12804 1952 12832
rect 1903 12801 1915 12804
rect 1857 12795 1915 12801
rect 1946 12792 1952 12804
rect 2004 12832 2010 12844
rect 2130 12832 2136 12844
rect 2004 12804 2136 12832
rect 2004 12792 2010 12804
rect 2130 12792 2136 12804
rect 2188 12792 2194 12844
rect 2406 12792 2412 12844
rect 2464 12832 2470 12844
rect 2593 12835 2651 12841
rect 2593 12832 2605 12835
rect 2464 12804 2605 12832
rect 2464 12792 2470 12804
rect 2593 12801 2605 12804
rect 2639 12801 2651 12835
rect 2593 12795 2651 12801
rect 2777 12835 2835 12841
rect 2777 12801 2789 12835
rect 2823 12832 2835 12835
rect 3804 12832 3832 12928
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 9640 12872 11744 12900
rect 9640 12860 9646 12872
rect 5350 12832 5356 12844
rect 2823 12804 3832 12832
rect 5311 12804 5356 12832
rect 2823 12801 2835 12804
rect 2777 12795 2835 12801
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 6914 12832 6920 12844
rect 6875 12804 6920 12832
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 10229 12835 10287 12841
rect 10229 12832 10241 12835
rect 9824 12804 10241 12832
rect 9824 12792 9830 12804
rect 10229 12801 10241 12804
rect 10275 12801 10287 12835
rect 10229 12795 10287 12801
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12832 10747 12835
rect 11606 12832 11612 12844
rect 10735 12804 11612 12832
rect 10735 12801 10747 12804
rect 10689 12795 10747 12801
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 11716 12841 11744 12872
rect 13354 12860 13360 12912
rect 13412 12900 13418 12912
rect 16942 12900 16948 12912
rect 13412 12872 16948 12900
rect 13412 12860 13418 12872
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 18322 12860 18328 12912
rect 18380 12900 18386 12912
rect 20622 12900 20628 12912
rect 18380 12872 20628 12900
rect 18380 12860 18386 12872
rect 20622 12860 20628 12872
rect 20680 12860 20686 12912
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12832 14335 12835
rect 14366 12832 14372 12844
rect 14323 12804 14372 12832
rect 14323 12801 14335 12804
rect 14277 12795 14335 12801
rect 14366 12792 14372 12804
rect 14424 12792 14430 12844
rect 14918 12792 14924 12844
rect 14976 12832 14982 12844
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 14976 12804 15209 12832
rect 14976 12792 14982 12804
rect 15197 12801 15209 12804
rect 15243 12832 15255 12835
rect 15286 12832 15292 12844
rect 15243 12804 15292 12832
rect 15243 12801 15255 12804
rect 15197 12795 15255 12801
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 18969 12835 19027 12841
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 2041 12767 2099 12773
rect 2041 12733 2053 12767
rect 2087 12764 2099 12767
rect 2958 12764 2964 12776
rect 2087 12736 2964 12764
rect 2087 12733 2099 12736
rect 2041 12727 2099 12733
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 3602 12724 3608 12776
rect 3660 12764 3666 12776
rect 8205 12767 8263 12773
rect 3660 12736 7788 12764
rect 3660 12724 3666 12736
rect 1949 12699 2007 12705
rect 1949 12665 1961 12699
rect 1995 12696 2007 12699
rect 3050 12696 3056 12708
rect 1995 12668 3056 12696
rect 1995 12665 2007 12668
rect 1949 12659 2007 12665
rect 3050 12656 3056 12668
rect 3108 12656 3114 12708
rect 5442 12656 5448 12708
rect 5500 12696 5506 12708
rect 7101 12699 7159 12705
rect 7101 12696 7113 12699
rect 5500 12668 7113 12696
rect 5500 12656 5506 12668
rect 7101 12665 7113 12668
rect 7147 12665 7159 12699
rect 7101 12659 7159 12665
rect 7193 12699 7251 12705
rect 7193 12665 7205 12699
rect 7239 12696 7251 12699
rect 7653 12699 7711 12705
rect 7653 12696 7665 12699
rect 7239 12668 7665 12696
rect 7239 12665 7251 12668
rect 7193 12659 7251 12665
rect 7653 12665 7665 12668
rect 7699 12665 7711 12699
rect 7653 12659 7711 12665
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 2869 12631 2927 12637
rect 2869 12628 2881 12631
rect 2832 12600 2881 12628
rect 2832 12588 2838 12600
rect 2869 12597 2881 12600
rect 2915 12597 2927 12631
rect 3234 12628 3240 12640
rect 3195 12600 3240 12628
rect 2869 12591 2927 12597
rect 3234 12588 3240 12600
rect 3292 12588 3298 12640
rect 4706 12628 4712 12640
rect 4667 12600 4712 12628
rect 4706 12588 4712 12600
rect 4764 12588 4770 12640
rect 5074 12628 5080 12640
rect 5035 12600 5080 12628
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12628 5227 12631
rect 6546 12628 6552 12640
rect 5215 12600 6552 12628
rect 5215 12597 5227 12600
rect 5169 12591 5227 12597
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 7760 12628 7788 12736
rect 8205 12733 8217 12767
rect 8251 12764 8263 12767
rect 8754 12764 8760 12776
rect 8251 12736 8760 12764
rect 8251 12733 8263 12736
rect 8205 12727 8263 12733
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 10042 12764 10048 12776
rect 10003 12736 10048 12764
rect 10042 12724 10048 12736
rect 10100 12764 10106 12776
rect 10873 12767 10931 12773
rect 10873 12764 10885 12767
rect 10100 12736 10885 12764
rect 10100 12724 10106 12736
rect 10873 12733 10885 12736
rect 10919 12733 10931 12767
rect 10873 12727 10931 12733
rect 11790 12724 11796 12776
rect 11848 12764 11854 12776
rect 11957 12767 12015 12773
rect 11957 12764 11969 12767
rect 11848 12736 11969 12764
rect 11848 12724 11854 12736
rect 11957 12733 11969 12736
rect 12003 12733 12015 12767
rect 16850 12764 16856 12776
rect 11957 12727 12015 12733
rect 12268 12736 16856 12764
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 8450 12699 8508 12705
rect 8450 12696 8462 12699
rect 8352 12668 8462 12696
rect 8352 12656 8358 12668
rect 8450 12665 8462 12668
rect 8496 12665 8508 12699
rect 12268 12696 12296 12736
rect 16850 12724 16856 12736
rect 16908 12724 16914 12776
rect 17034 12724 17040 12776
rect 17092 12764 17098 12776
rect 18325 12767 18383 12773
rect 18325 12764 18337 12767
rect 17092 12736 18337 12764
rect 17092 12724 17098 12736
rect 18325 12733 18337 12736
rect 18371 12733 18383 12767
rect 18325 12727 18383 12733
rect 18414 12724 18420 12776
rect 18472 12724 18478 12776
rect 14093 12699 14151 12705
rect 14093 12696 14105 12699
rect 8450 12659 8508 12665
rect 8588 12668 12296 12696
rect 12406 12668 14105 12696
rect 8588 12628 8616 12668
rect 7760 12600 8616 12628
rect 9490 12588 9496 12640
rect 9548 12628 9554 12640
rect 9585 12631 9643 12637
rect 9585 12628 9597 12631
rect 9548 12600 9597 12628
rect 9548 12588 9554 12600
rect 9585 12597 9597 12600
rect 9631 12597 9643 12631
rect 9585 12591 9643 12597
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10134 12628 10140 12640
rect 9732 12600 9777 12628
rect 10095 12600 10140 12628
rect 9732 12588 9738 12600
rect 10134 12588 10140 12600
rect 10192 12628 10198 12640
rect 10781 12631 10839 12637
rect 10781 12628 10793 12631
rect 10192 12600 10793 12628
rect 10192 12588 10198 12600
rect 10781 12597 10793 12600
rect 10827 12597 10839 12631
rect 10781 12591 10839 12597
rect 11241 12631 11299 12637
rect 11241 12597 11253 12631
rect 11287 12628 11299 12631
rect 12406 12628 12434 12668
rect 14093 12665 14105 12668
rect 14139 12665 14151 12699
rect 14093 12659 14151 12665
rect 14274 12656 14280 12708
rect 14332 12696 14338 12708
rect 14829 12699 14887 12705
rect 14829 12696 14841 12699
rect 14332 12668 14841 12696
rect 14332 12656 14338 12668
rect 14829 12665 14841 12668
rect 14875 12696 14887 12699
rect 15289 12699 15347 12705
rect 15289 12696 15301 12699
rect 14875 12668 15301 12696
rect 14875 12665 14887 12668
rect 14829 12659 14887 12665
rect 15289 12665 15301 12668
rect 15335 12665 15347 12699
rect 15289 12659 15347 12665
rect 15381 12699 15439 12705
rect 15381 12665 15393 12699
rect 15427 12696 15439 12699
rect 15841 12699 15899 12705
rect 15841 12696 15853 12699
rect 15427 12668 15853 12696
rect 15427 12665 15439 12668
rect 15381 12659 15439 12665
rect 15841 12665 15853 12668
rect 15887 12665 15899 12699
rect 15841 12659 15899 12665
rect 18080 12699 18138 12705
rect 18080 12665 18092 12699
rect 18126 12696 18138 12699
rect 18432 12696 18460 12724
rect 18984 12696 19012 12795
rect 20438 12792 20444 12844
rect 20496 12832 20502 12844
rect 20717 12835 20775 12841
rect 20717 12832 20729 12835
rect 20496 12804 20729 12832
rect 20496 12792 20502 12804
rect 20717 12801 20729 12804
rect 20763 12801 20775 12835
rect 20717 12795 20775 12801
rect 20898 12792 20904 12844
rect 20956 12832 20962 12844
rect 20993 12835 21051 12841
rect 20993 12832 21005 12835
rect 20956 12804 21005 12832
rect 20956 12792 20962 12804
rect 20993 12801 21005 12804
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12764 20131 12767
rect 21450 12764 21456 12776
rect 20119 12736 21456 12764
rect 20119 12733 20131 12736
rect 20073 12727 20131 12733
rect 21450 12724 21456 12736
rect 21508 12724 21514 12776
rect 18126 12668 19012 12696
rect 18126 12665 18138 12668
rect 18080 12659 18138 12665
rect 20438 12656 20444 12708
rect 20496 12696 20502 12708
rect 20625 12699 20683 12705
rect 20625 12696 20637 12699
rect 20496 12668 20637 12696
rect 20496 12656 20502 12668
rect 20625 12665 20637 12668
rect 20671 12665 20683 12699
rect 20625 12659 20683 12665
rect 13998 12628 14004 12640
rect 11287 12600 12434 12628
rect 13959 12600 14004 12628
rect 11287 12597 11299 12600
rect 11241 12591 11299 12597
rect 13998 12588 14004 12600
rect 14056 12588 14062 12640
rect 15746 12628 15752 12640
rect 15707 12600 15752 12628
rect 15746 12588 15752 12600
rect 15804 12588 15810 12640
rect 18417 12631 18475 12637
rect 18417 12597 18429 12631
rect 18463 12628 18475 12631
rect 18598 12628 18604 12640
rect 18463 12600 18604 12628
rect 18463 12597 18475 12600
rect 18417 12591 18475 12597
rect 18598 12588 18604 12600
rect 18656 12588 18662 12640
rect 18782 12628 18788 12640
rect 18743 12600 18788 12628
rect 18782 12588 18788 12600
rect 18840 12588 18846 12640
rect 18874 12588 18880 12640
rect 18932 12628 18938 12640
rect 18932 12600 18977 12628
rect 18932 12588 18938 12600
rect 19610 12588 19616 12640
rect 19668 12628 19674 12640
rect 19889 12631 19947 12637
rect 19889 12628 19901 12631
rect 19668 12600 19901 12628
rect 19668 12588 19674 12600
rect 19889 12597 19901 12600
rect 19935 12628 19947 12631
rect 20533 12631 20591 12637
rect 20533 12628 20545 12631
rect 19935 12600 20545 12628
rect 19935 12597 19947 12600
rect 19889 12591 19947 12597
rect 20533 12597 20545 12600
rect 20579 12628 20591 12631
rect 20806 12628 20812 12640
rect 20579 12600 20812 12628
rect 20579 12597 20591 12600
rect 20533 12591 20591 12597
rect 20806 12588 20812 12600
rect 20864 12588 20870 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 2130 12424 2136 12436
rect 1627 12396 2136 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 2314 12384 2320 12436
rect 2372 12424 2378 12436
rect 2866 12424 2872 12436
rect 2372 12396 2872 12424
rect 2372 12384 2378 12396
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 3418 12384 3424 12436
rect 3476 12424 3482 12436
rect 3973 12427 4031 12433
rect 3973 12424 3985 12427
rect 3476 12396 3985 12424
rect 3476 12384 3482 12396
rect 3973 12393 3985 12396
rect 4019 12393 4031 12427
rect 3973 12387 4031 12393
rect 4433 12427 4491 12433
rect 4433 12393 4445 12427
rect 4479 12424 4491 12427
rect 4706 12424 4712 12436
rect 4479 12396 4712 12424
rect 4479 12393 4491 12396
rect 4433 12387 4491 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 8297 12427 8355 12433
rect 8297 12393 8309 12427
rect 8343 12424 8355 12427
rect 9766 12424 9772 12436
rect 8343 12396 9772 12424
rect 8343 12393 8355 12396
rect 8297 12387 8355 12393
rect 9766 12384 9772 12396
rect 9824 12424 9830 12436
rect 10042 12424 10048 12436
rect 9824 12396 10048 12424
rect 9824 12384 9830 12396
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 13814 12424 13820 12436
rect 11664 12396 13820 12424
rect 11664 12384 11670 12396
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 14369 12427 14427 12433
rect 14369 12424 14381 12427
rect 14056 12396 14381 12424
rect 14056 12384 14062 12396
rect 14369 12393 14381 12396
rect 14415 12393 14427 12427
rect 14369 12387 14427 12393
rect 17129 12427 17187 12433
rect 17129 12393 17141 12427
rect 17175 12424 17187 12427
rect 17681 12427 17739 12433
rect 17681 12424 17693 12427
rect 17175 12396 17693 12424
rect 17175 12393 17187 12396
rect 17129 12387 17187 12393
rect 17681 12393 17693 12396
rect 17727 12393 17739 12427
rect 17681 12387 17739 12393
rect 18509 12427 18567 12433
rect 18509 12393 18521 12427
rect 18555 12424 18567 12427
rect 18782 12424 18788 12436
rect 18555 12396 18788 12424
rect 18555 12393 18567 12396
rect 18509 12387 18567 12393
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 18877 12427 18935 12433
rect 18877 12393 18889 12427
rect 18923 12424 18935 12427
rect 19150 12424 19156 12436
rect 18923 12396 19156 12424
rect 18923 12393 18935 12396
rect 18877 12387 18935 12393
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 19610 12384 19616 12436
rect 19668 12424 19674 12436
rect 20165 12427 20223 12433
rect 19668 12396 20116 12424
rect 19668 12384 19674 12396
rect 1670 12316 1676 12368
rect 1728 12356 1734 12368
rect 11054 12356 11060 12368
rect 1728 12328 11060 12356
rect 1728 12316 1734 12328
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 14829 12359 14887 12365
rect 14829 12356 14841 12359
rect 14384 12328 14841 12356
rect 2682 12248 2688 12300
rect 2740 12297 2746 12300
rect 2740 12288 2752 12297
rect 2740 12260 2785 12288
rect 2740 12251 2752 12260
rect 2740 12248 2746 12251
rect 2866 12248 2872 12300
rect 2924 12288 2930 12300
rect 4338 12288 4344 12300
rect 2924 12260 3004 12288
rect 4299 12260 4344 12288
rect 2924 12248 2930 12260
rect 2976 12229 3004 12260
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 5166 12297 5172 12300
rect 5160 12288 5172 12297
rect 5127 12260 5172 12288
rect 5160 12251 5172 12260
rect 5166 12248 5172 12251
rect 5224 12248 5230 12300
rect 7173 12291 7231 12297
rect 7173 12288 7185 12291
rect 6288 12260 7185 12288
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3970 12220 3976 12232
rect 3007 12192 3976 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 3970 12180 3976 12192
rect 4028 12180 4034 12232
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 4632 12084 4660 12183
rect 4706 12180 4712 12232
rect 4764 12220 4770 12232
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4764 12192 4905 12220
rect 4764 12180 4770 12192
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 6288 12093 6316 12260
rect 7173 12257 7185 12260
rect 7219 12257 7231 12291
rect 7173 12251 7231 12257
rect 10042 12248 10048 12300
rect 10100 12288 10106 12300
rect 10330 12291 10388 12297
rect 10330 12288 10342 12291
rect 10100 12260 10342 12288
rect 10100 12248 10106 12260
rect 10330 12257 10342 12260
rect 10376 12257 10388 12291
rect 11698 12288 11704 12300
rect 11659 12260 11704 12288
rect 10330 12251 10388 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 11957 12291 12015 12297
rect 11957 12288 11969 12291
rect 11808 12260 11969 12288
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 6917 12223 6975 12229
rect 6917 12220 6929 12223
rect 6512 12192 6929 12220
rect 6512 12180 6518 12192
rect 6917 12189 6929 12192
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 9306 12180 9312 12232
rect 9364 12220 9370 12232
rect 9582 12220 9588 12232
rect 9364 12192 9588 12220
rect 9364 12180 9370 12192
rect 9582 12180 9588 12192
rect 9640 12180 9646 12232
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 10870 12220 10876 12232
rect 10643 12192 10876 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 11808 12220 11836 12260
rect 11957 12257 11969 12260
rect 12003 12257 12015 12291
rect 14384 12288 14412 12328
rect 14829 12325 14841 12328
rect 14875 12325 14887 12359
rect 14829 12319 14887 12325
rect 17221 12359 17279 12365
rect 17221 12325 17233 12359
rect 17267 12356 17279 12359
rect 18598 12356 18604 12368
rect 17267 12328 18604 12356
rect 17267 12325 17279 12328
rect 17221 12319 17279 12325
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 18690 12316 18696 12368
rect 18748 12356 18754 12368
rect 19705 12359 19763 12365
rect 18748 12328 19334 12356
rect 18748 12316 18754 12328
rect 11957 12251 12015 12257
rect 12820 12260 14412 12288
rect 14737 12291 14795 12297
rect 12820 12220 12848 12260
rect 14737 12257 14749 12291
rect 14783 12288 14795 12291
rect 15102 12288 15108 12300
rect 14783 12260 15108 12288
rect 14783 12257 14795 12260
rect 14737 12251 14795 12257
rect 15102 12248 15108 12260
rect 15160 12248 15166 12300
rect 15657 12291 15715 12297
rect 15657 12257 15669 12291
rect 15703 12288 15715 12291
rect 16114 12288 16120 12300
rect 15703 12260 16120 12288
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 16114 12248 16120 12260
rect 16172 12288 16178 12300
rect 17862 12288 17868 12300
rect 16172 12260 17868 12288
rect 16172 12248 16178 12260
rect 17862 12248 17868 12260
rect 17920 12248 17926 12300
rect 18046 12288 18052 12300
rect 18007 12260 18052 12288
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 11664 12192 11836 12220
rect 12728 12192 12848 12220
rect 11664 12180 11670 12192
rect 7926 12112 7932 12164
rect 7984 12152 7990 12164
rect 7984 12124 9352 12152
rect 7984 12112 7990 12124
rect 6273 12087 6331 12093
rect 6273 12084 6285 12087
rect 4632 12056 6285 12084
rect 6273 12053 6285 12056
rect 6319 12053 6331 12087
rect 9214 12084 9220 12096
rect 9175 12056 9220 12084
rect 6273 12047 6331 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 9324 12084 9352 12124
rect 10778 12084 10784 12096
rect 9324 12056 10784 12084
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 12066 12044 12072 12096
rect 12124 12084 12130 12096
rect 12434 12084 12440 12096
rect 12124 12056 12440 12084
rect 12124 12044 12130 12056
rect 12434 12044 12440 12056
rect 12492 12084 12498 12096
rect 12728 12084 12756 12192
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14921 12223 14979 12229
rect 14921 12220 14933 12223
rect 13872 12192 14933 12220
rect 13872 12180 13878 12192
rect 14921 12189 14933 12192
rect 14967 12220 14979 12223
rect 15286 12220 15292 12232
rect 14967 12192 15292 12220
rect 14967 12189 14979 12192
rect 14921 12183 14979 12189
rect 15286 12180 15292 12192
rect 15344 12220 15350 12232
rect 15381 12223 15439 12229
rect 15381 12220 15393 12223
rect 15344 12192 15393 12220
rect 15344 12180 15350 12192
rect 15381 12189 15393 12192
rect 15427 12189 15439 12223
rect 15381 12183 15439 12189
rect 15565 12223 15623 12229
rect 15565 12189 15577 12223
rect 15611 12220 15623 12223
rect 16758 12220 16764 12232
rect 15611 12192 16764 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 16942 12220 16948 12232
rect 16903 12192 16948 12220
rect 16942 12180 16948 12192
rect 17000 12180 17006 12232
rect 18138 12220 18144 12232
rect 18099 12192 18144 12220
rect 18138 12180 18144 12192
rect 18196 12180 18202 12232
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12220 18383 12223
rect 18414 12220 18420 12232
rect 18371 12192 18420 12220
rect 18371 12189 18383 12192
rect 18325 12183 18383 12189
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 18690 12180 18696 12232
rect 18748 12220 18754 12232
rect 18969 12223 19027 12229
rect 18969 12220 18981 12223
rect 18748 12192 18981 12220
rect 18748 12180 18754 12192
rect 18969 12189 18981 12192
rect 19015 12189 19027 12223
rect 19150 12220 19156 12232
rect 19111 12192 19156 12220
rect 18969 12183 19027 12189
rect 19150 12180 19156 12192
rect 19208 12180 19214 12232
rect 19306 12220 19334 12328
rect 19705 12325 19717 12359
rect 19751 12356 19763 12359
rect 19978 12356 19984 12368
rect 19751 12328 19984 12356
rect 19751 12325 19763 12328
rect 19705 12319 19763 12325
rect 19978 12316 19984 12328
rect 20036 12316 20042 12368
rect 20088 12356 20116 12396
rect 20165 12393 20177 12427
rect 20211 12424 20223 12427
rect 20346 12424 20352 12436
rect 20211 12396 20352 12424
rect 20211 12393 20223 12396
rect 20165 12387 20223 12393
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 20993 12427 21051 12433
rect 20993 12424 21005 12427
rect 20456 12396 21005 12424
rect 20456 12356 20484 12396
rect 20993 12393 21005 12396
rect 21039 12393 21051 12427
rect 20993 12387 21051 12393
rect 20088 12328 20484 12356
rect 20533 12359 20591 12365
rect 20533 12325 20545 12359
rect 20579 12356 20591 12359
rect 20622 12356 20628 12368
rect 20579 12328 20628 12356
rect 20579 12325 20591 12328
rect 20533 12319 20591 12325
rect 20622 12316 20628 12328
rect 20680 12316 20686 12368
rect 20714 12316 20720 12368
rect 20772 12356 20778 12368
rect 21269 12359 21327 12365
rect 21269 12356 21281 12359
rect 20772 12328 21281 12356
rect 20772 12316 20778 12328
rect 21269 12325 21281 12328
rect 21315 12325 21327 12359
rect 21269 12319 21327 12325
rect 20346 12248 20352 12300
rect 20404 12288 20410 12300
rect 21174 12288 21180 12300
rect 20404 12260 21180 12288
rect 20404 12248 20410 12260
rect 21174 12248 21180 12260
rect 21232 12248 21238 12300
rect 21450 12288 21456 12300
rect 21411 12260 21456 12288
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 19306 12192 20637 12220
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 20717 12223 20775 12229
rect 20717 12189 20729 12223
rect 20763 12189 20775 12223
rect 20717 12183 20775 12189
rect 13722 12112 13728 12164
rect 13780 12152 13786 12164
rect 19702 12152 19708 12164
rect 13780 12124 19708 12152
rect 13780 12112 13786 12124
rect 19702 12112 19708 12124
rect 19760 12112 19766 12164
rect 19889 12155 19947 12161
rect 19889 12121 19901 12155
rect 19935 12152 19947 12155
rect 19935 12124 20484 12152
rect 19935 12121 19947 12124
rect 19889 12115 19947 12121
rect 12492 12056 12756 12084
rect 13081 12087 13139 12093
rect 12492 12044 12498 12056
rect 13081 12053 13093 12087
rect 13127 12084 13139 12087
rect 13814 12084 13820 12096
rect 13127 12056 13820 12084
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 13814 12044 13820 12056
rect 13872 12084 13878 12096
rect 14366 12084 14372 12096
rect 13872 12056 14372 12084
rect 13872 12044 13878 12056
rect 14366 12044 14372 12056
rect 14424 12084 14430 12096
rect 15838 12084 15844 12096
rect 14424 12056 15844 12084
rect 14424 12044 14430 12056
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 16022 12084 16028 12096
rect 15983 12056 16028 12084
rect 16022 12044 16028 12056
rect 16080 12044 16086 12096
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 17589 12087 17647 12093
rect 16172 12056 16217 12084
rect 16172 12044 16178 12056
rect 17589 12053 17601 12087
rect 17635 12084 17647 12087
rect 19058 12084 19064 12096
rect 17635 12056 19064 12084
rect 17635 12053 17647 12056
rect 17589 12047 17647 12053
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 20073 12087 20131 12093
rect 20073 12053 20085 12087
rect 20119 12084 20131 12087
rect 20346 12084 20352 12096
rect 20119 12056 20352 12084
rect 20119 12053 20131 12056
rect 20073 12047 20131 12053
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 20456 12084 20484 12124
rect 20530 12112 20536 12164
rect 20588 12152 20594 12164
rect 20732 12152 20760 12183
rect 20588 12124 20760 12152
rect 20588 12112 20594 12124
rect 21450 12084 21456 12096
rect 20456 12056 21456 12084
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 2682 11880 2688 11892
rect 1627 11852 2688 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2682 11840 2688 11852
rect 2740 11880 2746 11892
rect 2740 11852 3004 11880
rect 2740 11840 2746 11852
rect 2976 11744 3004 11852
rect 4890 11840 4896 11892
rect 4948 11880 4954 11892
rect 5442 11880 5448 11892
rect 4948 11852 5448 11880
rect 4948 11840 4954 11852
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 5994 11840 6000 11892
rect 6052 11880 6058 11892
rect 6270 11880 6276 11892
rect 6052 11852 6276 11880
rect 6052 11840 6058 11852
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 6546 11880 6552 11892
rect 6507 11852 6552 11880
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 13446 11880 13452 11892
rect 8444 11852 13452 11880
rect 8444 11840 8450 11852
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 14090 11880 14096 11892
rect 14051 11852 14096 11880
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15657 11883 15715 11889
rect 15657 11880 15669 11883
rect 15528 11852 15669 11880
rect 15528 11840 15534 11852
rect 15657 11849 15669 11852
rect 15703 11849 15715 11883
rect 15657 11843 15715 11849
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 15896 11852 16252 11880
rect 15896 11840 15902 11852
rect 3050 11772 3056 11824
rect 3108 11812 3114 11824
rect 3108 11784 3153 11812
rect 3108 11772 3114 11784
rect 5166 11772 5172 11824
rect 5224 11812 5230 11824
rect 5350 11812 5356 11824
rect 5224 11784 5356 11812
rect 5224 11772 5230 11784
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 6638 11812 6644 11824
rect 6104 11784 6644 11812
rect 3510 11744 3516 11756
rect 2976 11716 3516 11744
rect 3510 11704 3516 11716
rect 3568 11744 3574 11756
rect 3605 11747 3663 11753
rect 3605 11744 3617 11747
rect 3568 11716 3617 11744
rect 3568 11704 3574 11716
rect 3605 11713 3617 11716
rect 3651 11713 3663 11747
rect 3970 11744 3976 11756
rect 3931 11716 3976 11744
rect 3605 11707 3663 11713
rect 3970 11704 3976 11716
rect 4028 11704 4034 11756
rect 4982 11704 4988 11756
rect 5040 11744 5046 11756
rect 6104 11753 6132 11784
rect 6638 11772 6644 11784
rect 6696 11772 6702 11824
rect 7742 11772 7748 11824
rect 7800 11812 7806 11824
rect 8297 11815 8355 11821
rect 8297 11812 8309 11815
rect 7800 11784 8309 11812
rect 7800 11772 7806 11784
rect 8297 11781 8309 11784
rect 8343 11781 8355 11815
rect 8297 11775 8355 11781
rect 9232 11784 9996 11812
rect 9232 11756 9260 11784
rect 5905 11747 5963 11753
rect 5905 11744 5917 11747
rect 5040 11716 5917 11744
rect 5040 11704 5046 11716
rect 5905 11713 5917 11716
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 6089 11747 6147 11753
rect 6089 11713 6101 11747
rect 6135 11713 6147 11747
rect 6089 11707 6147 11713
rect 6546 11704 6552 11756
rect 6604 11744 6610 11756
rect 7101 11747 7159 11753
rect 7101 11744 7113 11747
rect 6604 11716 7113 11744
rect 6604 11704 6610 11716
rect 7101 11713 7113 11716
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 7374 11704 7380 11756
rect 7432 11744 7438 11756
rect 7926 11744 7932 11756
rect 7432 11716 7932 11744
rect 7432 11704 7438 11716
rect 7926 11704 7932 11716
rect 7984 11704 7990 11756
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11744 8171 11747
rect 8202 11744 8208 11756
rect 8159 11716 8208 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 9214 11744 9220 11756
rect 8312 11716 9220 11744
rect 2866 11636 2872 11688
rect 2924 11676 2930 11688
rect 2961 11679 3019 11685
rect 2961 11676 2973 11679
rect 2924 11648 2973 11676
rect 2924 11636 2930 11648
rect 2961 11645 2973 11648
rect 3007 11645 3019 11679
rect 2961 11639 3019 11645
rect 3234 11636 3240 11688
rect 3292 11676 3298 11688
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 3292 11648 3433 11676
rect 3292 11636 3298 11648
rect 3421 11645 3433 11648
rect 3467 11645 3479 11679
rect 8312 11676 8340 11716
rect 9214 11704 9220 11716
rect 9272 11704 9278 11756
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 9968 11753 9996 11784
rect 9861 11747 9919 11753
rect 9861 11744 9873 11747
rect 9732 11716 9873 11744
rect 9732 11704 9738 11716
rect 9861 11713 9873 11716
rect 9907 11713 9919 11747
rect 9861 11707 9919 11713
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 10686 11744 10692 11756
rect 10647 11716 10692 11744
rect 9953 11707 10011 11713
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 11974 11744 11980 11756
rect 10836 11716 10881 11744
rect 11935 11716 11980 11744
rect 10836 11704 10842 11716
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 14108 11744 14136 11840
rect 15565 11815 15623 11821
rect 15565 11781 15577 11815
rect 15611 11781 15623 11815
rect 15565 11775 15623 11781
rect 14108 11716 14320 11744
rect 8478 11676 8484 11688
rect 3421 11639 3479 11645
rect 4172 11648 8340 11676
rect 8439 11648 8484 11676
rect 2406 11568 2412 11620
rect 2464 11608 2470 11620
rect 2716 11611 2774 11617
rect 2716 11608 2728 11611
rect 2464 11580 2728 11608
rect 2464 11568 2470 11580
rect 2716 11577 2728 11580
rect 2762 11608 2774 11611
rect 4172 11608 4200 11648
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11676 9367 11679
rect 10502 11676 10508 11688
rect 9355 11648 10508 11676
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 10502 11636 10508 11648
rect 10560 11676 10566 11688
rect 10873 11679 10931 11685
rect 10873 11676 10885 11679
rect 10560 11648 10885 11676
rect 10560 11636 10566 11648
rect 10873 11645 10885 11648
rect 10919 11645 10931 11679
rect 10873 11639 10931 11645
rect 11698 11636 11704 11688
rect 11756 11676 11762 11688
rect 12713 11679 12771 11685
rect 12713 11676 12725 11679
rect 11756 11648 12725 11676
rect 11756 11636 11762 11648
rect 12713 11645 12725 11648
rect 12759 11645 12771 11679
rect 12713 11639 12771 11645
rect 12980 11679 13038 11685
rect 12980 11645 12992 11679
rect 13026 11676 13038 11679
rect 13814 11676 13820 11688
rect 13026 11648 13820 11676
rect 13026 11645 13038 11648
rect 12980 11639 13038 11645
rect 2762 11580 4200 11608
rect 4240 11611 4298 11617
rect 2762 11577 2774 11580
rect 2716 11571 2774 11577
rect 4240 11577 4252 11611
rect 4286 11608 4298 11611
rect 4430 11608 4436 11620
rect 4286 11580 4436 11608
rect 4286 11577 4298 11580
rect 4240 11571 4298 11577
rect 4430 11568 4436 11580
rect 4488 11568 4494 11620
rect 9769 11611 9827 11617
rect 5184 11580 9444 11608
rect 1394 11540 1400 11552
rect 1355 11512 1400 11540
rect 1394 11500 1400 11512
rect 1452 11500 1458 11552
rect 3513 11543 3571 11549
rect 3513 11509 3525 11543
rect 3559 11540 3571 11543
rect 5184 11540 5212 11580
rect 3559 11512 5212 11540
rect 3559 11509 3571 11512
rect 3513 11503 3571 11509
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 5810 11540 5816 11552
rect 5500 11512 5545 11540
rect 5771 11512 5816 11540
rect 5500 11500 5506 11512
rect 5810 11500 5816 11512
rect 5868 11500 5874 11552
rect 6914 11540 6920 11552
rect 6875 11512 6920 11540
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 9416 11549 9444 11580
rect 9769 11577 9781 11611
rect 9815 11608 9827 11611
rect 12434 11608 12440 11620
rect 9815 11580 12440 11608
rect 9815 11577 9827 11580
rect 9769 11571 9827 11577
rect 12434 11568 12440 11580
rect 12492 11568 12498 11620
rect 12728 11608 12756 11639
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11645 14243 11679
rect 14292 11676 14320 11716
rect 14441 11679 14499 11685
rect 14441 11676 14453 11679
rect 14292 11648 14453 11676
rect 14185 11639 14243 11645
rect 14441 11645 14453 11648
rect 14487 11645 14499 11679
rect 15580 11676 15608 11775
rect 16022 11772 16028 11824
rect 16080 11812 16086 11824
rect 16080 11784 16160 11812
rect 16080 11772 16086 11784
rect 16132 11753 16160 11784
rect 16224 11753 16252 11852
rect 16758 11840 16764 11892
rect 16816 11880 16822 11892
rect 18325 11883 18383 11889
rect 16816 11852 17908 11880
rect 16816 11840 16822 11852
rect 17880 11812 17908 11852
rect 18325 11849 18337 11883
rect 18371 11880 18383 11883
rect 18598 11880 18604 11892
rect 18371 11852 18604 11880
rect 18371 11849 18383 11852
rect 18325 11843 18383 11849
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 20349 11883 20407 11889
rect 20349 11880 20361 11883
rect 19576 11852 20361 11880
rect 19576 11840 19582 11852
rect 20349 11849 20361 11852
rect 20395 11849 20407 11883
rect 20349 11843 20407 11849
rect 20809 11883 20867 11889
rect 20809 11849 20821 11883
rect 20855 11880 20867 11883
rect 20990 11880 20996 11892
rect 20855 11852 20996 11880
rect 20855 11849 20867 11852
rect 20809 11843 20867 11849
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 21361 11883 21419 11889
rect 21361 11849 21373 11883
rect 21407 11880 21419 11883
rect 21726 11880 21732 11892
rect 21407 11852 21732 11880
rect 21407 11849 21419 11852
rect 21361 11843 21419 11849
rect 21726 11840 21732 11852
rect 21784 11840 21790 11892
rect 18506 11812 18512 11824
rect 17880 11784 18512 11812
rect 18506 11772 18512 11784
rect 18564 11772 18570 11824
rect 19058 11772 19064 11824
rect 19116 11812 19122 11824
rect 20898 11812 20904 11824
rect 19116 11784 19288 11812
rect 19116 11772 19122 11784
rect 19260 11753 19288 11784
rect 19904 11784 20904 11812
rect 19904 11753 19932 11784
rect 20898 11772 20904 11784
rect 20956 11772 20962 11824
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 16209 11747 16267 11753
rect 16209 11713 16221 11747
rect 16255 11713 16267 11747
rect 16209 11707 16267 11713
rect 19245 11747 19303 11753
rect 19245 11713 19257 11747
rect 19291 11713 19303 11747
rect 19245 11707 19303 11713
rect 19889 11747 19947 11753
rect 19889 11713 19901 11747
rect 19935 11713 19947 11747
rect 19889 11707 19947 11713
rect 19978 11704 19984 11756
rect 20036 11744 20042 11756
rect 20036 11716 20081 11744
rect 20036 11704 20042 11716
rect 14441 11639 14499 11645
rect 14568 11648 15608 11676
rect 13078 11608 13084 11620
rect 12728 11580 13084 11608
rect 13078 11568 13084 11580
rect 13136 11608 13142 11620
rect 14200 11608 14228 11639
rect 13136 11580 14228 11608
rect 13136 11568 13142 11580
rect 14274 11568 14280 11620
rect 14332 11608 14338 11620
rect 14568 11608 14596 11648
rect 15746 11636 15752 11688
rect 15804 11676 15810 11688
rect 16025 11679 16083 11685
rect 16025 11676 16037 11679
rect 15804 11648 16037 11676
rect 15804 11636 15810 11648
rect 16025 11645 16037 11648
rect 16071 11645 16083 11679
rect 16025 11639 16083 11645
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 16942 11676 16948 11688
rect 16816 11648 16948 11676
rect 16816 11636 16822 11648
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 20533 11679 20591 11685
rect 20533 11676 20545 11679
rect 17052 11648 20545 11676
rect 17052 11608 17080 11648
rect 20533 11645 20545 11648
rect 20579 11645 20591 11679
rect 20990 11676 20996 11688
rect 20951 11648 20996 11676
rect 20533 11639 20591 11645
rect 20990 11636 20996 11648
rect 21048 11636 21054 11688
rect 21450 11676 21456 11688
rect 21411 11648 21456 11676
rect 21450 11636 21456 11648
rect 21508 11636 21514 11688
rect 14332 11580 14596 11608
rect 16960 11580 17080 11608
rect 17190 11611 17248 11617
rect 14332 11568 14338 11580
rect 7009 11543 7067 11549
rect 7009 11509 7021 11543
rect 7055 11540 7067 11543
rect 7469 11543 7527 11549
rect 7469 11540 7481 11543
rect 7055 11512 7481 11540
rect 7055 11509 7067 11512
rect 7009 11503 7067 11509
rect 7469 11509 7481 11512
rect 7515 11509 7527 11543
rect 7469 11503 7527 11509
rect 7837 11543 7895 11549
rect 7837 11509 7849 11543
rect 7883 11540 7895 11543
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 7883 11512 9321 11540
rect 7883 11509 7895 11512
rect 7837 11503 7895 11509
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 9309 11503 9367 11509
rect 9401 11543 9459 11549
rect 9401 11509 9413 11543
rect 9447 11509 9459 11543
rect 11238 11540 11244 11552
rect 11199 11512 11244 11540
rect 9401 11503 9459 11509
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 12158 11540 12164 11552
rect 12119 11512 12164 11540
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12253 11543 12311 11549
rect 12253 11509 12265 11543
rect 12299 11540 12311 11543
rect 12526 11540 12532 11552
rect 12299 11512 12532 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 12621 11543 12679 11549
rect 12621 11509 12633 11543
rect 12667 11540 12679 11543
rect 16960 11540 16988 11580
rect 17190 11577 17202 11611
rect 17236 11577 17248 11611
rect 17190 11571 17248 11577
rect 12667 11512 16988 11540
rect 12667 11509 12679 11512
rect 12621 11503 12679 11509
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 17205 11540 17233 11571
rect 17862 11568 17868 11620
rect 17920 11608 17926 11620
rect 18782 11608 18788 11620
rect 17920 11580 18788 11608
rect 17920 11568 17926 11580
rect 18782 11568 18788 11580
rect 18840 11568 18846 11620
rect 18969 11611 19027 11617
rect 18969 11577 18981 11611
rect 19015 11608 19027 11611
rect 20162 11608 20168 11620
rect 19015 11580 20168 11608
rect 19015 11577 19027 11580
rect 18969 11571 19027 11577
rect 20162 11568 20168 11580
rect 20220 11568 20226 11620
rect 20717 11611 20775 11617
rect 20717 11577 20729 11611
rect 20763 11608 20775 11611
rect 21542 11608 21548 11620
rect 20763 11580 21548 11608
rect 20763 11577 20775 11580
rect 20717 11571 20775 11577
rect 21542 11568 21548 11580
rect 21600 11568 21606 11620
rect 17092 11512 17233 11540
rect 17092 11500 17098 11512
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18601 11543 18659 11549
rect 18601 11540 18613 11543
rect 18104 11512 18613 11540
rect 18104 11500 18110 11512
rect 18601 11509 18613 11512
rect 18647 11509 18659 11543
rect 19058 11540 19064 11552
rect 19019 11512 19064 11540
rect 18601 11503 18659 11509
rect 19058 11500 19064 11512
rect 19116 11500 19122 11552
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 19392 11512 19441 11540
rect 19392 11500 19398 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19429 11503 19487 11509
rect 19797 11543 19855 11549
rect 19797 11509 19809 11543
rect 19843 11540 19855 11543
rect 20070 11540 20076 11552
rect 19843 11512 20076 11540
rect 19843 11509 19855 11512
rect 19797 11503 19855 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 21177 11543 21235 11549
rect 21177 11509 21189 11543
rect 21223 11540 21235 11543
rect 21450 11540 21456 11552
rect 21223 11512 21456 11540
rect 21223 11509 21235 11512
rect 21177 11503 21235 11509
rect 21450 11500 21456 11512
rect 21508 11500 21514 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 1670 11336 1676 11348
rect 1627 11308 1676 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 1946 11336 1952 11348
rect 1907 11308 1952 11336
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 3237 11339 3295 11345
rect 3237 11336 3249 11339
rect 2823 11308 3249 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 3237 11305 3249 11308
rect 3283 11305 3295 11339
rect 3237 11299 3295 11305
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 4709 11339 4767 11345
rect 4709 11336 4721 11339
rect 4396 11308 4721 11336
rect 4396 11296 4402 11308
rect 4709 11305 4721 11308
rect 4755 11305 4767 11339
rect 4709 11299 4767 11305
rect 4801 11339 4859 11345
rect 4801 11305 4813 11339
rect 4847 11336 4859 11339
rect 5074 11336 5080 11348
rect 4847 11308 5080 11336
rect 4847 11305 4859 11308
rect 4801 11299 4859 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 5629 11339 5687 11345
rect 5629 11336 5641 11339
rect 5307 11308 5641 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5629 11305 5641 11308
rect 5675 11305 5687 11339
rect 5629 11299 5687 11305
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 6089 11339 6147 11345
rect 6089 11336 6101 11339
rect 5776 11308 6101 11336
rect 5776 11296 5782 11308
rect 6089 11305 6101 11308
rect 6135 11305 6147 11339
rect 6089 11299 6147 11305
rect 6914 11296 6920 11348
rect 6972 11336 6978 11348
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 6972 11308 7297 11336
rect 6972 11296 6978 11308
rect 7285 11305 7297 11308
rect 7331 11305 7343 11339
rect 7285 11299 7343 11305
rect 7745 11339 7803 11345
rect 7745 11305 7757 11339
rect 7791 11336 7803 11339
rect 8386 11336 8392 11348
rect 7791 11308 8392 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 9674 11336 9680 11348
rect 9635 11308 9680 11336
rect 9674 11296 9680 11308
rect 9732 11336 9738 11348
rect 10594 11336 10600 11348
rect 9732 11308 10600 11336
rect 9732 11296 9738 11308
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 11790 11336 11796 11348
rect 10980 11308 11796 11336
rect 3142 11268 3148 11280
rect 1780 11240 3148 11268
rect 1780 11212 1808 11240
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 5169 11271 5227 11277
rect 5169 11237 5181 11271
rect 5215 11268 5227 11271
rect 5442 11268 5448 11280
rect 5215 11240 5448 11268
rect 5215 11237 5227 11240
rect 5169 11231 5227 11237
rect 5442 11228 5448 11240
rect 5500 11228 5506 11280
rect 7466 11228 7472 11280
rect 7524 11268 7530 11280
rect 7653 11271 7711 11277
rect 7653 11268 7665 11271
rect 7524 11240 7665 11268
rect 7524 11228 7530 11240
rect 7653 11237 7665 11240
rect 7699 11268 7711 11271
rect 8205 11271 8263 11277
rect 8205 11268 8217 11271
rect 7699 11240 8217 11268
rect 7699 11237 7711 11240
rect 7653 11231 7711 11237
rect 8205 11237 8217 11240
rect 8251 11268 8263 11271
rect 8251 11240 8800 11268
rect 8251 11237 8263 11240
rect 8205 11231 8263 11237
rect 1486 11200 1492 11212
rect 1447 11172 1492 11200
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 1762 11200 1768 11212
rect 1723 11172 1768 11200
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2409 11203 2467 11209
rect 2409 11169 2421 11203
rect 2455 11200 2467 11203
rect 2866 11200 2872 11212
rect 2455 11172 2872 11200
rect 2455 11169 2467 11172
rect 2409 11163 2467 11169
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 4338 11200 4344 11212
rect 4299 11172 4344 11200
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 5902 11160 5908 11212
rect 5960 11200 5966 11212
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 5960 11172 6009 11200
rect 5960 11160 5966 11172
rect 5997 11169 6009 11172
rect 6043 11169 6055 11203
rect 6546 11200 6552 11212
rect 5997 11163 6055 11169
rect 6104 11172 6552 11200
rect 2225 11135 2283 11141
rect 2225 11101 2237 11135
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 3326 11132 3332 11144
rect 2363 11104 2636 11132
rect 3287 11104 3332 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2240 11064 2268 11095
rect 2406 11064 2412 11076
rect 2240 11036 2412 11064
rect 2406 11024 2412 11036
rect 2464 11024 2470 11076
rect 2608 10996 2636 11104
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 3510 11132 3516 11144
rect 3471 11104 3516 11132
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4246 11132 4252 11144
rect 4207 11104 4252 11132
rect 4065 11095 4123 11101
rect 2869 11067 2927 11073
rect 2869 11033 2881 11067
rect 2915 11064 2927 11067
rect 2958 11064 2964 11076
rect 2915 11036 2964 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 2958 11024 2964 11036
rect 3016 11024 3022 11076
rect 4080 11064 4108 11095
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 4430 11092 4436 11144
rect 4488 11132 4494 11144
rect 5442 11132 5448 11144
rect 4488 11104 5448 11132
rect 4488 11092 4494 11104
rect 5442 11092 5448 11104
rect 5500 11132 5506 11144
rect 6104 11132 6132 11172
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 7834 11160 7840 11212
rect 7892 11200 7898 11212
rect 8665 11203 8723 11209
rect 8665 11200 8677 11203
rect 7892 11172 8677 11200
rect 7892 11160 7898 11172
rect 8665 11169 8677 11172
rect 8711 11169 8723 11203
rect 8772 11200 8800 11240
rect 8938 11228 8944 11280
rect 8996 11268 9002 11280
rect 9398 11268 9404 11280
rect 8996 11240 9404 11268
rect 8996 11228 9002 11240
rect 9398 11228 9404 11240
rect 9456 11268 9462 11280
rect 9585 11271 9643 11277
rect 9585 11268 9597 11271
rect 9456 11240 9597 11268
rect 9456 11228 9462 11240
rect 9585 11237 9597 11240
rect 9631 11237 9643 11271
rect 10980 11268 11008 11308
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 12158 11296 12164 11348
rect 12216 11336 12222 11348
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 12216 11308 12265 11336
rect 12216 11296 12222 11308
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 12253 11299 12311 11305
rect 12621 11339 12679 11345
rect 12621 11305 12633 11339
rect 12667 11336 12679 11339
rect 13081 11339 13139 11345
rect 13081 11336 13093 11339
rect 12667 11308 13093 11336
rect 12667 11305 12679 11308
rect 12621 11299 12679 11305
rect 13081 11305 13093 11308
rect 13127 11305 13139 11339
rect 13538 11336 13544 11348
rect 13499 11308 13544 11336
rect 13081 11299 13139 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 15378 11336 15384 11348
rect 13740 11308 15384 11336
rect 9585 11231 9643 11237
rect 9876 11240 11008 11268
rect 9876 11200 9904 11240
rect 11238 11228 11244 11280
rect 11296 11268 11302 11280
rect 12713 11271 12771 11277
rect 12713 11268 12725 11271
rect 11296 11240 12725 11268
rect 11296 11228 11302 11240
rect 12713 11237 12725 11240
rect 12759 11237 12771 11271
rect 12713 11231 12771 11237
rect 13449 11271 13507 11277
rect 13449 11237 13461 11271
rect 13495 11268 13507 11271
rect 13740 11268 13768 11308
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 15565 11339 15623 11345
rect 15565 11305 15577 11339
rect 15611 11336 15623 11339
rect 16850 11336 16856 11348
rect 15611 11308 16856 11336
rect 15611 11305 15623 11308
rect 15565 11299 15623 11305
rect 13495 11240 13768 11268
rect 13495 11237 13507 11240
rect 13449 11231 13507 11237
rect 13814 11228 13820 11280
rect 13872 11268 13878 11280
rect 15010 11268 15016 11280
rect 13872 11240 15016 11268
rect 13872 11228 13878 11240
rect 15010 11228 15016 11240
rect 15068 11228 15074 11280
rect 15488 11268 15516 11299
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 17034 11336 17040 11348
rect 16947 11308 17040 11336
rect 17034 11296 17040 11308
rect 17092 11336 17098 11348
rect 18601 11339 18659 11345
rect 17092 11308 17724 11336
rect 17092 11296 17098 11308
rect 15902 11271 15960 11277
rect 15902 11268 15914 11271
rect 15488 11240 15914 11268
rect 15902 11237 15914 11240
rect 15948 11237 15960 11271
rect 17589 11271 17647 11277
rect 17589 11268 17601 11271
rect 15902 11231 15960 11237
rect 16040 11240 17601 11268
rect 8772 11172 9904 11200
rect 8665 11163 8723 11169
rect 10686 11160 10692 11212
rect 10744 11200 10750 11212
rect 11048 11203 11106 11209
rect 11048 11200 11060 11203
rect 10744 11172 11060 11200
rect 10744 11160 10750 11172
rect 11048 11169 11060 11172
rect 11094 11200 11106 11203
rect 13906 11200 13912 11212
rect 11094 11172 13768 11200
rect 13867 11172 13912 11200
rect 11094 11169 11106 11172
rect 11048 11163 11106 11169
rect 5500 11104 6132 11132
rect 6273 11135 6331 11141
rect 5500 11092 5506 11104
rect 6273 11101 6285 11135
rect 6319 11132 6331 11135
rect 6638 11132 6644 11144
rect 6319 11104 6644 11132
rect 6319 11101 6331 11104
rect 6273 11095 6331 11101
rect 5350 11064 5356 11076
rect 4080 11036 5356 11064
rect 5350 11024 5356 11036
rect 5408 11024 5414 11076
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 6288 11064 6316 11095
rect 6638 11092 6644 11104
rect 6696 11132 6702 11144
rect 7101 11135 7159 11141
rect 7101 11132 7113 11135
rect 6696 11104 7113 11132
rect 6696 11092 6702 11104
rect 7101 11101 7113 11104
rect 7147 11132 7159 11135
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 7147 11104 7941 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7929 11101 7941 11104
rect 7975 11132 7987 11135
rect 8202 11132 8208 11144
rect 7975 11104 8208 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 9490 11092 9496 11144
rect 9548 11132 9554 11144
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9548 11104 9781 11132
rect 9548 11092 9554 11104
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 10778 11132 10784 11144
rect 10739 11104 10784 11132
rect 9769 11095 9827 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 13740 11141 13768 11172
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 14056 11172 14412 11200
rect 14056 11160 14062 11172
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12492 11104 12817 11132
rect 12492 11092 12498 11104
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 14274 11132 14280 11144
rect 13771 11104 14280 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14384 11132 14412 11172
rect 14550 11160 14556 11212
rect 14608 11200 14614 11212
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 14608 11172 14657 11200
rect 14608 11160 14614 11172
rect 14645 11169 14657 11172
rect 14691 11169 14703 11203
rect 16040 11200 16068 11240
rect 17589 11237 17601 11240
rect 17635 11237 17647 11271
rect 17696 11268 17724 11308
rect 18601 11305 18613 11339
rect 18647 11336 18659 11339
rect 18874 11336 18880 11348
rect 18647 11308 18880 11336
rect 18647 11305 18659 11308
rect 18601 11299 18659 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 19058 11296 19064 11348
rect 19116 11336 19122 11348
rect 19613 11339 19671 11345
rect 19613 11336 19625 11339
rect 19116 11308 19625 11336
rect 19116 11296 19122 11308
rect 19613 11305 19625 11308
rect 19659 11305 19671 11339
rect 19613 11299 19671 11305
rect 19702 11296 19708 11348
rect 19760 11336 19766 11348
rect 21361 11339 21419 11345
rect 21361 11336 21373 11339
rect 19760 11308 21373 11336
rect 19760 11296 19766 11308
rect 21361 11305 21373 11308
rect 21407 11305 21419 11339
rect 21361 11299 21419 11305
rect 19150 11268 19156 11280
rect 17696 11240 19156 11268
rect 17589 11231 17647 11237
rect 19150 11228 19156 11240
rect 19208 11228 19214 11280
rect 19242 11228 19248 11280
rect 19300 11228 19306 11280
rect 19518 11228 19524 11280
rect 19576 11268 19582 11280
rect 19981 11271 20039 11277
rect 19981 11268 19993 11271
rect 19576 11240 19993 11268
rect 19576 11228 19582 11240
rect 19981 11237 19993 11240
rect 20027 11237 20039 11271
rect 19981 11231 20039 11237
rect 20073 11271 20131 11277
rect 20073 11237 20085 11271
rect 20119 11268 20131 11271
rect 20530 11268 20536 11280
rect 20119 11240 20536 11268
rect 20119 11237 20131 11240
rect 20073 11231 20131 11237
rect 20530 11228 20536 11240
rect 20588 11228 20594 11280
rect 20901 11271 20959 11277
rect 20901 11237 20913 11271
rect 20947 11268 20959 11271
rect 21634 11268 21640 11280
rect 20947 11240 21640 11268
rect 20947 11237 20959 11240
rect 20901 11231 20959 11237
rect 21634 11228 21640 11240
rect 21692 11228 21698 11280
rect 14645 11163 14703 11169
rect 14936 11172 16068 11200
rect 17497 11203 17555 11209
rect 14826 11132 14832 11144
rect 14384 11104 14832 11132
rect 14826 11092 14832 11104
rect 14884 11092 14890 11144
rect 5592 11036 6316 11064
rect 5592 11024 5598 11036
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 8849 11067 8907 11073
rect 8849 11064 8861 11067
rect 8812 11036 8861 11064
rect 8812 11024 8818 11036
rect 8849 11033 8861 11036
rect 8895 11064 8907 11067
rect 10796 11064 10824 11092
rect 12342 11064 12348 11076
rect 8895 11036 10824 11064
rect 11716 11036 12348 11064
rect 8895 11033 8907 11036
rect 8849 11027 8907 11033
rect 4154 10996 4160 11008
rect 2608 10968 4160 10996
rect 4154 10956 4160 10968
rect 4212 10956 4218 11008
rect 6638 10996 6644 11008
rect 6599 10968 6644 10996
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 9217 10999 9275 11005
rect 9217 10965 9229 10999
rect 9263 10996 9275 10999
rect 9582 10996 9588 11008
rect 9263 10968 9588 10996
rect 9263 10965 9275 10968
rect 9217 10959 9275 10965
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 11146 10956 11152 11008
rect 11204 10996 11210 11008
rect 11716 10996 11744 11036
rect 12342 11024 12348 11036
rect 12400 11064 12406 11076
rect 14936 11064 14964 11172
rect 17497 11169 17509 11203
rect 17543 11200 17555 11203
rect 17862 11200 17868 11212
rect 17543 11172 17868 11200
rect 17543 11169 17555 11172
rect 17497 11163 17555 11169
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18049 11203 18107 11209
rect 18049 11200 18061 11203
rect 18012 11172 18061 11200
rect 18012 11160 18018 11172
rect 18049 11169 18061 11172
rect 18095 11169 18107 11203
rect 19061 11203 19119 11209
rect 19061 11200 19073 11203
rect 18049 11163 18107 11169
rect 18248 11172 19073 11200
rect 15010 11092 15016 11144
rect 15068 11132 15074 11144
rect 15565 11135 15623 11141
rect 15565 11132 15577 11135
rect 15068 11104 15577 11132
rect 15068 11092 15074 11104
rect 15565 11101 15577 11104
rect 15611 11101 15623 11135
rect 15565 11095 15623 11101
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11101 15715 11135
rect 15657 11095 15715 11101
rect 12400 11036 14964 11064
rect 12400 11024 12406 11036
rect 11204 10968 11744 10996
rect 12161 10999 12219 11005
rect 11204 10956 11210 10968
rect 12161 10965 12173 10999
rect 12207 10996 12219 10999
rect 12434 10996 12440 11008
rect 12207 10968 12440 10996
rect 12207 10965 12219 10968
rect 12161 10959 12219 10965
rect 12434 10956 12440 10968
rect 12492 10956 12498 11008
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13814 10996 13820 11008
rect 12952 10968 13820 10996
rect 12952 10956 12958 10968
rect 13814 10956 13820 10968
rect 13872 10956 13878 11008
rect 14826 10996 14832 11008
rect 14787 10968 14832 10996
rect 14826 10956 14832 10968
rect 14884 10956 14890 11008
rect 15672 10996 15700 11095
rect 16850 11092 16856 11144
rect 16908 11132 16914 11144
rect 17586 11132 17592 11144
rect 16908 11104 17592 11132
rect 16908 11092 16914 11104
rect 17586 11092 17592 11104
rect 17644 11132 17650 11144
rect 17681 11135 17739 11141
rect 17681 11132 17693 11135
rect 17644 11104 17693 11132
rect 17644 11092 17650 11104
rect 17681 11101 17693 11104
rect 17727 11101 17739 11135
rect 17681 11095 17739 11101
rect 17770 11092 17776 11144
rect 17828 11132 17834 11144
rect 18248 11141 18276 11172
rect 19061 11169 19073 11172
rect 19107 11169 19119 11203
rect 19260 11200 19288 11228
rect 19061 11163 19119 11169
rect 19168 11172 19288 11200
rect 19168 11141 19196 11172
rect 20346 11160 20352 11212
rect 20404 11200 20410 11212
rect 20809 11203 20867 11209
rect 20809 11200 20821 11203
rect 20404 11172 20821 11200
rect 20404 11160 20410 11172
rect 20809 11169 20821 11172
rect 20855 11169 20867 11203
rect 20809 11163 20867 11169
rect 21453 11203 21511 11209
rect 21453 11169 21465 11203
rect 21499 11200 21511 11203
rect 21542 11200 21548 11212
rect 21499 11172 21548 11200
rect 21499 11169 21511 11172
rect 21453 11163 21511 11169
rect 21542 11160 21548 11172
rect 21600 11160 21606 11212
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 17828 11104 18245 11132
rect 17828 11092 17834 11104
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 19153 11135 19211 11141
rect 19153 11132 19165 11135
rect 18233 11095 18291 11101
rect 18340 11104 19165 11132
rect 17957 11067 18015 11073
rect 17957 11033 17969 11067
rect 18003 11064 18015 11067
rect 18340 11064 18368 11104
rect 19153 11101 19165 11104
rect 19199 11101 19211 11135
rect 19153 11095 19211 11101
rect 19245 11135 19303 11141
rect 19245 11101 19257 11135
rect 19291 11132 19303 11135
rect 19978 11132 19984 11144
rect 19291 11104 19984 11132
rect 19291 11101 19303 11104
rect 19245 11095 19303 11101
rect 18690 11064 18696 11076
rect 18003 11036 18368 11064
rect 18651 11036 18696 11064
rect 18003 11033 18015 11036
rect 17957 11027 18015 11033
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 19260 11064 19288 11095
rect 19978 11092 19984 11104
rect 20036 11132 20042 11144
rect 20165 11135 20223 11141
rect 20165 11132 20177 11135
rect 20036 11104 20177 11132
rect 20036 11092 20042 11104
rect 20165 11101 20177 11104
rect 20211 11132 20223 11135
rect 20714 11132 20720 11144
rect 20211 11104 20720 11132
rect 20211 11101 20223 11104
rect 20165 11095 20223 11101
rect 20714 11092 20720 11104
rect 20772 11132 20778 11144
rect 20993 11135 21051 11141
rect 20993 11132 21005 11135
rect 20772 11104 21005 11132
rect 20772 11092 20778 11104
rect 20993 11101 21005 11104
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 20898 11064 20904 11076
rect 18800 11036 19288 11064
rect 19637 11036 20904 11064
rect 16758 10996 16764 11008
rect 15672 10968 16764 10996
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 17126 10956 17132 11008
rect 17184 10996 17190 11008
rect 17184 10968 17229 10996
rect 17184 10956 17190 10968
rect 17586 10956 17592 11008
rect 17644 10996 17650 11008
rect 18800 10996 18828 11036
rect 17644 10968 18828 10996
rect 17644 10956 17650 10968
rect 18874 10956 18880 11008
rect 18932 10996 18938 11008
rect 19637 10996 19665 11036
rect 20898 11024 20904 11036
rect 20956 11064 20962 11076
rect 21910 11064 21916 11076
rect 20956 11036 21916 11064
rect 20956 11024 20962 11036
rect 21910 11024 21916 11036
rect 21968 11024 21974 11076
rect 18932 10968 19665 10996
rect 18932 10956 18938 10968
rect 19702 10956 19708 11008
rect 19760 10996 19766 11008
rect 20441 10999 20499 11005
rect 20441 10996 20453 10999
rect 19760 10968 20453 10996
rect 19760 10956 19766 10968
rect 20441 10965 20453 10968
rect 20487 10965 20499 10999
rect 20441 10959 20499 10965
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 2777 10795 2835 10801
rect 2777 10761 2789 10795
rect 2823 10792 2835 10795
rect 3326 10792 3332 10804
rect 2823 10764 3332 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 4246 10792 4252 10804
rect 4207 10764 4252 10792
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 4396 10764 5181 10792
rect 4396 10752 4402 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 5169 10755 5227 10761
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 6733 10795 6791 10801
rect 6733 10792 6745 10795
rect 5776 10764 6745 10792
rect 5776 10752 5782 10764
rect 6733 10761 6745 10764
rect 6779 10761 6791 10795
rect 6733 10755 6791 10761
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 7064 10764 7113 10792
rect 7064 10752 7070 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 7101 10755 7159 10761
rect 8294 10752 8300 10804
rect 8352 10792 8358 10804
rect 9122 10792 9128 10804
rect 8352 10764 9128 10792
rect 8352 10752 8358 10764
rect 9122 10752 9128 10764
rect 9180 10752 9186 10804
rect 11146 10792 11152 10804
rect 9968 10764 11152 10792
rect 3142 10724 3148 10736
rect 3103 10696 3148 10724
rect 3142 10684 3148 10696
rect 3200 10684 3206 10736
rect 3712 10696 5488 10724
rect 1486 10616 1492 10668
rect 1544 10656 1550 10668
rect 1765 10659 1823 10665
rect 1765 10656 1777 10659
rect 1544 10628 1777 10656
rect 1544 10616 1550 10628
rect 1765 10625 1777 10628
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10656 2283 10659
rect 2406 10656 2412 10668
rect 2271 10628 2412 10656
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 2866 10656 2872 10668
rect 2827 10628 2872 10656
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 3712 10665 3740 10696
rect 5460 10668 5488 10696
rect 3697 10659 3755 10665
rect 3697 10625 3709 10659
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 4706 10588 4712 10600
rect 2746 10560 4712 10588
rect 1394 10480 1400 10532
rect 1452 10520 1458 10532
rect 1489 10523 1547 10529
rect 1489 10520 1501 10523
rect 1452 10492 1501 10520
rect 1452 10480 1458 10492
rect 1489 10489 1501 10492
rect 1535 10489 1547 10523
rect 1670 10520 1676 10532
rect 1631 10492 1676 10520
rect 1489 10483 1547 10489
rect 1670 10480 1676 10492
rect 1728 10480 1734 10532
rect 2409 10523 2467 10529
rect 2409 10489 2421 10523
rect 2455 10520 2467 10523
rect 2746 10520 2774 10560
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 5000 10588 5028 10619
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 5721 10659 5779 10665
rect 5721 10656 5733 10659
rect 5500 10628 5733 10656
rect 5500 10616 5506 10628
rect 5721 10625 5733 10628
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 9968 10665 9996 10764
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 11698 10792 11704 10804
rect 11611 10764 11704 10792
rect 11698 10752 11704 10764
rect 11756 10792 11762 10804
rect 11974 10792 11980 10804
rect 11756 10764 11980 10792
rect 11756 10752 11762 10764
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 17218 10792 17224 10804
rect 12176 10764 17224 10792
rect 10134 10684 10140 10736
rect 10192 10724 10198 10736
rect 10410 10724 10416 10736
rect 10192 10696 10416 10724
rect 10192 10684 10198 10696
rect 10410 10684 10416 10696
rect 10468 10724 10474 10736
rect 11057 10727 11115 10733
rect 10468 10696 10824 10724
rect 10468 10684 10474 10696
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7156 10628 7665 10656
rect 7156 10616 7162 10628
rect 7653 10625 7665 10628
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 9953 10659 10011 10665
rect 9953 10625 9965 10659
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10625 10103 10659
rect 10045 10619 10103 10625
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 5534 10588 5540 10600
rect 5000 10560 5540 10588
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 7742 10588 7748 10600
rect 6687 10560 7748 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 7742 10548 7748 10560
rect 7800 10548 7806 10600
rect 7929 10591 7987 10597
rect 7929 10557 7941 10591
rect 7975 10588 7987 10591
rect 8754 10588 8760 10600
rect 7975 10560 8760 10588
rect 7975 10557 7987 10560
rect 7929 10551 7987 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 9490 10588 9496 10600
rect 9324 10560 9496 10588
rect 2455 10492 2774 10520
rect 2455 10489 2467 10492
rect 2409 10483 2467 10489
rect 4154 10480 4160 10532
rect 4212 10520 4218 10532
rect 4798 10520 4804 10532
rect 4212 10492 4804 10520
rect 4212 10480 4218 10492
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 7374 10480 7380 10532
rect 7432 10520 7438 10532
rect 8174 10523 8232 10529
rect 8174 10520 8186 10523
rect 7432 10492 8186 10520
rect 7432 10480 7438 10492
rect 8174 10489 8186 10492
rect 8220 10520 8232 10523
rect 9324 10520 9352 10560
rect 9490 10548 9496 10560
rect 9548 10588 9554 10600
rect 10060 10588 10088 10619
rect 9548 10560 10088 10588
rect 9548 10548 9554 10560
rect 8220 10492 9352 10520
rect 8220 10489 8232 10492
rect 8174 10483 8232 10489
rect 9398 10480 9404 10532
rect 9456 10520 9462 10532
rect 10520 10520 10548 10619
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 10796 10656 10824 10696
rect 11057 10693 11069 10727
rect 11103 10724 11115 10727
rect 12176 10724 12204 10764
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 17681 10795 17739 10801
rect 17681 10761 17693 10795
rect 17727 10792 17739 10795
rect 18138 10792 18144 10804
rect 17727 10764 18144 10792
rect 17727 10761 17739 10764
rect 17681 10755 17739 10761
rect 18138 10752 18144 10764
rect 18196 10752 18202 10804
rect 18509 10795 18567 10801
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 18966 10792 18972 10804
rect 18555 10764 18972 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 18966 10752 18972 10764
rect 19024 10752 19030 10804
rect 19058 10752 19064 10804
rect 19116 10792 19122 10804
rect 20162 10792 20168 10804
rect 19116 10764 19932 10792
rect 20123 10764 20168 10792
rect 19116 10752 19122 10764
rect 11103 10696 12204 10724
rect 11103 10693 11115 10696
rect 11057 10687 11115 10693
rect 13078 10684 13084 10736
rect 13136 10724 13142 10736
rect 13449 10727 13507 10733
rect 13449 10724 13461 10727
rect 13136 10696 13461 10724
rect 13136 10684 13142 10696
rect 13449 10693 13461 10696
rect 13495 10693 13507 10727
rect 13449 10687 13507 10693
rect 19702 10684 19708 10736
rect 19760 10724 19766 10736
rect 19760 10696 19840 10724
rect 19760 10684 19766 10696
rect 14274 10656 14280 10668
rect 10652 10628 10697 10656
rect 10796 10628 11284 10656
rect 14235 10628 14280 10656
rect 10652 10616 10658 10628
rect 11256 10597 11284 10628
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 15470 10656 15476 10668
rect 14752 10628 15476 10656
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10588 11299 10591
rect 12342 10588 12348 10600
rect 11287 10560 12348 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12814 10591 12872 10597
rect 12814 10588 12826 10591
rect 12492 10560 12826 10588
rect 12492 10548 12498 10560
rect 12814 10557 12826 10560
rect 12860 10557 12872 10591
rect 13078 10588 13084 10600
rect 13039 10560 13084 10588
rect 12814 10551 12872 10557
rect 13078 10548 13084 10560
rect 13136 10548 13142 10600
rect 13633 10591 13691 10597
rect 13633 10557 13645 10591
rect 13679 10588 13691 10591
rect 13998 10588 14004 10600
rect 13679 10560 14004 10588
rect 13679 10557 13691 10560
rect 13633 10551 13691 10557
rect 13998 10548 14004 10560
rect 14056 10548 14062 10600
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10588 14243 10591
rect 14752 10588 14780 10628
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 15838 10656 15844 10668
rect 15611 10628 15844 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 15838 10616 15844 10628
rect 15896 10656 15902 10668
rect 16301 10659 16359 10665
rect 16301 10656 16313 10659
rect 15896 10628 16313 10656
rect 15896 10616 15902 10628
rect 16301 10625 16313 10628
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 16390 10616 16396 10668
rect 16448 10656 16454 10668
rect 17034 10656 17040 10668
rect 16448 10628 16712 10656
rect 16995 10628 17040 10656
rect 16448 10616 16454 10628
rect 14231 10560 14780 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 14826 10548 14832 10600
rect 14884 10588 14890 10600
rect 16577 10591 16635 10597
rect 16577 10588 16589 10591
rect 14884 10560 16589 10588
rect 14884 10548 14890 10560
rect 16577 10557 16589 10560
rect 16623 10557 16635 10591
rect 16684 10588 16712 10628
rect 17034 10616 17040 10628
rect 17092 10616 17098 10668
rect 17218 10656 17224 10668
rect 17179 10628 17224 10656
rect 17218 10616 17224 10628
rect 17276 10616 17282 10668
rect 18874 10616 18880 10668
rect 18932 10616 18938 10668
rect 19150 10656 19156 10668
rect 19111 10628 19156 10656
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 19429 10659 19487 10665
rect 19429 10625 19441 10659
rect 19475 10625 19487 10659
rect 19429 10619 19487 10625
rect 16684 10560 17080 10588
rect 16577 10551 16635 10557
rect 12894 10520 12900 10532
rect 9456 10492 10088 10520
rect 10520 10492 12900 10520
rect 9456 10480 9462 10492
rect 2314 10452 2320 10464
rect 2275 10424 2320 10452
rect 2314 10412 2320 10424
rect 2372 10412 2378 10464
rect 3786 10452 3792 10464
rect 3747 10424 3792 10452
rect 3786 10412 3792 10424
rect 3844 10412 3850 10464
rect 3881 10455 3939 10461
rect 3881 10421 3893 10455
rect 3927 10452 3939 10455
rect 4341 10455 4399 10461
rect 4341 10452 4353 10455
rect 3927 10424 4353 10452
rect 3927 10421 3939 10424
rect 3881 10415 3939 10421
rect 4341 10421 4353 10424
rect 4387 10421 4399 10455
rect 4341 10415 4399 10421
rect 4709 10455 4767 10461
rect 4709 10421 4721 10455
rect 4755 10452 4767 10455
rect 4890 10452 4896 10464
rect 4755 10424 4896 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5534 10452 5540 10464
rect 5495 10424 5540 10452
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 5626 10412 5632 10464
rect 5684 10452 5690 10464
rect 6454 10452 6460 10464
rect 5684 10424 5729 10452
rect 6415 10424 6460 10452
rect 5684 10412 5690 10424
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 7466 10452 7472 10464
rect 7427 10424 7472 10452
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 7561 10455 7619 10461
rect 7561 10421 7573 10455
rect 7607 10452 7619 10455
rect 9122 10452 9128 10464
rect 7607 10424 9128 10452
rect 7607 10421 7619 10424
rect 7561 10415 7619 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9306 10452 9312 10464
rect 9267 10424 9312 10452
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 9490 10452 9496 10464
rect 9451 10424 9496 10452
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 9861 10455 9919 10461
rect 9861 10421 9873 10455
rect 9907 10452 9919 10455
rect 9950 10452 9956 10464
rect 9907 10424 9956 10452
rect 9907 10421 9919 10424
rect 9861 10415 9919 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10060 10452 10088 10492
rect 12894 10480 12900 10492
rect 12952 10480 12958 10532
rect 13262 10480 13268 10532
rect 13320 10520 13326 10532
rect 15381 10523 15439 10529
rect 15381 10520 15393 10523
rect 13320 10492 15393 10520
rect 13320 10480 13326 10492
rect 15381 10489 15393 10492
rect 15427 10489 15439 10523
rect 15381 10483 15439 10489
rect 15470 10480 15476 10532
rect 15528 10520 15534 10532
rect 15930 10520 15936 10532
rect 15528 10492 15936 10520
rect 15528 10480 15534 10492
rect 15930 10480 15936 10492
rect 15988 10480 15994 10532
rect 16117 10523 16175 10529
rect 16117 10489 16129 10523
rect 16163 10520 16175 10523
rect 16942 10520 16948 10532
rect 16163 10492 16948 10520
rect 16163 10489 16175 10492
rect 16117 10483 16175 10489
rect 16942 10480 16948 10492
rect 17000 10480 17006 10532
rect 17052 10520 17080 10560
rect 17126 10548 17132 10600
rect 17184 10588 17190 10600
rect 17313 10591 17371 10597
rect 17313 10588 17325 10591
rect 17184 10560 17325 10588
rect 17184 10548 17190 10560
rect 17313 10557 17325 10560
rect 17359 10557 17371 10591
rect 18892 10588 18920 10616
rect 17313 10551 17371 10557
rect 17420 10560 18920 10588
rect 18969 10591 19027 10597
rect 17420 10520 17448 10560
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19334 10588 19340 10600
rect 19015 10560 19340 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 19334 10548 19340 10560
rect 19392 10548 19398 10600
rect 19444 10588 19472 10619
rect 19518 10588 19524 10600
rect 19444 10560 19524 10588
rect 19518 10548 19524 10560
rect 19576 10548 19582 10600
rect 19610 10548 19616 10600
rect 19668 10588 19674 10600
rect 19668 10560 19713 10588
rect 19668 10548 19674 10560
rect 17052 10492 17448 10520
rect 18877 10523 18935 10529
rect 18877 10489 18889 10523
rect 18923 10520 18935 10523
rect 19812 10520 19840 10696
rect 18923 10492 19840 10520
rect 19904 10520 19932 10764
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 20990 10792 20996 10804
rect 20951 10764 20996 10792
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 20073 10727 20131 10733
rect 20073 10693 20085 10727
rect 20119 10724 20131 10727
rect 21174 10724 21180 10736
rect 20119 10696 21180 10724
rect 20119 10693 20131 10696
rect 20073 10687 20131 10693
rect 21174 10684 21180 10696
rect 21232 10684 21238 10736
rect 20714 10656 20720 10668
rect 20675 10628 20720 10656
rect 20714 10616 20720 10628
rect 20772 10616 20778 10668
rect 20533 10591 20591 10597
rect 20533 10557 20545 10591
rect 20579 10588 20591 10591
rect 20622 10588 20628 10600
rect 20579 10560 20628 10588
rect 20579 10557 20591 10560
rect 20533 10551 20591 10557
rect 20622 10548 20628 10560
rect 20680 10548 20686 10600
rect 20898 10548 20904 10600
rect 20956 10588 20962 10600
rect 21177 10591 21235 10597
rect 21177 10588 21189 10591
rect 20956 10560 21189 10588
rect 20956 10548 20962 10560
rect 21177 10557 21189 10560
rect 21223 10557 21235 10591
rect 21177 10551 21235 10557
rect 21269 10523 21327 10529
rect 21269 10520 21281 10523
rect 19904 10492 21281 10520
rect 18923 10489 18935 10492
rect 18877 10483 18935 10489
rect 21269 10489 21281 10492
rect 21315 10489 21327 10523
rect 21450 10520 21456 10532
rect 21411 10492 21456 10520
rect 21269 10483 21327 10489
rect 21450 10480 21456 10492
rect 21508 10480 21514 10532
rect 10689 10455 10747 10461
rect 10689 10452 10701 10455
rect 10060 10424 10701 10452
rect 10689 10421 10701 10424
rect 10735 10421 10747 10455
rect 10689 10415 10747 10421
rect 12066 10412 12072 10464
rect 12124 10452 12130 10464
rect 13173 10455 13231 10461
rect 13173 10452 13185 10455
rect 12124 10424 13185 10452
rect 12124 10412 12130 10424
rect 13173 10421 13185 10424
rect 13219 10421 13231 10455
rect 13173 10415 13231 10421
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 13725 10455 13783 10461
rect 13725 10452 13737 10455
rect 13596 10424 13737 10452
rect 13596 10412 13602 10424
rect 13725 10421 13737 10424
rect 13771 10421 13783 10455
rect 13725 10415 13783 10421
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14090 10452 14096 10464
rect 13964 10424 14096 10452
rect 13964 10412 13970 10424
rect 14090 10412 14096 10424
rect 14148 10412 14154 10464
rect 14274 10412 14280 10464
rect 14332 10452 14338 10464
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 14332 10424 14933 10452
rect 14332 10412 14338 10424
rect 14921 10421 14933 10424
rect 14967 10421 14979 10455
rect 15286 10452 15292 10464
rect 15247 10424 15292 10452
rect 14921 10415 14979 10421
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 15746 10452 15752 10464
rect 15707 10424 15752 10452
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 16206 10452 16212 10464
rect 16167 10424 16212 10452
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16758 10452 16764 10464
rect 16671 10424 16764 10452
rect 16758 10412 16764 10424
rect 16816 10452 16822 10464
rect 17126 10452 17132 10464
rect 16816 10424 17132 10452
rect 16816 10412 16822 10424
rect 17126 10412 17132 10424
rect 17184 10412 17190 10464
rect 19702 10452 19708 10464
rect 19663 10424 19708 10452
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 20162 10412 20168 10464
rect 20220 10452 20226 10464
rect 20625 10455 20683 10461
rect 20625 10452 20637 10455
rect 20220 10424 20637 10452
rect 20220 10412 20226 10424
rect 20625 10421 20637 10424
rect 20671 10421 20683 10455
rect 20625 10415 20683 10421
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 1765 10251 1823 10257
rect 1765 10248 1777 10251
rect 1636 10220 1777 10248
rect 1636 10208 1642 10220
rect 1765 10217 1777 10220
rect 1811 10217 1823 10251
rect 2222 10248 2228 10260
rect 2183 10220 2228 10248
rect 1765 10211 1823 10217
rect 2222 10208 2228 10220
rect 2280 10208 2286 10260
rect 3786 10208 3792 10260
rect 3844 10248 3850 10260
rect 4525 10251 4583 10257
rect 4525 10248 4537 10251
rect 3844 10220 4537 10248
rect 3844 10208 3850 10220
rect 4525 10217 4537 10220
rect 4571 10217 4583 10251
rect 5442 10248 5448 10260
rect 5403 10220 5448 10248
rect 4525 10211 4583 10217
rect 5442 10208 5448 10220
rect 5500 10208 5506 10260
rect 7101 10251 7159 10257
rect 7101 10217 7113 10251
rect 7147 10248 7159 10251
rect 8386 10248 8392 10260
rect 7147 10220 8392 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 9122 10248 9128 10260
rect 9083 10220 9128 10248
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 9490 10248 9496 10260
rect 9451 10220 9496 10248
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 12437 10251 12495 10257
rect 9640 10220 9685 10248
rect 9784 10220 12296 10248
rect 9640 10208 9646 10220
rect 4433 10183 4491 10189
rect 4433 10149 4445 10183
rect 4479 10180 4491 10183
rect 5534 10180 5540 10192
rect 4479 10152 5540 10180
rect 4479 10149 4491 10152
rect 4433 10143 4491 10149
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 6638 10189 6644 10192
rect 6580 10183 6644 10189
rect 6580 10149 6592 10183
rect 6626 10149 6644 10183
rect 6580 10143 6644 10149
rect 6638 10140 6644 10143
rect 6696 10140 6702 10192
rect 9784 10180 9812 10220
rect 6748 10152 9812 10180
rect 11088 10183 11146 10189
rect 1486 10112 1492 10124
rect 1447 10084 1492 10112
rect 1486 10072 1492 10084
rect 1544 10072 1550 10124
rect 1946 10112 1952 10124
rect 1907 10084 1952 10112
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 2038 10072 2044 10124
rect 2096 10112 2102 10124
rect 2317 10115 2375 10121
rect 2317 10112 2329 10115
rect 2096 10084 2329 10112
rect 2096 10072 2102 10084
rect 2317 10081 2329 10084
rect 2363 10081 2375 10115
rect 2317 10075 2375 10081
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 4893 10115 4951 10121
rect 4893 10112 4905 10115
rect 4856 10084 4905 10112
rect 4856 10072 4862 10084
rect 4893 10081 4905 10084
rect 4939 10081 4951 10115
rect 6748 10112 6776 10152
rect 11088 10149 11100 10183
rect 11134 10180 11146 10183
rect 11698 10180 11704 10192
rect 11134 10152 11704 10180
rect 11134 10149 11146 10152
rect 11088 10143 11146 10149
rect 11698 10140 11704 10152
rect 11756 10140 11762 10192
rect 11977 10183 12035 10189
rect 11977 10149 11989 10183
rect 12023 10180 12035 10183
rect 12268 10180 12296 10220
rect 12437 10217 12449 10251
rect 12483 10248 12495 10251
rect 12526 10248 12532 10260
rect 12483 10220 12532 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 13262 10248 13268 10260
rect 12636 10220 13124 10248
rect 13223 10220 13268 10248
rect 12636 10180 12664 10220
rect 13096 10180 13124 10220
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13725 10251 13783 10257
rect 13725 10217 13737 10251
rect 13771 10248 13783 10251
rect 14274 10248 14280 10260
rect 13771 10220 14280 10248
rect 13771 10217 13783 10220
rect 13725 10211 13783 10217
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 14366 10208 14372 10260
rect 14424 10248 14430 10260
rect 14737 10251 14795 10257
rect 14737 10248 14749 10251
rect 14424 10220 14749 10248
rect 14424 10208 14430 10220
rect 14737 10217 14749 10220
rect 14783 10248 14795 10251
rect 14783 10220 15884 10248
rect 14783 10217 14795 10220
rect 14737 10211 14795 10217
rect 13817 10183 13875 10189
rect 12023 10152 12204 10180
rect 12268 10152 12664 10180
rect 12728 10152 13032 10180
rect 13096 10152 13308 10180
rect 12023 10149 12035 10152
rect 11977 10143 12035 10149
rect 4893 10075 4951 10081
rect 5828 10084 6776 10112
rect 8317 10115 8375 10121
rect 4982 10044 4988 10056
rect 4943 10016 4988 10044
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 5718 10044 5724 10056
rect 5215 10016 5724 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9976 1731 9979
rect 5828 9976 5856 10084
rect 8317 10081 8329 10115
rect 8363 10112 8375 10115
rect 8662 10112 8668 10124
rect 8363 10084 8668 10112
rect 8363 10081 8375 10084
rect 8317 10075 8375 10081
rect 8662 10072 8668 10084
rect 8720 10112 8726 10124
rect 12066 10112 12072 10124
rect 8720 10084 9352 10112
rect 12027 10084 12072 10112
rect 8720 10072 8726 10084
rect 9324 10056 9352 10084
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 12176 10112 12204 10152
rect 12728 10112 12756 10152
rect 12894 10112 12900 10124
rect 12176 10084 12756 10112
rect 12855 10084 12900 10112
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 8573 10047 8631 10053
rect 6871 10016 7604 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 1719 9948 5856 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 1854 9868 1860 9920
rect 1912 9908 1918 9920
rect 2501 9911 2559 9917
rect 2501 9908 2513 9911
rect 1912 9880 2513 9908
rect 1912 9868 1918 9880
rect 2501 9877 2513 9880
rect 2547 9877 2559 9911
rect 2501 9871 2559 9877
rect 7098 9868 7104 9920
rect 7156 9908 7162 9920
rect 7193 9911 7251 9917
rect 7193 9908 7205 9911
rect 7156 9880 7205 9908
rect 7156 9868 7162 9880
rect 7193 9877 7205 9880
rect 7239 9877 7251 9911
rect 7576 9908 7604 10016
rect 8573 10013 8585 10047
rect 8619 10044 8631 10047
rect 8754 10044 8760 10056
rect 8619 10016 8760 10044
rect 8619 10013 8631 10016
rect 8573 10007 8631 10013
rect 8588 9908 8616 10007
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 9306 10004 9312 10056
rect 9364 10044 9370 10056
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9364 10016 9689 10044
rect 9364 10004 9370 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10013 11943 10047
rect 12434 10044 12440 10056
rect 11885 10007 11943 10013
rect 12084 10016 12440 10044
rect 9582 9908 9588 9920
rect 7576 9880 9588 9908
rect 7193 9871 7251 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9953 9911 10011 9917
rect 9953 9908 9965 9911
rect 9732 9880 9965 9908
rect 9732 9868 9738 9880
rect 9953 9877 9965 9880
rect 9999 9877 10011 9911
rect 11348 9908 11376 10007
rect 11900 9976 11928 10007
rect 12084 9976 12112 10016
rect 12434 10004 12440 10016
rect 12492 10004 12498 10056
rect 12618 10044 12624 10056
rect 12579 10016 12624 10044
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 12802 10044 12808 10056
rect 12763 10016 12808 10044
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 13004 10044 13032 10152
rect 13280 10112 13308 10152
rect 13817 10149 13829 10183
rect 13863 10180 13875 10183
rect 15746 10180 15752 10192
rect 13863 10152 15752 10180
rect 13863 10149 13875 10152
rect 13817 10143 13875 10149
rect 15746 10140 15752 10152
rect 15804 10140 15810 10192
rect 15856 10180 15884 10220
rect 15930 10208 15936 10260
rect 15988 10248 15994 10260
rect 17586 10248 17592 10260
rect 15988 10220 17264 10248
rect 17547 10220 17592 10248
rect 15988 10208 15994 10220
rect 16454 10183 16512 10189
rect 16454 10180 16466 10183
rect 15856 10152 16466 10180
rect 16454 10149 16466 10152
rect 16500 10149 16512 10183
rect 16454 10143 16512 10149
rect 17126 10140 17132 10192
rect 17184 10140 17190 10192
rect 17236 10180 17264 10220
rect 17586 10208 17592 10220
rect 17644 10208 17650 10260
rect 19610 10248 19616 10260
rect 19571 10220 19616 10248
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 20993 10251 21051 10257
rect 19873 10220 20852 10248
rect 19334 10180 19340 10192
rect 17236 10152 19340 10180
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 14182 10112 14188 10124
rect 13280 10084 14188 10112
rect 14182 10072 14188 10084
rect 14240 10072 14246 10124
rect 15562 10112 15568 10124
rect 15120 10084 15568 10112
rect 13538 10044 13544 10056
rect 13004 10016 13544 10044
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10044 13691 10047
rect 14366 10044 14372 10056
rect 13679 10016 14372 10044
rect 13679 10013 13691 10016
rect 13633 10007 13691 10013
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 11900 9948 12112 9976
rect 12986 9936 12992 9988
rect 13044 9976 13050 9988
rect 15120 9976 15148 10084
rect 15562 10072 15568 10084
rect 15620 10072 15626 10124
rect 15838 10072 15844 10124
rect 15896 10121 15902 10124
rect 15896 10112 15908 10121
rect 16117 10115 16175 10121
rect 15896 10084 15941 10112
rect 15896 10075 15908 10084
rect 16117 10081 16129 10115
rect 16163 10112 16175 10115
rect 16209 10115 16267 10121
rect 16209 10112 16221 10115
rect 16163 10084 16221 10112
rect 16163 10081 16175 10084
rect 16117 10075 16175 10081
rect 16209 10081 16221 10084
rect 16255 10112 16267 10115
rect 17144 10112 17172 10140
rect 16255 10084 17172 10112
rect 16255 10081 16267 10084
rect 16209 10075 16267 10081
rect 15896 10072 15902 10075
rect 17218 10072 17224 10124
rect 17276 10112 17282 10124
rect 19873 10112 19901 10220
rect 20824 10180 20852 10220
rect 20993 10217 21005 10251
rect 21039 10248 21051 10251
rect 21266 10248 21272 10260
rect 21039 10220 21272 10248
rect 21039 10217 21051 10220
rect 20993 10211 21051 10217
rect 21266 10208 21272 10220
rect 21324 10208 21330 10260
rect 20824 10152 21312 10180
rect 19978 10112 19984 10124
rect 17276 10084 19901 10112
rect 19939 10084 19984 10112
rect 17276 10072 17282 10084
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 20806 10112 20812 10124
rect 20767 10084 20812 10112
rect 20806 10072 20812 10084
rect 20864 10072 20870 10124
rect 21284 10121 21312 10152
rect 21269 10115 21327 10121
rect 21269 10081 21281 10115
rect 21315 10081 21327 10115
rect 21450 10112 21456 10124
rect 21411 10084 21456 10112
rect 21269 10075 21327 10081
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 20073 10047 20131 10053
rect 20073 10044 20085 10047
rect 19392 10016 20085 10044
rect 19392 10004 19398 10016
rect 20073 10013 20085 10016
rect 20119 10013 20131 10047
rect 20073 10007 20131 10013
rect 20257 10047 20315 10053
rect 20257 10013 20269 10047
rect 20303 10044 20315 10047
rect 20438 10044 20444 10056
rect 20303 10016 20444 10044
rect 20303 10013 20315 10016
rect 20257 10007 20315 10013
rect 20438 10004 20444 10016
rect 20496 10004 20502 10056
rect 20717 10047 20775 10053
rect 20717 10013 20729 10047
rect 20763 10044 20775 10047
rect 21468 10044 21496 10072
rect 20763 10016 21496 10044
rect 20763 10013 20775 10016
rect 20717 10007 20775 10013
rect 20898 9976 20904 9988
rect 13044 9948 15148 9976
rect 17512 9948 20904 9976
rect 13044 9936 13050 9948
rect 13078 9908 13084 9920
rect 11348 9880 13084 9908
rect 9953 9871 10011 9877
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 14185 9911 14243 9917
rect 14185 9877 14197 9911
rect 14231 9908 14243 9911
rect 17512 9908 17540 9948
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 21177 9979 21235 9985
rect 21177 9945 21189 9979
rect 21223 9976 21235 9979
rect 21542 9976 21548 9988
rect 21223 9948 21548 9976
rect 21223 9945 21235 9948
rect 21177 9939 21235 9945
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 14231 9880 17540 9908
rect 14231 9877 14243 9880
rect 14185 9871 14243 9877
rect 18138 9868 18144 9920
rect 18196 9908 18202 9920
rect 20530 9908 20536 9920
rect 18196 9880 20536 9908
rect 18196 9868 18202 9880
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 1946 9664 1952 9716
rect 2004 9704 2010 9716
rect 2409 9707 2467 9713
rect 2409 9704 2421 9707
rect 2004 9676 2421 9704
rect 2004 9664 2010 9676
rect 2409 9673 2421 9676
rect 2455 9673 2467 9707
rect 2409 9667 2467 9673
rect 2884 9676 3832 9704
rect 2130 9636 2136 9648
rect 2091 9608 2136 9636
rect 2130 9596 2136 9608
rect 2188 9596 2194 9648
rect 2314 9596 2320 9648
rect 2372 9636 2378 9648
rect 2884 9636 2912 9676
rect 2372 9608 2912 9636
rect 2372 9596 2378 9608
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 1504 9540 2697 9568
rect 1504 9444 1532 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2832 9540 2881 9568
rect 2832 9528 2838 9540
rect 2869 9537 2881 9540
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 2317 9503 2375 9509
rect 2317 9500 2329 9503
rect 1636 9472 2329 9500
rect 1636 9460 1642 9472
rect 2317 9469 2329 9472
rect 2363 9469 2375 9503
rect 2590 9500 2596 9512
rect 2551 9472 2596 9500
rect 2317 9463 2375 9469
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 3142 9500 3148 9512
rect 2792 9472 3013 9500
rect 3103 9472 3148 9500
rect 1486 9432 1492 9444
rect 1447 9404 1492 9432
rect 1486 9392 1492 9404
rect 1544 9392 1550 9444
rect 1854 9432 1860 9444
rect 1815 9404 1860 9432
rect 1854 9392 1860 9404
rect 1912 9392 1918 9444
rect 2041 9435 2099 9441
rect 2041 9401 2053 9435
rect 2087 9432 2099 9435
rect 2792 9432 2820 9472
rect 2087 9404 2820 9432
rect 2087 9401 2099 9404
rect 2041 9395 2099 9401
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 2866 9364 2872 9376
rect 1627 9336 2872 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 2866 9324 2872 9336
rect 2924 9324 2930 9376
rect 2985 9364 3013 9472
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 3804 9500 3832 9676
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 4396 9676 4936 9704
rect 4396 9664 4402 9676
rect 4522 9568 4528 9580
rect 4483 9540 4528 9568
rect 4522 9528 4528 9540
rect 4580 9568 4586 9580
rect 4908 9577 4936 9676
rect 4982 9664 4988 9716
rect 5040 9704 5046 9716
rect 5040 9676 5764 9704
rect 5040 9664 5046 9676
rect 5353 9639 5411 9645
rect 5353 9605 5365 9639
rect 5399 9636 5411 9639
rect 5626 9636 5632 9648
rect 5399 9608 5632 9636
rect 5399 9605 5411 9608
rect 5353 9599 5411 9605
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 5736 9636 5764 9676
rect 7466 9664 7472 9716
rect 7524 9704 7530 9716
rect 8021 9707 8079 9713
rect 8021 9704 8033 9707
rect 7524 9676 8033 9704
rect 7524 9664 7530 9676
rect 8021 9673 8033 9676
rect 8067 9673 8079 9707
rect 8021 9667 8079 9673
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 13170 9704 13176 9716
rect 12584 9676 13176 9704
rect 12584 9664 12590 9676
rect 13170 9664 13176 9676
rect 13228 9704 13234 9716
rect 15102 9704 15108 9716
rect 13228 9676 15108 9704
rect 13228 9664 13234 9676
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 15473 9707 15531 9713
rect 15473 9704 15485 9707
rect 15344 9676 15485 9704
rect 15344 9664 15350 9676
rect 15473 9673 15485 9676
rect 15519 9673 15531 9707
rect 15473 9667 15531 9673
rect 15562 9664 15568 9716
rect 15620 9704 15626 9716
rect 15620 9676 17908 9704
rect 15620 9664 15626 9676
rect 5736 9608 5856 9636
rect 4755 9571 4813 9577
rect 4755 9568 4767 9571
rect 4580 9540 4767 9568
rect 4580 9528 4586 9540
rect 4755 9537 4767 9540
rect 4801 9537 4813 9571
rect 4755 9531 4813 9537
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9537 4951 9571
rect 5828 9568 5856 9608
rect 6730 9596 6736 9648
rect 6788 9636 6794 9648
rect 6788 9608 9352 9636
rect 6788 9596 6794 9608
rect 5828 9540 6040 9568
rect 4893 9531 4951 9537
rect 5902 9500 5908 9512
rect 3804 9472 5908 9500
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6012 9500 6040 9540
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 6362 9568 6368 9580
rect 6236 9540 6368 9568
rect 6236 9528 6242 9540
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 7374 9568 7380 9580
rect 7335 9540 7380 9568
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 8662 9568 8668 9580
rect 8623 9540 8668 9568
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 7469 9503 7527 9509
rect 7469 9500 7481 9503
rect 6012 9472 7481 9500
rect 7469 9469 7481 9472
rect 7515 9469 7527 9503
rect 8386 9500 8392 9512
rect 8347 9472 8392 9500
rect 7469 9463 7527 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 4246 9392 4252 9444
rect 4304 9432 4310 9444
rect 4706 9432 4712 9444
rect 4304 9404 4712 9432
rect 4304 9392 4310 9404
rect 4706 9392 4712 9404
rect 4764 9432 4770 9444
rect 4985 9435 5043 9441
rect 4985 9432 4997 9435
rect 4764 9404 4997 9432
rect 4764 9392 4770 9404
rect 4985 9401 4997 9404
rect 5031 9401 5043 9435
rect 7190 9432 7196 9444
rect 4985 9395 5043 9401
rect 5276 9404 7196 9432
rect 5276 9364 5304 9404
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 8481 9435 8539 9441
rect 8481 9432 8493 9435
rect 7944 9404 8493 9432
rect 7558 9364 7564 9376
rect 2985 9336 5304 9364
rect 7519 9336 7564 9364
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 7944 9373 7972 9404
rect 8481 9401 8493 9404
rect 8527 9401 8539 9435
rect 9324 9432 9352 9608
rect 9398 9596 9404 9648
rect 9456 9636 9462 9648
rect 11238 9636 11244 9648
rect 9456 9608 11244 9636
rect 9456 9596 9462 9608
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 14829 9639 14887 9645
rect 14829 9605 14841 9639
rect 14875 9636 14887 9639
rect 15838 9636 15844 9648
rect 14875 9608 15844 9636
rect 14875 9605 14887 9608
rect 14829 9599 14887 9605
rect 15838 9596 15844 9608
rect 15896 9596 15902 9648
rect 16666 9636 16672 9648
rect 16627 9608 16672 9636
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 16942 9636 16948 9648
rect 16903 9608 16948 9636
rect 16942 9596 16948 9608
rect 17000 9596 17006 9648
rect 9674 9528 9680 9580
rect 9732 9568 9738 9580
rect 10321 9571 10379 9577
rect 10321 9568 10333 9571
rect 9732 9540 10333 9568
rect 9732 9528 9738 9540
rect 10321 9537 10333 9540
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9568 10839 9571
rect 10827 9540 11836 9568
rect 10827 9537 10839 9540
rect 10781 9531 10839 9537
rect 10134 9500 10140 9512
rect 10095 9472 10140 9500
rect 10134 9460 10140 9472
rect 10192 9500 10198 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10192 9472 10977 9500
rect 10192 9460 10198 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 10229 9435 10287 9441
rect 10229 9432 10241 9435
rect 9324 9404 10241 9432
rect 8481 9395 8539 9401
rect 10229 9401 10241 9404
rect 10275 9432 10287 9435
rect 10873 9435 10931 9441
rect 10873 9432 10885 9435
rect 10275 9404 10885 9432
rect 10275 9401 10287 9404
rect 10229 9395 10287 9401
rect 10873 9401 10885 9404
rect 10919 9401 10931 9435
rect 11808 9432 11836 9540
rect 13078 9528 13084 9580
rect 13136 9568 13142 9580
rect 13262 9568 13268 9580
rect 13136 9540 13268 9568
rect 13136 9528 13142 9540
rect 13262 9528 13268 9540
rect 13320 9568 13326 9580
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 13320 9540 13461 9568
rect 13320 9528 13326 9540
rect 13449 9537 13461 9540
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 15470 9528 15476 9580
rect 15528 9568 15534 9580
rect 16117 9571 16175 9577
rect 16117 9568 16129 9571
rect 15528 9540 16129 9568
rect 15528 9528 15534 9540
rect 16117 9537 16129 9540
rect 16163 9568 16175 9571
rect 17497 9571 17555 9577
rect 17497 9568 17509 9571
rect 16163 9540 17509 9568
rect 16163 9537 16175 9540
rect 16117 9531 16175 9537
rect 17497 9537 17509 9540
rect 17543 9537 17555 9571
rect 17497 9531 17555 9537
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9500 11943 9503
rect 13096 9500 13124 9528
rect 13716 9503 13774 9509
rect 13716 9500 13728 9503
rect 11931 9472 13124 9500
rect 13648 9472 13728 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 12158 9441 12164 9444
rect 12152 9432 12164 9441
rect 11808 9404 12164 9432
rect 10873 9395 10931 9401
rect 12152 9395 12164 9404
rect 12158 9392 12164 9395
rect 12216 9392 12222 9444
rect 12618 9392 12624 9444
rect 12676 9432 12682 9444
rect 12676 9404 13308 9432
rect 12676 9392 12682 9404
rect 7929 9367 7987 9373
rect 7929 9333 7941 9367
rect 7975 9333 7987 9367
rect 9766 9364 9772 9376
rect 9727 9336 9772 9364
rect 7929 9327 7987 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 11333 9367 11391 9373
rect 11333 9333 11345 9367
rect 11379 9364 11391 9367
rect 12802 9364 12808 9376
rect 11379 9336 12808 9364
rect 11379 9333 11391 9336
rect 11333 9327 11391 9333
rect 12802 9324 12808 9336
rect 12860 9324 12866 9376
rect 13280 9373 13308 9404
rect 13265 9367 13323 9373
rect 13265 9333 13277 9367
rect 13311 9364 13323 9367
rect 13648 9364 13676 9472
rect 13716 9469 13728 9472
rect 13762 9500 13774 9503
rect 15488 9500 15516 9528
rect 13762 9472 15516 9500
rect 15841 9503 15899 9509
rect 13762 9469 13774 9472
rect 13716 9463 13774 9469
rect 15841 9469 15853 9503
rect 15887 9500 15899 9503
rect 16390 9500 16396 9512
rect 15887 9472 16396 9500
rect 15887 9469 15899 9472
rect 15841 9463 15899 9469
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 17405 9503 17463 9509
rect 17405 9500 17417 9503
rect 16724 9472 17417 9500
rect 16724 9460 16730 9472
rect 17405 9469 17417 9472
rect 17451 9469 17463 9503
rect 17880 9500 17908 9676
rect 19426 9664 19432 9716
rect 19484 9704 19490 9716
rect 19484 9676 20024 9704
rect 19484 9664 19490 9676
rect 19996 9645 20024 9676
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 20993 9707 21051 9713
rect 20993 9704 21005 9707
rect 20864 9676 21005 9704
rect 20864 9664 20870 9676
rect 20993 9673 21005 9676
rect 21039 9673 21051 9707
rect 20993 9667 21051 9673
rect 19889 9639 19947 9645
rect 19889 9605 19901 9639
rect 19935 9636 19947 9639
rect 19981 9639 20039 9645
rect 19981 9636 19993 9639
rect 19935 9608 19993 9636
rect 19935 9605 19947 9608
rect 19889 9599 19947 9605
rect 19981 9605 19993 9608
rect 20027 9605 20039 9639
rect 21082 9636 21088 9648
rect 19981 9599 20039 9605
rect 20548 9608 21088 9636
rect 20548 9568 20576 9608
rect 21082 9596 21088 9608
rect 21140 9596 21146 9648
rect 21358 9636 21364 9648
rect 21319 9608 21364 9636
rect 21358 9596 21364 9608
rect 21416 9596 21422 9648
rect 20714 9568 20720 9580
rect 19628 9540 20576 9568
rect 20675 9540 20720 9568
rect 19628 9500 19656 9540
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 17880 9472 19656 9500
rect 19705 9503 19763 9509
rect 17405 9463 17463 9469
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 19797 9503 19855 9509
rect 19797 9500 19809 9503
rect 19751 9472 19809 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 19797 9469 19809 9472
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9500 19947 9503
rect 20625 9503 20683 9509
rect 20625 9500 20637 9503
rect 19935 9472 20637 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 20625 9469 20637 9472
rect 20671 9469 20683 9503
rect 21174 9500 21180 9512
rect 21135 9472 21180 9500
rect 20625 9463 20683 9469
rect 21174 9460 21180 9472
rect 21232 9460 21238 9512
rect 21542 9500 21548 9512
rect 21503 9472 21548 9500
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 14550 9392 14556 9444
rect 14608 9432 14614 9444
rect 16485 9435 16543 9441
rect 14608 9404 16436 9432
rect 14608 9392 14614 9404
rect 13311 9336 13676 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 15378 9324 15384 9376
rect 15436 9364 15442 9376
rect 15933 9367 15991 9373
rect 15933 9364 15945 9367
rect 15436 9336 15945 9364
rect 15436 9324 15442 9336
rect 15933 9333 15945 9336
rect 15979 9364 15991 9367
rect 16298 9364 16304 9376
rect 15979 9336 16304 9364
rect 15979 9333 15991 9336
rect 15933 9327 15991 9333
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 16408 9364 16436 9404
rect 16485 9401 16497 9435
rect 16531 9432 16543 9435
rect 17313 9435 17371 9441
rect 17313 9432 17325 9435
rect 16531 9404 17325 9432
rect 16531 9401 16543 9404
rect 16485 9395 16543 9401
rect 17313 9401 17325 9404
rect 17359 9401 17371 9435
rect 17313 9395 17371 9401
rect 17586 9392 17592 9444
rect 17644 9432 17650 9444
rect 19426 9432 19432 9444
rect 19484 9441 19490 9444
rect 19484 9435 19518 9441
rect 17644 9404 18460 9432
rect 19370 9404 19432 9432
rect 17644 9392 17650 9404
rect 18138 9364 18144 9376
rect 16408 9336 18144 9364
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 18230 9324 18236 9376
rect 18288 9364 18294 9376
rect 18325 9367 18383 9373
rect 18325 9364 18337 9367
rect 18288 9336 18337 9364
rect 18288 9324 18294 9336
rect 18325 9333 18337 9336
rect 18371 9333 18383 9367
rect 18432 9364 18460 9404
rect 19426 9392 19432 9404
rect 19506 9432 19518 9435
rect 20438 9432 20444 9444
rect 19506 9404 20444 9432
rect 19506 9401 19518 9404
rect 19484 9395 19518 9401
rect 19484 9392 19490 9395
rect 20438 9392 20444 9404
rect 20496 9392 20502 9444
rect 19610 9364 19616 9376
rect 18432 9336 19616 9364
rect 18325 9327 18383 9333
rect 19610 9324 19616 9336
rect 19668 9364 19674 9376
rect 19797 9367 19855 9373
rect 19797 9364 19809 9367
rect 19668 9336 19809 9364
rect 19668 9324 19674 9336
rect 19797 9333 19809 9336
rect 19843 9333 19855 9367
rect 19797 9327 19855 9333
rect 20070 9324 20076 9376
rect 20128 9364 20134 9376
rect 20165 9367 20223 9373
rect 20165 9364 20177 9367
rect 20128 9336 20177 9364
rect 20128 9324 20134 9336
rect 20165 9333 20177 9336
rect 20211 9333 20223 9367
rect 20530 9364 20536 9376
rect 20491 9336 20536 9364
rect 20165 9327 20223 9333
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 2590 9120 2596 9172
rect 2648 9160 2654 9172
rect 3881 9163 3939 9169
rect 3881 9160 3893 9163
rect 2648 9132 3893 9160
rect 2648 9120 2654 9132
rect 3881 9129 3893 9132
rect 3927 9129 3939 9163
rect 3881 9123 3939 9129
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 5350 9160 5356 9172
rect 4764 9132 5356 9160
rect 4764 9120 4770 9132
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 5813 9163 5871 9169
rect 5813 9160 5825 9163
rect 5491 9132 5825 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 5813 9129 5825 9132
rect 5859 9129 5871 9163
rect 6178 9160 6184 9172
rect 6139 9132 6184 9160
rect 5813 9123 5871 9129
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 6273 9163 6331 9169
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 9309 9163 9367 9169
rect 9309 9160 9321 9163
rect 6319 9132 9321 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 9309 9129 9321 9132
rect 9355 9129 9367 9163
rect 9766 9160 9772 9172
rect 9727 9132 9772 9160
rect 9309 9123 9367 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 10413 9163 10471 9169
rect 10413 9129 10425 9163
rect 10459 9129 10471 9163
rect 10413 9123 10471 9129
rect 10873 9163 10931 9169
rect 10873 9129 10885 9163
rect 10919 9160 10931 9163
rect 11882 9160 11888 9172
rect 10919 9132 11888 9160
rect 10919 9129 10931 9132
rect 10873 9123 10931 9129
rect 1412 9064 4568 9092
rect 1412 9033 1440 9064
rect 1946 9033 1952 9036
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 1940 8987 1952 9033
rect 2004 9024 2010 9036
rect 2004 8996 2040 9024
rect 1946 8984 1952 8987
rect 2004 8984 2010 8996
rect 2406 8984 2412 9036
rect 2464 9024 2470 9036
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 2464 8996 4261 9024
rect 2464 8984 2470 8996
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 1688 8820 1716 8919
rect 3234 8916 3240 8968
rect 3292 8956 3298 8968
rect 4341 8959 4399 8965
rect 4341 8956 4353 8959
rect 3292 8928 4353 8956
rect 3292 8916 3298 8928
rect 4341 8925 4353 8928
rect 4387 8925 4399 8959
rect 4341 8919 4399 8925
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 3053 8891 3111 8897
rect 3053 8857 3065 8891
rect 3099 8888 3111 8891
rect 3142 8888 3148 8900
rect 3099 8860 3148 8888
rect 3099 8857 3111 8860
rect 3053 8851 3111 8857
rect 3142 8848 3148 8860
rect 3200 8888 3206 8900
rect 4448 8888 4476 8919
rect 3200 8860 4476 8888
rect 4540 8888 4568 9064
rect 5902 9052 5908 9104
rect 5960 9092 5966 9104
rect 7101 9095 7159 9101
rect 7101 9092 7113 9095
rect 5960 9064 7113 9092
rect 5960 9052 5966 9064
rect 7101 9061 7113 9064
rect 7147 9061 7159 9095
rect 7101 9055 7159 9061
rect 7190 9052 7196 9104
rect 7248 9092 7254 9104
rect 7248 9064 8524 9092
rect 7248 9052 7254 9064
rect 5353 9027 5411 9033
rect 5353 8993 5365 9027
rect 5399 9024 5411 9027
rect 5442 9024 5448 9036
rect 5399 8996 5448 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 8202 9024 8208 9036
rect 5776 8996 8208 9024
rect 5776 8984 5782 8996
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8386 9024 8392 9036
rect 8347 8996 8392 9024
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 8496 9024 8524 9064
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 9030 9092 9036 9104
rect 8628 9064 9036 9092
rect 8628 9052 8634 9064
rect 9030 9052 9036 9064
rect 9088 9092 9094 9104
rect 9125 9095 9183 9101
rect 9125 9092 9137 9095
rect 9088 9064 9137 9092
rect 9088 9052 9094 9064
rect 9125 9061 9137 9064
rect 9171 9061 9183 9095
rect 9125 9055 9183 9061
rect 9677 9095 9735 9101
rect 9677 9061 9689 9095
rect 9723 9092 9735 9095
rect 10428 9092 10456 9123
rect 11882 9120 11888 9132
rect 11940 9120 11946 9172
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 13357 9163 13415 9169
rect 13357 9160 13369 9163
rect 12952 9132 13369 9160
rect 12952 9120 12958 9132
rect 13357 9129 13369 9132
rect 13403 9129 13415 9163
rect 13357 9123 13415 9129
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 13504 9132 13737 9160
rect 13504 9120 13510 9132
rect 13725 9129 13737 9132
rect 13771 9160 13783 9163
rect 14461 9163 14519 9169
rect 14461 9160 14473 9163
rect 13771 9132 14473 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 14461 9129 14473 9132
rect 14507 9160 14519 9163
rect 14550 9160 14556 9172
rect 14507 9132 14556 9160
rect 14507 9129 14519 9132
rect 14461 9123 14519 9129
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 15565 9163 15623 9169
rect 15565 9129 15577 9163
rect 15611 9160 15623 9163
rect 15930 9160 15936 9172
rect 15611 9132 15936 9160
rect 15611 9129 15623 9132
rect 15565 9123 15623 9129
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 16025 9163 16083 9169
rect 16025 9129 16037 9163
rect 16071 9160 16083 9163
rect 16206 9160 16212 9172
rect 16071 9132 16212 9160
rect 16071 9129 16083 9132
rect 16025 9123 16083 9129
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 16298 9120 16304 9172
rect 16356 9160 16362 9172
rect 18969 9163 19027 9169
rect 16356 9132 18368 9160
rect 16356 9120 16362 9132
rect 11900 9092 11928 9120
rect 13817 9095 13875 9101
rect 13817 9092 13829 9095
rect 9723 9064 10456 9092
rect 10520 9064 10916 9092
rect 11900 9064 13829 9092
rect 9723 9061 9735 9064
rect 9677 9055 9735 9061
rect 10520 9024 10548 9064
rect 10778 9024 10784 9036
rect 8496 8996 10548 9024
rect 10739 8996 10784 9024
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 10888 9024 10916 9064
rect 13817 9061 13829 9064
rect 13863 9061 13875 9095
rect 18230 9092 18236 9104
rect 13817 9055 13875 9061
rect 15580 9064 18236 9092
rect 12710 9024 12716 9036
rect 10888 8996 12716 9024
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 13009 9027 13067 9033
rect 13009 8993 13021 9027
rect 13055 9024 13067 9027
rect 15580 9024 15608 9064
rect 18230 9052 18236 9064
rect 18288 9052 18294 9104
rect 13055 8996 15608 9024
rect 15657 9027 15715 9033
rect 13055 8993 13067 8996
rect 13009 8987 13067 8993
rect 15657 8993 15669 9027
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 17037 9027 17095 9033
rect 17037 8993 17049 9027
rect 17083 8993 17095 9027
rect 17037 8987 17095 8993
rect 5626 8956 5632 8968
rect 5587 8928 5632 8956
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 6365 8959 6423 8965
rect 6365 8956 6377 8959
rect 6144 8928 6377 8956
rect 6144 8916 6150 8928
rect 6365 8925 6377 8928
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8925 7251 8959
rect 7374 8956 7380 8968
rect 7335 8928 7380 8956
rect 7193 8919 7251 8925
rect 4985 8891 5043 8897
rect 4985 8888 4997 8891
rect 4540 8860 4997 8888
rect 3200 8848 3206 8860
rect 4985 8857 4997 8860
rect 5031 8857 5043 8891
rect 7208 8888 7236 8919
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 8478 8956 8484 8968
rect 8439 8928 8484 8956
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 8628 8928 8673 8956
rect 8628 8916 8634 8928
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 8812 8928 9873 8956
rect 8812 8916 8818 8928
rect 9861 8925 9873 8928
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8925 11023 8959
rect 11330 8956 11336 8968
rect 11291 8928 11336 8956
rect 10965 8919 11023 8925
rect 7653 8891 7711 8897
rect 7653 8888 7665 8891
rect 7208 8860 7665 8888
rect 4985 8851 5043 8857
rect 7653 8857 7665 8860
rect 7699 8888 7711 8891
rect 8662 8888 8668 8900
rect 7699 8860 8668 8888
rect 7699 8857 7711 8860
rect 7653 8851 7711 8857
rect 8662 8848 8668 8860
rect 8720 8848 8726 8900
rect 8941 8891 8999 8897
rect 8941 8857 8953 8891
rect 8987 8888 8999 8891
rect 9398 8888 9404 8900
rect 8987 8860 9404 8888
rect 8987 8857 8999 8860
rect 8941 8851 8999 8857
rect 2774 8820 2780 8832
rect 1688 8792 2780 8820
rect 2774 8780 2780 8792
rect 2832 8820 2838 8832
rect 3418 8820 3424 8832
rect 2832 8792 3424 8820
rect 2832 8780 2838 8792
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 5810 8780 5816 8832
rect 5868 8820 5874 8832
rect 6733 8823 6791 8829
rect 6733 8820 6745 8823
rect 5868 8792 6745 8820
rect 5868 8780 5874 8792
rect 6733 8789 6745 8792
rect 6779 8789 6791 8823
rect 6733 8783 6791 8789
rect 8021 8823 8079 8829
rect 8021 8789 8033 8823
rect 8067 8820 8079 8823
rect 8202 8820 8208 8832
rect 8067 8792 8208 8820
rect 8067 8789 8079 8792
rect 8021 8783 8079 8789
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 8956 8820 8984 8851
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 10980 8888 11008 8919
rect 11330 8916 11336 8928
rect 11388 8916 11394 8968
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 13909 8959 13967 8965
rect 13909 8925 13921 8959
rect 13955 8925 13967 8959
rect 15470 8956 15476 8968
rect 15431 8928 15476 8956
rect 13909 8919 13967 8925
rect 9732 8860 11008 8888
rect 9732 8848 9738 8860
rect 8444 8792 8984 8820
rect 8444 8780 8450 8792
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 9766 8820 9772 8832
rect 9088 8792 9772 8820
rect 9088 8780 9094 8792
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 11885 8823 11943 8829
rect 11885 8789 11897 8823
rect 11931 8820 11943 8823
rect 12158 8820 12164 8832
rect 11931 8792 12164 8820
rect 11931 8789 11943 8792
rect 11885 8783 11943 8789
rect 12158 8780 12164 8792
rect 12216 8820 12222 8832
rect 13924 8820 13952 8919
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 15672 8888 15700 8987
rect 16850 8956 16856 8968
rect 16811 8928 16856 8956
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 16945 8959 17003 8965
rect 16945 8925 16957 8959
rect 16991 8925 17003 8959
rect 16945 8919 17003 8925
rect 16960 8888 16988 8919
rect 15212 8860 15700 8888
rect 16316 8860 16988 8888
rect 12216 8792 13952 8820
rect 12216 8780 12222 8792
rect 14642 8780 14648 8832
rect 14700 8820 14706 8832
rect 15212 8829 15240 8860
rect 16316 8832 16344 8860
rect 15197 8823 15255 8829
rect 15197 8820 15209 8823
rect 14700 8792 15209 8820
rect 14700 8780 14706 8792
rect 15197 8789 15209 8792
rect 15243 8789 15255 8823
rect 16298 8820 16304 8832
rect 16259 8792 16304 8820
rect 15197 8783 15255 8789
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 16574 8820 16580 8832
rect 16535 8792 16580 8820
rect 16574 8780 16580 8792
rect 16632 8820 16638 8832
rect 17052 8820 17080 8987
rect 17126 8984 17132 9036
rect 17184 9024 17190 9036
rect 17586 9024 17592 9036
rect 17184 8996 17592 9024
rect 17184 8984 17190 8996
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 17856 9027 17914 9033
rect 17856 8993 17868 9027
rect 17902 9024 17914 9027
rect 18138 9024 18144 9036
rect 17902 8996 18144 9024
rect 17902 8993 17914 8996
rect 17856 8987 17914 8993
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 18340 9024 18368 9132
rect 18969 9129 18981 9163
rect 19015 9160 19027 9163
rect 19426 9160 19432 9172
rect 19015 9132 19432 9160
rect 19015 9129 19027 9132
rect 18969 9123 19027 9129
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 20162 9160 20168 9172
rect 19720 9132 20168 9160
rect 18414 9052 18420 9104
rect 18472 9092 18478 9104
rect 19518 9092 19524 9104
rect 18472 9064 19524 9092
rect 18472 9052 18478 9064
rect 19518 9052 19524 9064
rect 19576 9052 19582 9104
rect 19426 9024 19432 9036
rect 18340 8996 19432 9024
rect 19426 8984 19432 8996
rect 19484 9024 19490 9036
rect 19720 9024 19748 9132
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 20530 9120 20536 9172
rect 20588 9160 20594 9172
rect 20993 9163 21051 9169
rect 20993 9160 21005 9163
rect 20588 9132 21005 9160
rect 20588 9120 20594 9132
rect 20993 9129 21005 9132
rect 21039 9129 21051 9163
rect 20993 9123 21051 9129
rect 21082 9120 21088 9172
rect 21140 9160 21146 9172
rect 21361 9163 21419 9169
rect 21361 9160 21373 9163
rect 21140 9132 21373 9160
rect 21140 9120 21146 9132
rect 21361 9129 21373 9132
rect 21407 9129 21419 9163
rect 21361 9123 21419 9129
rect 19886 9092 19892 9104
rect 19847 9064 19892 9092
rect 19886 9052 19892 9064
rect 19944 9052 19950 9104
rect 20073 9095 20131 9101
rect 20073 9061 20085 9095
rect 20119 9092 20131 9095
rect 20119 9064 21496 9092
rect 20119 9061 20131 9064
rect 20073 9055 20131 9061
rect 19484 8996 19748 9024
rect 19904 9024 19932 9052
rect 21468 9036 21496 9064
rect 20533 9027 20591 9033
rect 20533 9024 20545 9027
rect 19904 8996 20545 9024
rect 19484 8984 19490 8996
rect 20533 8993 20545 8996
rect 20579 8993 20591 9027
rect 21450 9024 21456 9036
rect 21411 8996 21456 9024
rect 20533 8987 20591 8993
rect 21450 8984 21456 8996
rect 21508 8984 21514 9036
rect 19886 8916 19892 8968
rect 19944 8956 19950 8968
rect 20346 8956 20352 8968
rect 19944 8928 20352 8956
rect 19944 8916 19950 8928
rect 20346 8916 20352 8928
rect 20404 8956 20410 8968
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 20404 8928 20637 8956
rect 20404 8916 20410 8928
rect 20625 8925 20637 8928
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 20714 8916 20720 8968
rect 20772 8956 20778 8968
rect 20772 8928 20817 8956
rect 20772 8916 20778 8928
rect 18598 8848 18604 8900
rect 18656 8888 18662 8900
rect 20898 8888 20904 8900
rect 18656 8860 20904 8888
rect 18656 8848 18662 8860
rect 20898 8848 20904 8860
rect 20956 8848 20962 8900
rect 16632 8792 17080 8820
rect 17405 8823 17463 8829
rect 16632 8780 16638 8792
rect 17405 8789 17417 8823
rect 17451 8820 17463 8823
rect 18874 8820 18880 8832
rect 17451 8792 18880 8820
rect 17451 8789 17463 8792
rect 17405 8783 17463 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 20162 8820 20168 8832
rect 20123 8792 20168 8820
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 2406 8616 2412 8628
rect 2367 8588 2412 8616
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 2866 8616 2872 8628
rect 2700 8588 2872 8616
rect 2700 8548 2728 8588
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 3068 8588 3341 8616
rect 1780 8520 2728 8548
rect 1780 8412 1808 8520
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8480 1915 8483
rect 1946 8480 1952 8492
rect 1903 8452 1952 8480
rect 1903 8449 1915 8452
rect 1857 8443 1915 8449
rect 1946 8440 1952 8452
rect 2004 8480 2010 8492
rect 2593 8483 2651 8489
rect 2593 8480 2605 8483
rect 2004 8452 2605 8480
rect 2004 8440 2010 8452
rect 2593 8449 2605 8452
rect 2639 8449 2651 8483
rect 2774 8480 2780 8492
rect 2735 8452 2780 8480
rect 2593 8443 2651 8449
rect 2774 8440 2780 8452
rect 2832 8440 2838 8492
rect 2041 8415 2099 8421
rect 1780 8384 1992 8412
rect 1964 8353 1992 8384
rect 2041 8381 2053 8415
rect 2087 8412 2099 8415
rect 2869 8415 2927 8421
rect 2087 8384 2820 8412
rect 2087 8381 2099 8384
rect 2041 8375 2099 8381
rect 1949 8347 2007 8353
rect 1949 8313 1961 8347
rect 1995 8313 2007 8347
rect 2792 8344 2820 8384
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 3068 8412 3096 8588
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 3329 8579 3387 8585
rect 4157 8619 4215 8625
rect 4157 8585 4169 8619
rect 4203 8616 4215 8619
rect 5442 8616 5448 8628
rect 4203 8588 5304 8616
rect 5403 8588 5448 8616
rect 4203 8585 4215 8588
rect 4157 8579 4215 8585
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 3292 8520 3337 8548
rect 3292 8508 3298 8520
rect 3510 8440 3516 8492
rect 3568 8480 3574 8492
rect 3881 8483 3939 8489
rect 3881 8480 3893 8483
rect 3568 8452 3893 8480
rect 3568 8440 3574 8452
rect 3881 8449 3893 8452
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 2915 8384 3096 8412
rect 3789 8415 3847 8421
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 4172 8412 4200 8579
rect 4246 8508 4252 8560
rect 4304 8548 4310 8560
rect 4982 8548 4988 8560
rect 4304 8520 4988 8548
rect 4304 8508 4310 8520
rect 4982 8508 4988 8520
rect 5040 8508 5046 8560
rect 5276 8548 5304 8588
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 5592 8588 6132 8616
rect 5592 8576 5598 8588
rect 5718 8548 5724 8560
rect 5276 8520 5724 8548
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 6104 8548 6132 8588
rect 6178 8576 6184 8628
rect 6236 8616 6242 8628
rect 6273 8619 6331 8625
rect 6273 8616 6285 8619
rect 6236 8588 6285 8616
rect 6236 8576 6242 8588
rect 6273 8585 6285 8588
rect 6319 8585 6331 8619
rect 7929 8619 7987 8625
rect 6273 8579 6331 8585
rect 6380 8588 7512 8616
rect 6380 8548 6408 8588
rect 6104 8520 6408 8548
rect 7484 8548 7512 8588
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 8570 8616 8576 8628
rect 7975 8588 8576 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 8662 8576 8668 8628
rect 8720 8616 8726 8628
rect 12526 8616 12532 8628
rect 8720 8588 12532 8616
rect 8720 8576 8726 8588
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 16114 8616 16120 8628
rect 12768 8588 16120 8616
rect 12768 8576 12774 8588
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 19334 8616 19340 8628
rect 19295 8588 19340 8616
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 20036 8588 20085 8616
rect 20036 8576 20042 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 20990 8616 20996 8628
rect 20951 8588 20996 8616
rect 20073 8579 20131 8585
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8616 21419 8619
rect 21726 8616 21732 8628
rect 21407 8588 21732 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 21726 8576 21732 8588
rect 21784 8576 21790 8628
rect 8389 8551 8447 8557
rect 8389 8548 8401 8551
rect 7484 8520 8401 8548
rect 8389 8517 8401 8520
rect 8435 8548 8447 8551
rect 8754 8548 8760 8560
rect 8435 8520 8760 8548
rect 8435 8517 8447 8520
rect 8389 8511 8447 8517
rect 8754 8508 8760 8520
rect 8812 8508 8818 8560
rect 9766 8508 9772 8560
rect 9824 8548 9830 8560
rect 16298 8548 16304 8560
rect 9824 8520 16304 8548
rect 9824 8508 9830 8520
rect 16298 8508 16304 8520
rect 16356 8508 16362 8560
rect 18138 8508 18144 8560
rect 18196 8548 18202 8560
rect 18509 8551 18567 8557
rect 18509 8548 18521 8551
rect 18196 8520 18521 8548
rect 18196 8508 18202 8520
rect 18509 8517 18521 8520
rect 18555 8548 18567 8551
rect 18555 8520 20668 8548
rect 18555 8517 18567 8520
rect 18509 8511 18567 8517
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 4939 8452 5488 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 3835 8384 4200 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 5074 8372 5080 8424
rect 5132 8372 5138 8424
rect 5460 8412 5488 8452
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 5629 8483 5687 8489
rect 5629 8480 5641 8483
rect 5592 8452 5641 8480
rect 5592 8440 5598 8452
rect 5629 8449 5641 8452
rect 5675 8449 5687 8483
rect 5810 8480 5816 8492
rect 5771 8452 5816 8480
rect 5629 8443 5687 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 11238 8440 11244 8492
rect 11296 8480 11302 8492
rect 16574 8480 16580 8492
rect 11296 8452 16580 8480
rect 11296 8440 11302 8452
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 17126 8440 17132 8492
rect 17184 8480 17190 8492
rect 18708 8489 18736 8520
rect 20640 8492 20668 8520
rect 18693 8483 18751 8489
rect 17184 8452 17229 8480
rect 17184 8440 17190 8452
rect 18693 8449 18705 8483
rect 18739 8449 18751 8483
rect 18874 8480 18880 8492
rect 18835 8452 18880 8480
rect 18693 8443 18751 8449
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 19981 8483 20039 8489
rect 19981 8449 19993 8483
rect 20027 8480 20039 8483
rect 20346 8480 20352 8492
rect 20027 8452 20352 8480
rect 20027 8449 20039 8452
rect 19981 8443 20039 8449
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 20622 8480 20628 8492
rect 20583 8452 20628 8480
rect 20622 8440 20628 8452
rect 20680 8440 20686 8492
rect 6086 8412 6092 8424
rect 5460 8384 6092 8412
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 6178 8372 6184 8424
rect 6236 8412 6242 8424
rect 6454 8412 6460 8424
rect 6236 8384 6460 8412
rect 6236 8372 6242 8384
rect 6454 8372 6460 8384
rect 6512 8412 6518 8424
rect 6549 8415 6607 8421
rect 6549 8412 6561 8415
rect 6512 8384 6561 8412
rect 6512 8372 6518 8384
rect 6549 8381 6561 8384
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 9502 8415 9560 8421
rect 9502 8412 9514 8415
rect 7432 8384 9514 8412
rect 7432 8372 7438 8384
rect 9502 8381 9514 8384
rect 9548 8412 9560 8415
rect 9674 8412 9680 8424
rect 9548 8384 9680 8412
rect 9548 8381 9560 8384
rect 9502 8375 9560 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 19797 8415 19855 8421
rect 9824 8384 9869 8412
rect 9824 8372 9830 8384
rect 19797 8381 19809 8415
rect 19843 8412 19855 8415
rect 19843 8384 21496 8412
rect 19843 8381 19855 8384
rect 19797 8375 19855 8381
rect 3142 8344 3148 8356
rect 2792 8316 3148 8344
rect 1949 8307 2007 8313
rect 3142 8304 3148 8316
rect 3200 8304 3206 8356
rect 5092 8344 5120 8372
rect 21468 8356 21496 8384
rect 3712 8316 5120 8344
rect 1394 8276 1400 8288
rect 1355 8248 1400 8276
rect 1394 8236 1400 8248
rect 1452 8236 1458 8288
rect 2682 8236 2688 8288
rect 2740 8276 2746 8288
rect 3712 8285 3740 8316
rect 5626 8304 5632 8356
rect 5684 8344 5690 8356
rect 6822 8353 6828 8356
rect 6794 8347 6828 8353
rect 6794 8344 6806 8347
rect 5684 8316 6806 8344
rect 5684 8304 5690 8316
rect 6794 8313 6806 8316
rect 6880 8344 6886 8356
rect 6880 8316 6942 8344
rect 6794 8307 6828 8313
rect 6822 8304 6828 8307
rect 6880 8304 6886 8316
rect 7006 8304 7012 8356
rect 7064 8344 7070 8356
rect 14090 8344 14096 8356
rect 7064 8316 14096 8344
rect 7064 8304 7070 8316
rect 14090 8304 14096 8316
rect 14148 8304 14154 8356
rect 16850 8304 16856 8356
rect 16908 8344 16914 8356
rect 17374 8347 17432 8353
rect 17374 8344 17386 8347
rect 16908 8316 17386 8344
rect 16908 8304 16914 8316
rect 17374 8313 17386 8316
rect 17420 8344 17432 8347
rect 17678 8344 17684 8356
rect 17420 8316 17684 8344
rect 17420 8313 17432 8316
rect 17374 8307 17432 8313
rect 17678 8304 17684 8316
rect 17736 8304 17742 8356
rect 19613 8347 19671 8353
rect 19613 8313 19625 8347
rect 19659 8344 19671 8347
rect 21082 8344 21088 8356
rect 19659 8316 21088 8344
rect 19659 8313 19671 8316
rect 19613 8307 19671 8313
rect 21082 8304 21088 8316
rect 21140 8304 21146 8356
rect 21450 8344 21456 8356
rect 21411 8316 21456 8344
rect 21450 8304 21456 8316
rect 21508 8304 21514 8356
rect 3697 8279 3755 8285
rect 3697 8276 3709 8279
rect 2740 8248 3709 8276
rect 2740 8236 2746 8248
rect 3697 8245 3709 8248
rect 3743 8245 3755 8279
rect 3697 8239 3755 8245
rect 4890 8236 4896 8288
rect 4948 8276 4954 8288
rect 4985 8279 5043 8285
rect 4985 8276 4997 8279
rect 4948 8248 4997 8276
rect 4948 8236 4954 8248
rect 4985 8245 4997 8248
rect 5031 8245 5043 8279
rect 4985 8239 5043 8245
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5902 8276 5908 8288
rect 5132 8248 5177 8276
rect 5863 8248 5908 8276
rect 5132 8236 5138 8248
rect 5902 8236 5908 8248
rect 5960 8236 5966 8288
rect 18966 8276 18972 8288
rect 18927 8248 18972 8276
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 19978 8236 19984 8288
rect 20036 8276 20042 8288
rect 20441 8279 20499 8285
rect 20441 8276 20453 8279
rect 20036 8248 20453 8276
rect 20036 8236 20042 8248
rect 20441 8245 20453 8248
rect 20487 8245 20499 8279
rect 20441 8239 20499 8245
rect 20530 8236 20536 8288
rect 20588 8276 20594 8288
rect 20588 8248 20633 8276
rect 20588 8236 20594 8248
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2041 8075 2099 8081
rect 2041 8072 2053 8075
rect 2004 8044 2053 8072
rect 2004 8032 2010 8044
rect 2041 8041 2053 8044
rect 2087 8041 2099 8075
rect 15194 8072 15200 8084
rect 2041 8035 2099 8041
rect 2746 8044 15200 8072
rect 1394 7964 1400 8016
rect 1452 8004 1458 8016
rect 1489 8007 1547 8013
rect 1489 8004 1501 8007
rect 1452 7976 1501 8004
rect 1452 7964 1458 7976
rect 1489 7973 1501 7976
rect 1535 7973 1547 8007
rect 1489 7967 1547 7973
rect 1673 8007 1731 8013
rect 1673 7973 1685 8007
rect 1719 8004 1731 8007
rect 2746 8004 2774 8044
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 17957 8075 18015 8081
rect 17957 8041 17969 8075
rect 18003 8072 18015 8075
rect 18046 8072 18052 8084
rect 18003 8044 18052 8072
rect 18003 8041 18015 8044
rect 17957 8035 18015 8041
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 18325 8075 18383 8081
rect 18325 8041 18337 8075
rect 18371 8072 18383 8075
rect 18966 8072 18972 8084
rect 18371 8044 18972 8072
rect 18371 8041 18383 8044
rect 18325 8035 18383 8041
rect 18966 8032 18972 8044
rect 19024 8032 19030 8084
rect 19702 8072 19708 8084
rect 19663 8044 19708 8072
rect 19702 8032 19708 8044
rect 19760 8032 19766 8084
rect 20162 8072 20168 8084
rect 20123 8044 20168 8072
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20254 8032 20260 8084
rect 20312 8072 20318 8084
rect 20533 8075 20591 8081
rect 20533 8072 20545 8075
rect 20312 8044 20545 8072
rect 20312 8032 20318 8044
rect 20533 8041 20545 8044
rect 20579 8041 20591 8075
rect 20533 8035 20591 8041
rect 21361 8075 21419 8081
rect 21361 8041 21373 8075
rect 21407 8072 21419 8075
rect 21818 8072 21824 8084
rect 21407 8044 21824 8072
rect 21407 8041 21419 8044
rect 21361 8035 21419 8041
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 1719 7976 2774 8004
rect 1719 7973 1731 7976
rect 1673 7967 1731 7973
rect 3418 7964 3424 8016
rect 3476 8004 3482 8016
rect 4976 8007 5034 8013
rect 3476 7976 4752 8004
rect 3476 7964 3482 7976
rect 1762 7936 1768 7948
rect 1723 7908 1768 7936
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 3165 7939 3223 7945
rect 3165 7905 3177 7939
rect 3211 7936 3223 7939
rect 3510 7936 3516 7948
rect 3211 7908 3516 7936
rect 3211 7905 3223 7908
rect 3165 7899 3223 7905
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 3878 7896 3884 7948
rect 3936 7936 3942 7948
rect 4724 7945 4752 7976
rect 4976 7973 4988 8007
rect 5022 8004 5034 8007
rect 5534 8004 5540 8016
rect 5022 7976 5540 8004
rect 5022 7973 5034 7976
rect 4976 7967 5034 7973
rect 5534 7964 5540 7976
rect 5592 7964 5598 8016
rect 6086 7964 6092 8016
rect 6144 8004 6150 8016
rect 6426 8007 6484 8013
rect 6426 8004 6438 8007
rect 6144 7976 6438 8004
rect 6144 7964 6150 7976
rect 6426 7973 6438 7976
rect 6472 7973 6484 8007
rect 6426 7967 6484 7973
rect 8113 8007 8171 8013
rect 8113 7973 8125 8007
rect 8159 8004 8171 8007
rect 8202 8004 8208 8016
rect 8159 7976 8208 8004
rect 8159 7973 8171 7976
rect 8113 7967 8171 7973
rect 8202 7964 8208 7976
rect 8260 7964 8266 8016
rect 8573 8007 8631 8013
rect 8573 7973 8585 8007
rect 8619 8004 8631 8007
rect 8846 8004 8852 8016
rect 8619 7976 8852 8004
rect 8619 7973 8631 7976
rect 8573 7967 8631 7973
rect 4249 7939 4307 7945
rect 4249 7936 4261 7939
rect 3936 7908 4261 7936
rect 3936 7896 3942 7908
rect 4249 7905 4261 7908
rect 4295 7905 4307 7939
rect 4249 7899 4307 7905
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 8021 7939 8079 7945
rect 8021 7905 8033 7939
rect 8067 7936 8079 7939
rect 8588 7936 8616 7967
rect 8846 7964 8852 7976
rect 8904 7964 8910 8016
rect 20070 8004 20076 8016
rect 20031 7976 20076 8004
rect 20070 7964 20076 7976
rect 20128 7964 20134 8016
rect 20346 7964 20352 8016
rect 20404 8004 20410 8016
rect 20404 7976 21220 8004
rect 20404 7964 20410 7976
rect 21192 7948 21220 7976
rect 8067 7908 8616 7936
rect 20717 7939 20775 7945
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 20717 7905 20729 7939
rect 20763 7936 20775 7939
rect 20806 7936 20812 7948
rect 20763 7908 20812 7936
rect 20763 7905 20775 7908
rect 20717 7899 20775 7905
rect 20806 7896 20812 7908
rect 20864 7896 20870 7948
rect 21174 7936 21180 7948
rect 21135 7908 21180 7936
rect 21174 7896 21180 7908
rect 21232 7896 21238 7948
rect 21450 7936 21456 7948
rect 21411 7908 21456 7936
rect 21450 7896 21456 7908
rect 21508 7896 21514 7948
rect 3418 7868 3424 7880
rect 3379 7840 3424 7868
rect 3418 7828 3424 7840
rect 3476 7828 3482 7880
rect 4338 7868 4344 7880
rect 4299 7840 4344 7868
rect 4338 7828 4344 7840
rect 4396 7828 4402 7880
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 6178 7868 6184 7880
rect 4571 7840 4660 7868
rect 6139 7840 6184 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 1949 7735 2007 7741
rect 1949 7701 1961 7735
rect 1995 7732 2007 7735
rect 3050 7732 3056 7744
rect 1995 7704 3056 7732
rect 1995 7701 2007 7704
rect 1949 7695 2007 7701
rect 3050 7692 3056 7704
rect 3108 7692 3114 7744
rect 3142 7692 3148 7744
rect 3200 7732 3206 7744
rect 3881 7735 3939 7741
rect 3881 7732 3893 7735
rect 3200 7704 3893 7732
rect 3200 7692 3206 7704
rect 3881 7701 3893 7704
rect 3927 7701 3939 7735
rect 4632 7732 4660 7840
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 7432 7840 8217 7868
rect 7432 7828 7438 7840
rect 8205 7837 8217 7840
rect 8251 7837 8263 7871
rect 17678 7868 17684 7880
rect 17639 7840 17684 7868
rect 8205 7831 8263 7837
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7868 17923 7871
rect 17954 7868 17960 7880
rect 17911 7840 17960 7868
rect 17911 7837 17923 7840
rect 17865 7831 17923 7837
rect 17954 7828 17960 7840
rect 18012 7868 18018 7880
rect 18138 7868 18144 7880
rect 18012 7840 18144 7868
rect 18012 7828 18018 7840
rect 18138 7828 18144 7840
rect 18196 7828 18202 7880
rect 20349 7871 20407 7877
rect 20349 7837 20361 7871
rect 20395 7868 20407 7871
rect 20438 7868 20444 7880
rect 20395 7840 20444 7868
rect 20395 7837 20407 7840
rect 20349 7831 20407 7837
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 20901 7871 20959 7877
rect 20901 7837 20913 7871
rect 20947 7868 20959 7871
rect 21468 7868 21496 7896
rect 20947 7840 21496 7868
rect 20947 7837 20959 7840
rect 20901 7831 20959 7837
rect 6086 7800 6092 7812
rect 6047 7772 6092 7800
rect 6086 7760 6092 7772
rect 6144 7760 6150 7812
rect 7650 7800 7656 7812
rect 7611 7772 7656 7800
rect 7650 7760 7656 7772
rect 7708 7760 7714 7812
rect 12250 7760 12256 7812
rect 12308 7800 12314 7812
rect 20993 7803 21051 7809
rect 20993 7800 21005 7803
rect 12308 7772 21005 7800
rect 12308 7760 12314 7772
rect 20993 7769 21005 7772
rect 21039 7769 21051 7803
rect 20993 7763 21051 7769
rect 4982 7732 4988 7744
rect 4632 7704 4988 7732
rect 3881 7695 3939 7701
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 6822 7692 6828 7744
rect 6880 7732 6886 7744
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 6880 7704 7573 7732
rect 6880 7692 6886 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 21082 7732 21088 7744
rect 8904 7704 21088 7732
rect 8904 7692 8910 7704
rect 21082 7692 21088 7704
rect 21140 7692 21146 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 2133 7531 2191 7537
rect 2133 7528 2145 7531
rect 1820 7500 2145 7528
rect 1820 7488 1826 7500
rect 2133 7497 2145 7500
rect 2179 7497 2191 7531
rect 14734 7528 14740 7540
rect 2133 7491 2191 7497
rect 2746 7500 14740 7528
rect 1673 7463 1731 7469
rect 1673 7429 1685 7463
rect 1719 7460 1731 7463
rect 2746 7460 2774 7500
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 16850 7488 16856 7540
rect 16908 7528 16914 7540
rect 16945 7531 17003 7537
rect 16945 7528 16957 7531
rect 16908 7500 16957 7528
rect 16908 7488 16914 7500
rect 16945 7497 16957 7500
rect 16991 7497 17003 7531
rect 20806 7528 20812 7540
rect 20767 7500 20812 7528
rect 16945 7491 17003 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 2866 7460 2872 7472
rect 1719 7432 2774 7460
rect 2827 7432 2872 7460
rect 1719 7429 1731 7432
rect 1673 7423 1731 7429
rect 2866 7420 2872 7432
rect 2924 7420 2930 7472
rect 4890 7460 4896 7472
rect 4851 7432 4896 7460
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 4982 7420 4988 7472
rect 5040 7460 5046 7472
rect 7374 7460 7380 7472
rect 5040 7432 7380 7460
rect 5040 7420 5046 7432
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 1765 7395 1823 7401
rect 1765 7392 1777 7395
rect 1544 7364 1777 7392
rect 1544 7352 1550 7364
rect 1765 7361 1777 7364
rect 1811 7361 1823 7395
rect 3510 7392 3516 7404
rect 3423 7364 3516 7392
rect 1765 7355 1823 7361
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 3878 7392 3884 7404
rect 3839 7364 3884 7392
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 3528 7324 3556 7352
rect 5000 7324 5028 7420
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5534 7392 5540 7404
rect 5491 7364 5540 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7392 8815 7395
rect 9582 7392 9588 7404
rect 8803 7364 9588 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 9582 7352 9588 7364
rect 9640 7352 9646 7404
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7361 21419 7395
rect 21361 7355 21419 7361
rect 3528 7296 5028 7324
rect 5258 7284 5264 7336
rect 5316 7324 5322 7336
rect 5353 7327 5411 7333
rect 5353 7324 5365 7327
rect 5316 7296 5365 7324
rect 5316 7284 5322 7296
rect 5353 7293 5365 7296
rect 5399 7293 5411 7327
rect 5353 7287 5411 7293
rect 18325 7327 18383 7333
rect 18325 7293 18337 7327
rect 18371 7324 18383 7327
rect 19334 7324 19340 7336
rect 18371 7296 19340 7324
rect 18371 7293 18383 7296
rect 18325 7287 18383 7293
rect 19334 7284 19340 7296
rect 19392 7284 19398 7336
rect 20990 7324 20996 7336
rect 19536 7296 20996 7324
rect 1394 7216 1400 7268
rect 1452 7256 1458 7268
rect 1489 7259 1547 7265
rect 1489 7256 1501 7259
rect 1452 7228 1501 7256
rect 1452 7216 1458 7228
rect 1489 7225 1501 7228
rect 1535 7256 1547 7259
rect 1949 7259 2007 7265
rect 1949 7256 1961 7259
rect 1535 7228 1961 7256
rect 1535 7225 1547 7228
rect 1489 7219 1547 7225
rect 1949 7225 1961 7228
rect 1995 7225 2007 7259
rect 1949 7219 2007 7225
rect 3237 7259 3295 7265
rect 3237 7225 3249 7259
rect 3283 7256 3295 7259
rect 4154 7256 4160 7268
rect 3283 7228 4160 7256
rect 3283 7225 3295 7228
rect 3237 7219 3295 7225
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 4798 7216 4804 7268
rect 4856 7256 4862 7268
rect 5276 7256 5304 7284
rect 8570 7265 8576 7268
rect 4856 7228 5304 7256
rect 8512 7259 8576 7265
rect 4856 7216 4862 7228
rect 8512 7225 8524 7259
rect 8558 7225 8576 7259
rect 8512 7219 8576 7225
rect 8570 7216 8576 7219
rect 8628 7216 8634 7268
rect 18080 7259 18138 7265
rect 18080 7225 18092 7259
rect 18126 7256 18138 7259
rect 19536 7256 19564 7296
rect 20990 7284 20996 7296
rect 21048 7324 21054 7336
rect 21376 7324 21404 7355
rect 21048 7296 21404 7324
rect 21048 7284 21054 7296
rect 18126 7228 19564 7256
rect 19604 7259 19662 7265
rect 18126 7225 18138 7228
rect 18080 7219 18138 7225
rect 19604 7225 19616 7259
rect 19650 7256 19662 7259
rect 19794 7256 19800 7268
rect 19650 7228 19800 7256
rect 19650 7225 19662 7228
rect 19604 7219 19662 7225
rect 19794 7216 19800 7228
rect 19852 7216 19858 7268
rect 3329 7191 3387 7197
rect 3329 7157 3341 7191
rect 3375 7188 3387 7191
rect 4246 7188 4252 7200
rect 3375 7160 4252 7188
rect 3375 7157 3387 7160
rect 3329 7151 3387 7157
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 5040 7160 5273 7188
rect 5040 7148 5046 7160
rect 5261 7157 5273 7160
rect 5307 7188 5319 7191
rect 5442 7188 5448 7200
rect 5307 7160 5448 7188
rect 5307 7157 5319 7160
rect 5261 7151 5319 7157
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5718 7188 5724 7200
rect 5679 7160 5724 7188
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 20714 7188 20720 7200
rect 20675 7160 20720 7188
rect 20714 7148 20720 7160
rect 20772 7148 20778 7200
rect 21174 7188 21180 7200
rect 21135 7160 21180 7188
rect 21174 7148 21180 7160
rect 21232 7148 21238 7200
rect 21266 7148 21272 7200
rect 21324 7188 21330 7200
rect 21324 7160 21369 7188
rect 21324 7148 21330 7160
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 1670 6984 1676 6996
rect 1452 6956 1676 6984
rect 1452 6944 1458 6956
rect 1670 6944 1676 6956
rect 1728 6944 1734 6996
rect 5261 6987 5319 6993
rect 5261 6953 5273 6987
rect 5307 6984 5319 6987
rect 5718 6984 5724 6996
rect 5307 6956 5724 6984
rect 5307 6953 5319 6956
rect 5261 6947 5319 6953
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 20990 6984 20996 6996
rect 20951 6956 20996 6984
rect 20990 6944 20996 6956
rect 21048 6944 21054 6996
rect 1486 6848 1492 6860
rect 1447 6820 1492 6848
rect 1486 6808 1492 6820
rect 1544 6808 1550 6860
rect 2958 6848 2964 6860
rect 3016 6857 3022 6860
rect 2928 6820 2964 6848
rect 2958 6808 2964 6820
rect 3016 6811 3028 6857
rect 3237 6851 3295 6857
rect 3237 6817 3249 6851
rect 3283 6848 3295 6851
rect 3418 6848 3424 6860
rect 3283 6820 3424 6848
rect 3283 6817 3295 6820
rect 3237 6811 3295 6817
rect 3016 6808 3022 6811
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 19610 6848 19616 6860
rect 19392 6820 19616 6848
rect 19392 6808 19398 6820
rect 19610 6808 19616 6820
rect 19668 6808 19674 6860
rect 19880 6851 19938 6857
rect 19880 6817 19892 6851
rect 19926 6848 19938 6851
rect 20714 6848 20720 6860
rect 19926 6820 20720 6848
rect 19926 6817 19938 6820
rect 19880 6811 19938 6817
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 21177 6851 21235 6857
rect 21177 6817 21189 6851
rect 21223 6848 21235 6851
rect 21450 6848 21456 6860
rect 21223 6820 21456 6848
rect 21223 6817 21235 6820
rect 21177 6811 21235 6817
rect 21450 6808 21456 6820
rect 21508 6808 21514 6860
rect 5350 6780 5356 6792
rect 5311 6752 5356 6780
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 5445 6783 5503 6789
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 5534 6780 5540 6792
rect 5491 6752 5540 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 4893 6715 4951 6721
rect 4893 6681 4905 6715
rect 4939 6712 4951 6715
rect 5074 6712 5080 6724
rect 4939 6684 5080 6712
rect 4939 6681 4951 6684
rect 4893 6675 4951 6681
rect 5074 6672 5080 6684
rect 5132 6672 5138 6724
rect 21269 6715 21327 6721
rect 21269 6712 21281 6715
rect 20548 6684 21281 6712
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 1857 6647 1915 6653
rect 1857 6613 1869 6647
rect 1903 6644 1915 6647
rect 3694 6644 3700 6656
rect 1903 6616 3700 6644
rect 1903 6613 1915 6616
rect 1857 6607 1915 6613
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 20548 6644 20576 6684
rect 21269 6681 21281 6684
rect 21315 6681 21327 6715
rect 21269 6675 21327 6681
rect 11848 6616 20576 6644
rect 11848 6604 11854 6616
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 1578 6400 1584 6452
rect 1636 6440 1642 6452
rect 10502 6440 10508 6452
rect 1636 6412 10508 6440
rect 1636 6400 1642 6412
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 21082 6332 21088 6384
rect 21140 6372 21146 6384
rect 21269 6375 21327 6381
rect 21269 6372 21281 6375
rect 21140 6344 21281 6372
rect 21140 6332 21146 6344
rect 21269 6341 21281 6344
rect 21315 6341 21327 6375
rect 21269 6335 21327 6341
rect 20717 6307 20775 6313
rect 20717 6273 20729 6307
rect 20763 6304 20775 6307
rect 21174 6304 21180 6316
rect 20763 6276 21180 6304
rect 20763 6273 20775 6276
rect 20717 6267 20775 6273
rect 21174 6264 21180 6276
rect 21232 6264 21238 6316
rect 1486 6168 1492 6180
rect 1447 6140 1492 6168
rect 1486 6128 1492 6140
rect 1544 6128 1550 6180
rect 1673 6171 1731 6177
rect 1673 6137 1685 6171
rect 1719 6168 1731 6171
rect 14642 6168 14648 6180
rect 1719 6140 14648 6168
rect 1719 6137 1731 6140
rect 1673 6131 1731 6137
rect 14642 6128 14648 6140
rect 14700 6128 14706 6180
rect 21177 6171 21235 6177
rect 21177 6137 21189 6171
rect 21223 6168 21235 6171
rect 21450 6168 21456 6180
rect 21223 6140 21456 6168
rect 21223 6137 21235 6140
rect 21177 6131 21235 6137
rect 21450 6128 21456 6140
rect 21508 6128 21514 6180
rect 1504 6100 1532 6128
rect 1765 6103 1823 6109
rect 1765 6100 1777 6103
rect 1504 6072 1777 6100
rect 1765 6069 1777 6072
rect 1811 6069 1823 6103
rect 1765 6063 1823 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 1581 5899 1639 5905
rect 1581 5896 1593 5899
rect 1452 5868 1593 5896
rect 1452 5856 1458 5868
rect 1581 5865 1593 5868
rect 1627 5865 1639 5899
rect 1581 5859 1639 5865
rect 21085 5899 21143 5905
rect 21085 5865 21097 5899
rect 21131 5896 21143 5899
rect 21266 5896 21272 5908
rect 21131 5868 21272 5896
rect 21131 5865 21143 5868
rect 21085 5859 21143 5865
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 21361 5899 21419 5905
rect 21361 5865 21373 5899
rect 21407 5865 21419 5899
rect 21361 5859 21419 5865
rect 9214 5788 9220 5840
rect 9272 5828 9278 5840
rect 21376 5828 21404 5859
rect 9272 5800 21404 5828
rect 9272 5788 9278 5800
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5760 1458 5772
rect 1673 5763 1731 5769
rect 1673 5760 1685 5763
rect 1452 5732 1685 5760
rect 1452 5720 1458 5732
rect 1673 5729 1685 5732
rect 1719 5729 1731 5763
rect 1673 5723 1731 5729
rect 20162 5720 20168 5772
rect 20220 5760 20226 5772
rect 20717 5763 20775 5769
rect 20717 5760 20729 5763
rect 20220 5732 20729 5760
rect 20220 5720 20226 5732
rect 20717 5729 20729 5732
rect 20763 5729 20775 5763
rect 20717 5723 20775 5729
rect 21269 5763 21327 5769
rect 21269 5729 21281 5763
rect 21315 5760 21327 5763
rect 21542 5760 21548 5772
rect 21315 5732 21548 5760
rect 21315 5729 21327 5732
rect 21269 5723 21327 5729
rect 21542 5720 21548 5732
rect 21600 5720 21606 5772
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 20625 5695 20683 5701
rect 20625 5661 20637 5695
rect 20671 5692 20683 5695
rect 21358 5692 21364 5704
rect 20671 5664 21364 5692
rect 20671 5661 20683 5664
rect 20625 5655 20683 5661
rect 20548 5624 20576 5655
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 20714 5624 20720 5636
rect 20548 5596 20720 5624
rect 20714 5584 20720 5596
rect 20772 5584 20778 5636
rect 20162 5556 20168 5568
rect 20123 5528 20168 5556
rect 20162 5516 20168 5528
rect 20220 5516 20226 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5284 1731 5287
rect 6270 5284 6276 5296
rect 1719 5256 6276 5284
rect 1719 5253 1731 5256
rect 1673 5247 1731 5253
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 20898 5244 20904 5296
rect 20956 5284 20962 5296
rect 21269 5287 21327 5293
rect 21269 5284 21281 5287
rect 20956 5256 21281 5284
rect 20956 5244 20962 5256
rect 21269 5253 21281 5256
rect 21315 5253 21327 5287
rect 21269 5247 21327 5253
rect 1486 5148 1492 5160
rect 1447 5120 1492 5148
rect 1486 5108 1492 5120
rect 1544 5148 1550 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1544 5120 1777 5148
rect 1544 5108 1550 5120
rect 1765 5117 1777 5120
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 21177 5151 21235 5157
rect 21177 5117 21189 5151
rect 21223 5148 21235 5151
rect 21450 5148 21456 5160
rect 21223 5120 21456 5148
rect 21223 5117 21235 5120
rect 21177 5111 21235 5117
rect 21450 5108 21456 5120
rect 21508 5108 21514 5160
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 3326 4808 3332 4820
rect 1627 4780 3332 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 21358 4808 21364 4820
rect 21319 4780 21364 4808
rect 21358 4768 21364 4780
rect 21416 4768 21422 4820
rect 1949 4743 2007 4749
rect 1949 4740 1961 4743
rect 1412 4712 1961 4740
rect 1412 4684 1440 4712
rect 1949 4709 1961 4712
rect 1995 4709 2007 4743
rect 1949 4703 2007 4709
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 1670 4672 1676 4684
rect 1631 4644 1676 4672
rect 1670 4632 1676 4644
rect 1728 4672 1734 4684
rect 2133 4675 2191 4681
rect 2133 4672 2145 4675
rect 1728 4644 2145 4672
rect 1728 4632 1734 4644
rect 2133 4641 2145 4644
rect 2179 4641 2191 4675
rect 2133 4635 2191 4641
rect 20809 4675 20867 4681
rect 20809 4641 20821 4675
rect 20855 4672 20867 4675
rect 21266 4672 21272 4684
rect 20855 4644 21272 4672
rect 20855 4641 20867 4644
rect 20809 4635 20867 4641
rect 21266 4632 21272 4644
rect 21324 4632 21330 4684
rect 21542 4672 21548 4684
rect 21503 4644 21548 4672
rect 21542 4632 21548 4644
rect 21600 4632 21606 4684
rect 20162 4604 20168 4616
rect 1872 4576 20168 4604
rect 1872 4545 1900 4576
rect 20162 4564 20168 4576
rect 20220 4564 20226 4616
rect 20993 4607 21051 4613
rect 20993 4573 21005 4607
rect 21039 4604 21051 4607
rect 21560 4604 21588 4632
rect 21039 4576 21588 4604
rect 21039 4573 21051 4576
rect 20993 4567 21051 4573
rect 1857 4539 1915 4545
rect 1857 4505 1869 4539
rect 1903 4505 1915 4539
rect 1857 4499 1915 4505
rect 6362 4496 6368 4548
rect 6420 4536 6426 4548
rect 21085 4539 21143 4545
rect 21085 4536 21097 4539
rect 6420 4508 21097 4536
rect 6420 4496 6426 4508
rect 21085 4505 21097 4508
rect 21131 4505 21143 4539
rect 21085 4499 21143 4505
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 1581 4267 1639 4273
rect 1581 4233 1593 4267
rect 1627 4264 1639 4267
rect 5350 4264 5356 4276
rect 1627 4236 5356 4264
rect 1627 4233 1639 4236
rect 1581 4227 1639 4233
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 1394 4060 1400 4072
rect 1355 4032 1400 4060
rect 1394 4020 1400 4032
rect 1452 4060 1458 4072
rect 1673 4063 1731 4069
rect 1673 4060 1685 4063
rect 1452 4032 1685 4060
rect 1452 4020 1458 4032
rect 1673 4029 1685 4032
rect 1719 4029 1731 4063
rect 1673 4023 1731 4029
rect 21269 4063 21327 4069
rect 21269 4029 21281 4063
rect 21315 4060 21327 4063
rect 21542 4060 21548 4072
rect 21315 4032 21548 4060
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 21542 4020 21548 4032
rect 21600 4020 21606 4072
rect 19886 3884 19892 3936
rect 19944 3924 19950 3936
rect 21361 3927 21419 3933
rect 21361 3924 21373 3927
rect 19944 3896 21373 3924
rect 19944 3884 19950 3896
rect 21361 3893 21373 3896
rect 21407 3893 21419 3927
rect 21361 3887 21419 3893
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 4338 3720 4344 3732
rect 1627 3692 4344 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 4338 3680 4344 3692
rect 4396 3680 4402 3732
rect 21361 3723 21419 3729
rect 21361 3689 21373 3723
rect 21407 3720 21419 3723
rect 21634 3720 21640 3732
rect 21407 3692 21640 3720
rect 21407 3689 21419 3692
rect 21361 3683 21419 3689
rect 21634 3680 21640 3692
rect 21692 3680 21698 3732
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3584 1458 3596
rect 1857 3587 1915 3593
rect 1857 3584 1869 3587
rect 1452 3556 1869 3584
rect 1452 3544 1458 3556
rect 1857 3553 1869 3556
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 21085 3587 21143 3593
rect 21085 3553 21097 3587
rect 21131 3584 21143 3587
rect 21542 3584 21548 3596
rect 21131 3556 21548 3584
rect 21131 3553 21143 3556
rect 21085 3547 21143 3553
rect 21542 3544 21548 3556
rect 21600 3544 21606 3596
rect 20901 3519 20959 3525
rect 20901 3485 20913 3519
rect 20947 3516 20959 3519
rect 21450 3516 21456 3528
rect 20947 3488 21456 3516
rect 20947 3485 20959 3488
rect 20901 3479 20959 3485
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 1486 3408 1492 3460
rect 1544 3448 1550 3460
rect 1673 3451 1731 3457
rect 1673 3448 1685 3451
rect 1544 3420 1685 3448
rect 1544 3408 1550 3420
rect 1673 3417 1685 3420
rect 1719 3417 1731 3451
rect 1673 3411 1731 3417
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 2225 3451 2283 3457
rect 2225 3448 2237 3451
rect 2004 3420 2237 3448
rect 2004 3408 2010 3420
rect 2225 3417 2237 3420
rect 2271 3417 2283 3451
rect 2225 3411 2283 3417
rect 19978 3408 19984 3460
rect 20036 3448 20042 3460
rect 20990 3448 20996 3460
rect 20036 3420 20996 3448
rect 20036 3408 20042 3420
rect 20990 3408 20996 3420
rect 21048 3408 21054 3460
rect 21269 3451 21327 3457
rect 21269 3417 21281 3451
rect 21315 3448 21327 3451
rect 21315 3420 21588 3448
rect 21315 3417 21327 3420
rect 21269 3411 21327 3417
rect 21560 3392 21588 3420
rect 1762 3340 1768 3392
rect 1820 3380 1826 3392
rect 2041 3383 2099 3389
rect 2041 3380 2053 3383
rect 1820 3352 2053 3380
rect 1820 3340 1826 3352
rect 2041 3349 2053 3352
rect 2087 3349 2099 3383
rect 20622 3380 20628 3392
rect 20583 3352 20628 3380
rect 2041 3343 2099 3349
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 21542 3340 21548 3392
rect 21600 3340 21606 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 2133 3179 2191 3185
rect 2133 3145 2145 3179
rect 2179 3176 2191 3179
rect 4246 3176 4252 3188
rect 2179 3148 4252 3176
rect 2179 3145 2191 3148
rect 2133 3139 2191 3145
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4801 3179 4859 3185
rect 4801 3145 4813 3179
rect 4847 3176 4859 3179
rect 5166 3176 5172 3188
rect 4847 3148 5172 3176
rect 4847 3145 4859 3148
rect 4801 3139 4859 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5629 3179 5687 3185
rect 5629 3145 5641 3179
rect 5675 3176 5687 3179
rect 6730 3176 6736 3188
rect 5675 3148 6736 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 20438 3136 20444 3188
rect 20496 3176 20502 3188
rect 20809 3179 20867 3185
rect 20809 3176 20821 3179
rect 20496 3148 20821 3176
rect 20496 3136 20502 3148
rect 20809 3145 20821 3148
rect 20855 3145 20867 3179
rect 20809 3139 20867 3145
rect 20990 3136 20996 3188
rect 21048 3176 21054 3188
rect 21361 3179 21419 3185
rect 21361 3176 21373 3179
rect 21048 3148 21373 3176
rect 21048 3136 21054 3148
rect 21361 3145 21373 3148
rect 21407 3145 21419 3179
rect 21361 3139 21419 3145
rect 1581 3111 1639 3117
rect 1581 3077 1593 3111
rect 1627 3108 1639 3111
rect 4982 3108 4988 3120
rect 1627 3080 4988 3108
rect 1627 3077 1639 3080
rect 1581 3071 1639 3077
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 20533 3111 20591 3117
rect 20533 3077 20545 3111
rect 20579 3108 20591 3111
rect 20579 3080 21312 3108
rect 20579 3077 20591 3080
rect 20533 3071 20591 3077
rect 5902 3040 5908 3052
rect 2746 3012 5908 3040
rect 1394 2972 1400 2984
rect 1355 2944 1400 2972
rect 1394 2932 1400 2944
rect 1452 2932 1458 2984
rect 1670 2972 1676 2984
rect 1631 2944 1676 2972
rect 1670 2932 1676 2944
rect 1728 2932 1734 2984
rect 1946 2972 1952 2984
rect 1907 2944 1952 2972
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 2746 2972 2774 3012
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 20622 3040 20628 3052
rect 20548 3012 20628 3040
rect 20548 2984 20576 3012
rect 20622 3000 20628 3012
rect 20680 3040 20686 3052
rect 20680 3012 21036 3040
rect 20680 3000 20686 3012
rect 4982 2972 4988 2984
rect 2424 2944 2774 2972
rect 4943 2944 4988 2972
rect 1412 2904 1440 2932
rect 2225 2907 2283 2913
rect 2225 2904 2237 2907
rect 1412 2876 2237 2904
rect 2225 2873 2237 2876
rect 2271 2873 2283 2907
rect 2225 2867 2283 2873
rect 1857 2839 1915 2845
rect 1857 2805 1869 2839
rect 1903 2836 1915 2839
rect 2424 2836 2452 2944
rect 4982 2932 4988 2944
rect 5040 2932 5046 2984
rect 5813 2975 5871 2981
rect 5813 2941 5825 2975
rect 5859 2972 5871 2975
rect 11514 2972 11520 2984
rect 5859 2944 11520 2972
rect 5859 2941 5871 2944
rect 5813 2935 5871 2941
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 20530 2932 20536 2984
rect 20588 2932 20594 2984
rect 20717 2975 20775 2981
rect 20717 2941 20729 2975
rect 20763 2972 20775 2975
rect 20806 2972 20812 2984
rect 20763 2944 20812 2972
rect 20763 2941 20775 2944
rect 20717 2935 20775 2941
rect 20806 2932 20812 2944
rect 20864 2932 20870 2984
rect 21008 2981 21036 3012
rect 21284 2984 21312 3080
rect 20993 2975 21051 2981
rect 20993 2941 21005 2975
rect 21039 2941 21051 2975
rect 21266 2972 21272 2984
rect 21179 2944 21272 2972
rect 20993 2935 21051 2941
rect 21266 2932 21272 2944
rect 21324 2932 21330 2984
rect 21542 2972 21548 2984
rect 21503 2944 21548 2972
rect 21542 2932 21548 2944
rect 21600 2932 21606 2984
rect 2501 2907 2559 2913
rect 2501 2873 2513 2907
rect 2547 2904 2559 2907
rect 2866 2904 2872 2916
rect 2547 2876 2872 2904
rect 2547 2873 2559 2876
rect 2501 2867 2559 2873
rect 2866 2864 2872 2876
rect 2924 2864 2930 2916
rect 5442 2864 5448 2916
rect 5500 2904 5506 2916
rect 15381 2907 15439 2913
rect 15381 2904 15393 2907
rect 5500 2876 15393 2904
rect 5500 2864 5506 2876
rect 15381 2873 15393 2876
rect 15427 2873 15439 2907
rect 15562 2904 15568 2916
rect 15523 2876 15568 2904
rect 15381 2867 15439 2873
rect 15562 2864 15568 2876
rect 15620 2864 15626 2916
rect 20349 2907 20407 2913
rect 20349 2873 20361 2907
rect 20395 2904 20407 2907
rect 20622 2904 20628 2916
rect 20395 2876 20628 2904
rect 20395 2873 20407 2876
rect 20349 2867 20407 2873
rect 20622 2864 20628 2876
rect 20680 2864 20686 2916
rect 1903 2808 2452 2836
rect 2685 2839 2743 2845
rect 1903 2805 1915 2808
rect 1857 2799 1915 2805
rect 2685 2805 2697 2839
rect 2731 2836 2743 2839
rect 2774 2836 2780 2848
rect 2731 2808 2780 2836
rect 2731 2805 2743 2808
rect 2685 2799 2743 2805
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 18138 2796 18144 2848
rect 18196 2836 18202 2848
rect 21085 2839 21143 2845
rect 21085 2836 21097 2839
rect 18196 2808 21097 2836
rect 18196 2796 18202 2808
rect 21085 2805 21097 2808
rect 21131 2805 21143 2839
rect 21085 2799 21143 2805
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 2038 2632 2044 2644
rect 1903 2604 2044 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 2682 2632 2688 2644
rect 2179 2604 2688 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 2958 2632 2964 2644
rect 2919 2604 2964 2632
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 5166 2632 5172 2644
rect 3375 2604 5172 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 11514 2632 11520 2644
rect 11475 2604 11520 2632
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 15562 2592 15568 2644
rect 15620 2632 15626 2644
rect 16117 2635 16175 2641
rect 16117 2632 16129 2635
rect 15620 2604 16129 2632
rect 15620 2592 15626 2604
rect 16117 2601 16129 2604
rect 16163 2601 16175 2635
rect 16117 2595 16175 2601
rect 19426 2592 19432 2644
rect 19484 2632 19490 2644
rect 20165 2635 20223 2641
rect 20165 2632 20177 2635
rect 19484 2604 20177 2632
rect 19484 2592 19490 2604
rect 20165 2601 20177 2604
rect 20211 2601 20223 2635
rect 20165 2595 20223 2601
rect 20441 2635 20499 2641
rect 20441 2601 20453 2635
rect 20487 2601 20499 2635
rect 20441 2595 20499 2601
rect 20993 2635 21051 2641
rect 20993 2601 21005 2635
rect 21039 2632 21051 2635
rect 21910 2632 21916 2644
rect 21039 2604 21916 2632
rect 21039 2601 21051 2604
rect 20993 2595 21051 2601
rect 2774 2564 2780 2576
rect 1964 2536 2780 2564
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 1964 2505 1992 2536
rect 2774 2524 2780 2536
rect 2832 2524 2838 2576
rect 7098 2564 7104 2576
rect 7059 2536 7104 2564
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 17954 2524 17960 2576
rect 18012 2564 18018 2576
rect 20456 2564 20484 2595
rect 21910 2592 21916 2604
rect 21968 2592 21974 2644
rect 18012 2536 20484 2564
rect 18012 2524 18018 2536
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2465 1731 2499
rect 1673 2459 1731 2465
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2465 2007 2499
rect 2317 2499 2375 2505
rect 2317 2496 2329 2499
rect 1949 2459 2007 2465
rect 2240 2468 2329 2496
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 1688 2292 1716 2459
rect 2240 2360 2268 2468
rect 2317 2465 2329 2468
rect 2363 2465 2375 2499
rect 2317 2459 2375 2465
rect 2406 2456 2412 2508
rect 2464 2496 2470 2508
rect 3237 2499 3295 2505
rect 3237 2496 3249 2499
rect 2464 2468 3249 2496
rect 2464 2456 2470 2468
rect 3237 2465 3249 2468
rect 3283 2465 3295 2499
rect 3510 2496 3516 2508
rect 3471 2468 3516 2496
rect 3237 2459 3295 2465
rect 3252 2428 3280 2459
rect 3510 2456 3516 2468
rect 3568 2496 3574 2508
rect 3881 2499 3939 2505
rect 3881 2496 3893 2499
rect 3568 2468 3893 2496
rect 3568 2456 3574 2468
rect 3881 2465 3893 2468
rect 3927 2465 3939 2499
rect 11698 2496 11704 2508
rect 11659 2468 11704 2496
rect 3881 2459 3939 2465
rect 11698 2456 11704 2468
rect 11756 2496 11762 2508
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11756 2468 11897 2496
rect 11756 2456 11762 2468
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 16114 2456 16120 2508
rect 16172 2496 16178 2508
rect 16301 2499 16359 2505
rect 16301 2496 16313 2499
rect 16172 2468 16313 2496
rect 16172 2456 16178 2468
rect 16301 2465 16313 2468
rect 16347 2465 16359 2499
rect 16301 2459 16359 2465
rect 19705 2499 19763 2505
rect 19705 2465 19717 2499
rect 19751 2496 19763 2499
rect 20346 2496 20352 2508
rect 19751 2468 20352 2496
rect 19751 2465 19763 2468
rect 19705 2459 19763 2465
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 20622 2496 20628 2508
rect 20583 2468 20628 2496
rect 20622 2456 20628 2468
rect 20680 2456 20686 2508
rect 20714 2456 20720 2508
rect 20772 2496 20778 2508
rect 20901 2499 20959 2505
rect 20901 2496 20913 2499
rect 20772 2468 20913 2496
rect 20772 2456 20778 2468
rect 20901 2465 20913 2468
rect 20947 2465 20959 2499
rect 21174 2496 21180 2508
rect 21135 2468 21180 2496
rect 20901 2459 20959 2465
rect 21174 2456 21180 2468
rect 21232 2456 21238 2508
rect 21450 2496 21456 2508
rect 21411 2468 21456 2496
rect 21450 2456 21456 2468
rect 21508 2456 21514 2508
rect 3605 2431 3663 2437
rect 3605 2428 3617 2431
rect 3252 2400 3617 2428
rect 3605 2397 3617 2400
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 20073 2431 20131 2437
rect 5040 2400 16574 2428
rect 5040 2388 5046 2400
rect 3053 2363 3111 2369
rect 3053 2360 3065 2363
rect 2240 2332 3065 2360
rect 3053 2329 3065 2332
rect 3099 2329 3111 2363
rect 3053 2323 3111 2329
rect 6914 2320 6920 2372
rect 6972 2360 6978 2372
rect 16546 2360 16574 2400
rect 20073 2397 20085 2431
rect 20119 2428 20131 2431
rect 21192 2428 21220 2456
rect 20119 2400 21220 2428
rect 20119 2397 20131 2400
rect 20073 2391 20131 2397
rect 20717 2363 20775 2369
rect 20717 2360 20729 2363
rect 6972 2332 7017 2360
rect 16546 2332 20729 2360
rect 6972 2320 6978 2332
rect 20717 2329 20729 2332
rect 20763 2329 20775 2363
rect 20717 2323 20775 2329
rect 2866 2292 2872 2304
rect 1688 2264 2872 2292
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16393 2295 16451 2301
rect 16393 2292 16405 2295
rect 16172 2264 16405 2292
rect 16172 2252 16178 2264
rect 16393 2261 16405 2264
rect 16439 2261 16451 2295
rect 16393 2255 16451 2261
rect 20438 2252 20444 2304
rect 20496 2292 20502 2304
rect 21361 2295 21419 2301
rect 21361 2292 21373 2295
rect 20496 2264 21373 2292
rect 20496 2252 20502 2264
rect 21361 2261 21373 2264
rect 21407 2261 21419 2295
rect 21361 2255 21419 2261
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 1578 2048 1584 2100
rect 1636 2088 1642 2100
rect 4154 2088 4160 2100
rect 1636 2060 4160 2088
rect 1636 2048 1642 2060
rect 4154 2048 4160 2060
rect 4212 2048 4218 2100
<< via1 >>
rect 2688 20884 2740 20936
rect 3516 20884 3568 20936
rect 1860 20816 1912 20868
rect 3424 20816 3476 20868
rect 1400 20748 1452 20800
rect 2872 20748 2924 20800
rect 17960 20748 18012 20800
rect 21456 20748 21508 20800
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 2780 20544 2832 20596
rect 2964 20587 3016 20596
rect 2964 20553 2973 20587
rect 2973 20553 3007 20587
rect 3007 20553 3016 20587
rect 2964 20544 3016 20553
rect 3332 20587 3384 20596
rect 3332 20553 3341 20587
rect 3341 20553 3375 20587
rect 3375 20553 3384 20587
rect 3332 20544 3384 20553
rect 3792 20544 3844 20596
rect 9404 20544 9456 20596
rect 9956 20544 10008 20596
rect 1492 20476 1544 20528
rect 3884 20519 3936 20528
rect 3884 20485 3893 20519
rect 3893 20485 3927 20519
rect 3927 20485 3936 20519
rect 3884 20476 3936 20485
rect 4344 20476 4396 20528
rect 4804 20519 4856 20528
rect 4804 20485 4813 20519
rect 4813 20485 4847 20519
rect 4847 20485 4856 20519
rect 4804 20476 4856 20485
rect 5264 20519 5316 20528
rect 5264 20485 5273 20519
rect 5273 20485 5307 20519
rect 5307 20485 5316 20519
rect 5264 20476 5316 20485
rect 6736 20476 6788 20528
rect 7472 20476 7524 20528
rect 1032 20340 1084 20392
rect 2596 20408 2648 20460
rect 2780 20408 2832 20460
rect 10048 20476 10100 20528
rect 9864 20408 9916 20460
rect 572 20272 624 20324
rect 1492 20315 1544 20324
rect 1492 20281 1501 20315
rect 1501 20281 1535 20315
rect 1535 20281 1544 20315
rect 1492 20272 1544 20281
rect 2136 20315 2188 20324
rect 2136 20281 2145 20315
rect 2145 20281 2179 20315
rect 2179 20281 2188 20315
rect 2136 20272 2188 20281
rect 2504 20272 2556 20324
rect 2228 20204 2280 20256
rect 3884 20340 3936 20392
rect 5080 20340 5132 20392
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 6092 20383 6144 20392
rect 6092 20349 6101 20383
rect 6101 20349 6135 20383
rect 6135 20349 6144 20383
rect 6092 20340 6144 20349
rect 6552 20383 6604 20392
rect 6552 20349 6561 20383
rect 6561 20349 6595 20383
rect 6595 20349 6604 20383
rect 6552 20340 6604 20349
rect 7012 20340 7064 20392
rect 7380 20383 7432 20392
rect 7380 20349 7389 20383
rect 7389 20349 7423 20383
rect 7423 20349 7432 20383
rect 7380 20340 7432 20349
rect 7840 20383 7892 20392
rect 7840 20349 7849 20383
rect 7849 20349 7883 20383
rect 7883 20349 7892 20383
rect 7840 20340 7892 20349
rect 8208 20383 8260 20392
rect 8208 20349 8217 20383
rect 8217 20349 8251 20383
rect 8251 20349 8260 20383
rect 8208 20340 8260 20349
rect 8668 20383 8720 20392
rect 8668 20349 8677 20383
rect 8677 20349 8711 20383
rect 8711 20349 8720 20383
rect 8668 20340 8720 20349
rect 9128 20340 9180 20392
rect 9496 20383 9548 20392
rect 9496 20349 9505 20383
rect 9505 20349 9539 20383
rect 9539 20349 9548 20383
rect 9496 20340 9548 20349
rect 11980 20544 12032 20596
rect 13360 20544 13412 20596
rect 15936 20544 15988 20596
rect 17960 20544 18012 20596
rect 18880 20544 18932 20596
rect 12164 20476 12216 20528
rect 12256 20476 12308 20528
rect 12808 20476 12860 20528
rect 13728 20476 13780 20528
rect 14188 20476 14240 20528
rect 14648 20476 14700 20528
rect 15200 20476 15252 20528
rect 15476 20476 15528 20528
rect 20168 20544 20220 20596
rect 20536 20544 20588 20596
rect 19708 20519 19760 20528
rect 19708 20485 19717 20519
rect 19717 20485 19751 20519
rect 19751 20485 19760 20519
rect 19708 20476 19760 20485
rect 20444 20519 20496 20528
rect 20444 20485 20453 20519
rect 20453 20485 20487 20519
rect 20487 20485 20496 20519
rect 20444 20476 20496 20485
rect 22744 20476 22796 20528
rect 10416 20340 10468 20392
rect 10784 20340 10836 20392
rect 11244 20340 11296 20392
rect 16304 20408 16356 20460
rect 19340 20408 19392 20460
rect 3056 20315 3108 20324
rect 3056 20281 3065 20315
rect 3065 20281 3099 20315
rect 3099 20281 3108 20315
rect 3056 20272 3108 20281
rect 3332 20272 3384 20324
rect 3700 20272 3752 20324
rect 4068 20315 4120 20324
rect 4068 20281 4077 20315
rect 4077 20281 4111 20315
rect 4111 20281 4120 20315
rect 4068 20272 4120 20281
rect 4896 20272 4948 20324
rect 3608 20204 3660 20256
rect 4252 20204 4304 20256
rect 6276 20247 6328 20256
rect 6276 20213 6285 20247
rect 6285 20213 6319 20247
rect 6319 20213 6328 20247
rect 6276 20204 6328 20213
rect 11796 20340 11848 20392
rect 12072 20340 12124 20392
rect 12532 20340 12584 20392
rect 12716 20383 12768 20392
rect 12716 20349 12725 20383
rect 12725 20349 12759 20383
rect 12759 20349 12768 20383
rect 12716 20340 12768 20349
rect 12900 20340 12952 20392
rect 16764 20340 16816 20392
rect 18420 20383 18472 20392
rect 11980 20272 12032 20324
rect 6644 20204 6696 20256
rect 6920 20204 6972 20256
rect 7196 20204 7248 20256
rect 8760 20204 8812 20256
rect 9036 20204 9088 20256
rect 9680 20247 9732 20256
rect 9680 20213 9689 20247
rect 9689 20213 9723 20247
rect 9723 20213 9732 20247
rect 9680 20204 9732 20213
rect 9956 20247 10008 20256
rect 9956 20213 9965 20247
rect 9965 20213 9999 20247
rect 9999 20213 10008 20247
rect 9956 20204 10008 20213
rect 10048 20204 10100 20256
rect 10508 20204 10560 20256
rect 11152 20204 11204 20256
rect 11888 20204 11940 20256
rect 12348 20247 12400 20256
rect 12348 20213 12357 20247
rect 12357 20213 12391 20247
rect 12391 20213 12400 20247
rect 12348 20204 12400 20213
rect 12624 20204 12676 20256
rect 14004 20272 14056 20324
rect 14096 20204 14148 20256
rect 14280 20272 14332 20324
rect 14832 20272 14884 20324
rect 15476 20315 15528 20324
rect 15476 20281 15485 20315
rect 15485 20281 15519 20315
rect 15519 20281 15528 20315
rect 15476 20272 15528 20281
rect 15844 20315 15896 20324
rect 15844 20281 15853 20315
rect 15853 20281 15887 20315
rect 15887 20281 15896 20315
rect 15844 20272 15896 20281
rect 15936 20272 15988 20324
rect 16212 20272 16264 20324
rect 16672 20315 16724 20324
rect 16672 20281 16681 20315
rect 16681 20281 16715 20315
rect 16715 20281 16724 20315
rect 16672 20272 16724 20281
rect 16028 20204 16080 20256
rect 16764 20204 16816 20256
rect 17684 20315 17736 20324
rect 17684 20281 17693 20315
rect 17693 20281 17727 20315
rect 17727 20281 17736 20315
rect 17684 20272 17736 20281
rect 18144 20272 18196 20324
rect 18420 20349 18429 20383
rect 18429 20349 18463 20383
rect 18463 20349 18472 20383
rect 18420 20340 18472 20349
rect 19616 20340 19668 20392
rect 19708 20340 19760 20392
rect 20720 20340 20772 20392
rect 18604 20315 18656 20324
rect 18604 20281 18613 20315
rect 18613 20281 18647 20315
rect 18647 20281 18656 20315
rect 18604 20272 18656 20281
rect 18972 20315 19024 20324
rect 18696 20204 18748 20256
rect 18972 20281 18981 20315
rect 18981 20281 19015 20315
rect 19015 20281 19024 20315
rect 18972 20272 19024 20281
rect 19156 20315 19208 20324
rect 19156 20281 19165 20315
rect 19165 20281 19199 20315
rect 19199 20281 19208 20315
rect 19156 20272 19208 20281
rect 19248 20204 19300 20256
rect 19432 20272 19484 20324
rect 19800 20204 19852 20256
rect 20444 20272 20496 20324
rect 20996 20315 21048 20324
rect 20996 20281 21005 20315
rect 21005 20281 21039 20315
rect 21039 20281 21048 20315
rect 20996 20272 21048 20281
rect 21180 20315 21232 20324
rect 21180 20281 21189 20315
rect 21189 20281 21223 20315
rect 21223 20281 21232 20315
rect 21180 20272 21232 20281
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 1860 20043 1912 20052
rect 1860 20009 1869 20043
rect 1869 20009 1903 20043
rect 1903 20009 1912 20043
rect 1860 20000 1912 20009
rect 4068 20000 4120 20052
rect 4160 20000 4212 20052
rect 6092 20000 6144 20052
rect 7012 20000 7064 20052
rect 8208 20000 8260 20052
rect 9404 20000 9456 20052
rect 9956 20000 10008 20052
rect 10876 20000 10928 20052
rect 2044 19932 2096 19984
rect 1584 19907 1636 19916
rect 1584 19873 1593 19907
rect 1593 19873 1627 19907
rect 1627 19873 1636 19907
rect 1584 19864 1636 19873
rect 1952 19907 2004 19916
rect 1952 19873 1961 19907
rect 1961 19873 1995 19907
rect 1995 19873 2004 19907
rect 1952 19864 2004 19873
rect 2136 19907 2188 19916
rect 2136 19873 2145 19907
rect 2145 19873 2179 19907
rect 2179 19873 2188 19907
rect 2136 19864 2188 19873
rect 2504 19932 2556 19984
rect 204 19796 256 19848
rect 2688 19796 2740 19848
rect 1400 19771 1452 19780
rect 1400 19737 1409 19771
rect 1409 19737 1443 19771
rect 1443 19737 1452 19771
rect 1400 19728 1452 19737
rect 1768 19728 1820 19780
rect 2596 19771 2648 19780
rect 2596 19737 2605 19771
rect 2605 19737 2639 19771
rect 2639 19737 2648 19771
rect 2596 19728 2648 19737
rect 3424 19864 3476 19916
rect 3516 19864 3568 19916
rect 8668 19932 8720 19984
rect 8852 19932 8904 19984
rect 9312 19932 9364 19984
rect 4252 19864 4304 19916
rect 8576 19907 8628 19916
rect 8576 19873 8585 19907
rect 8585 19873 8619 19907
rect 8619 19873 8628 19907
rect 8576 19864 8628 19873
rect 8760 19864 8812 19916
rect 9036 19864 9088 19916
rect 9220 19864 9272 19916
rect 10600 19932 10652 19984
rect 12440 19932 12492 19984
rect 12716 20000 12768 20052
rect 14188 20000 14240 20052
rect 15200 20000 15252 20052
rect 15844 20000 15896 20052
rect 16856 20000 16908 20052
rect 10692 19864 10744 19916
rect 2964 19728 3016 19780
rect 3424 19771 3476 19780
rect 3424 19737 3433 19771
rect 3433 19737 3467 19771
rect 3467 19737 3476 19771
rect 3424 19728 3476 19737
rect 3792 19728 3844 19780
rect 4068 19771 4120 19780
rect 4068 19737 4077 19771
rect 4077 19737 4111 19771
rect 4111 19737 4120 19771
rect 4068 19728 4120 19737
rect 4252 19728 4304 19780
rect 2780 19660 2832 19712
rect 6920 19728 6972 19780
rect 9128 19728 9180 19780
rect 9496 19728 9548 19780
rect 11244 19796 11296 19848
rect 11796 19839 11848 19848
rect 11796 19805 11805 19839
rect 11805 19805 11839 19839
rect 11839 19805 11848 19839
rect 11796 19796 11848 19805
rect 12808 19907 12860 19916
rect 12808 19873 12817 19907
rect 12817 19873 12851 19907
rect 12851 19873 12860 19907
rect 12808 19864 12860 19873
rect 17224 19975 17276 19984
rect 13636 19907 13688 19916
rect 13636 19873 13645 19907
rect 13645 19873 13679 19907
rect 13679 19873 13688 19907
rect 13636 19864 13688 19873
rect 14740 19907 14792 19916
rect 14740 19873 14749 19907
rect 14749 19873 14783 19907
rect 14783 19873 14792 19907
rect 14740 19864 14792 19873
rect 14832 19864 14884 19916
rect 15384 19864 15436 19916
rect 16120 19907 16172 19916
rect 16120 19873 16129 19907
rect 16129 19873 16163 19907
rect 16163 19873 16172 19907
rect 16120 19864 16172 19873
rect 16396 19907 16448 19916
rect 16396 19873 16405 19907
rect 16405 19873 16439 19907
rect 16439 19873 16448 19907
rect 16396 19864 16448 19873
rect 16488 19864 16540 19916
rect 17224 19941 17233 19975
rect 17233 19941 17267 19975
rect 17267 19941 17276 19975
rect 17224 19932 17276 19941
rect 17592 19975 17644 19984
rect 17592 19941 17601 19975
rect 17601 19941 17635 19975
rect 17635 19941 17644 19975
rect 17592 19932 17644 19941
rect 18052 19975 18104 19984
rect 18052 19941 18061 19975
rect 18061 19941 18095 19975
rect 18095 19941 18104 19975
rect 18052 19932 18104 19941
rect 18788 20000 18840 20052
rect 19156 20043 19208 20052
rect 19156 20009 19165 20043
rect 19165 20009 19199 20043
rect 19199 20009 19208 20043
rect 19156 20000 19208 20009
rect 19432 20043 19484 20052
rect 19432 20009 19441 20043
rect 19441 20009 19475 20043
rect 19475 20009 19484 20043
rect 19432 20000 19484 20009
rect 20444 20000 20496 20052
rect 17960 19864 18012 19916
rect 13360 19839 13412 19848
rect 4896 19660 4948 19712
rect 6276 19660 6328 19712
rect 8852 19660 8904 19712
rect 9956 19660 10008 19712
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 14556 19728 14608 19780
rect 14832 19728 14884 19780
rect 15568 19796 15620 19848
rect 17132 19796 17184 19848
rect 16672 19728 16724 19780
rect 12992 19660 13044 19712
rect 14004 19703 14056 19712
rect 14004 19669 14013 19703
rect 14013 19669 14047 19703
rect 14047 19669 14056 19703
rect 14004 19660 14056 19669
rect 14096 19660 14148 19712
rect 14924 19660 14976 19712
rect 15108 19703 15160 19712
rect 15108 19669 15117 19703
rect 15117 19669 15151 19703
rect 15151 19669 15160 19703
rect 15108 19660 15160 19669
rect 15292 19660 15344 19712
rect 18052 19728 18104 19780
rect 19064 19932 19116 19984
rect 20628 19975 20680 19984
rect 18880 19907 18932 19916
rect 18880 19873 18889 19907
rect 18889 19873 18923 19907
rect 18923 19873 18932 19907
rect 18880 19864 18932 19873
rect 19156 19864 19208 19916
rect 19248 19907 19300 19916
rect 19248 19873 19257 19907
rect 19257 19873 19291 19907
rect 19291 19873 19300 19907
rect 19248 19864 19300 19873
rect 19616 19864 19668 19916
rect 19984 19907 20036 19916
rect 19984 19873 19993 19907
rect 19993 19873 20027 19907
rect 20027 19873 20036 19907
rect 19984 19864 20036 19873
rect 20352 19907 20404 19916
rect 20352 19873 20361 19907
rect 20361 19873 20395 19907
rect 20395 19873 20404 19907
rect 20352 19864 20404 19873
rect 20628 19941 20637 19975
rect 20637 19941 20671 19975
rect 20671 19941 20680 19975
rect 20628 19932 20680 19941
rect 20904 19932 20956 19984
rect 20812 19907 20864 19916
rect 20812 19873 20821 19907
rect 20821 19873 20855 19907
rect 20855 19873 20864 19907
rect 20812 19864 20864 19873
rect 21088 19864 21140 19916
rect 20904 19796 20956 19848
rect 17132 19703 17184 19712
rect 17132 19669 17141 19703
rect 17141 19669 17175 19703
rect 17175 19669 17184 19703
rect 17132 19660 17184 19669
rect 17684 19660 17736 19712
rect 18788 19660 18840 19712
rect 18880 19660 18932 19712
rect 19524 19660 19576 19712
rect 20996 19728 21048 19780
rect 21548 19771 21600 19780
rect 21548 19737 21557 19771
rect 21557 19737 21591 19771
rect 21591 19737 21600 19771
rect 21548 19728 21600 19737
rect 20260 19660 20312 19712
rect 21916 19660 21968 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1952 19456 2004 19508
rect 3056 19456 3108 19508
rect 3240 19456 3292 19508
rect 3424 19456 3476 19508
rect 5448 19456 5500 19508
rect 9496 19456 9548 19508
rect 10600 19499 10652 19508
rect 10600 19465 10609 19499
rect 10609 19465 10643 19499
rect 10643 19465 10652 19499
rect 10600 19456 10652 19465
rect 11704 19456 11756 19508
rect 12900 19456 12952 19508
rect 15292 19456 15344 19508
rect 15476 19456 15528 19508
rect 17132 19456 17184 19508
rect 18788 19499 18840 19508
rect 1584 19388 1636 19440
rect 2688 19388 2740 19440
rect 4068 19388 4120 19440
rect 8116 19388 8168 19440
rect 12072 19388 12124 19440
rect 14648 19388 14700 19440
rect 2136 19320 2188 19372
rect 3240 19320 3292 19372
rect 3700 19320 3752 19372
rect 7748 19320 7800 19372
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 1768 19295 1820 19304
rect 1768 19261 1777 19295
rect 1777 19261 1811 19295
rect 1811 19261 1820 19295
rect 1768 19252 1820 19261
rect 2044 19184 2096 19236
rect 2412 19252 2464 19304
rect 2688 19252 2740 19304
rect 3056 19252 3108 19304
rect 3516 19295 3568 19304
rect 3516 19261 3525 19295
rect 3525 19261 3559 19295
rect 3559 19261 3568 19295
rect 3516 19252 3568 19261
rect 3608 19295 3660 19304
rect 3608 19261 3617 19295
rect 3617 19261 3651 19295
rect 3651 19261 3660 19295
rect 3976 19295 4028 19304
rect 3608 19252 3660 19261
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 1952 19159 2004 19168
rect 1952 19125 1961 19159
rect 1961 19125 1995 19159
rect 1995 19125 2004 19159
rect 1952 19116 2004 19125
rect 2964 19116 3016 19168
rect 5908 19184 5960 19236
rect 6460 19252 6512 19304
rect 9128 19295 9180 19304
rect 9128 19261 9137 19295
rect 9137 19261 9171 19295
rect 9171 19261 9180 19295
rect 9128 19252 9180 19261
rect 11244 19320 11296 19372
rect 11704 19320 11756 19372
rect 14924 19388 14976 19440
rect 16120 19388 16172 19440
rect 18144 19388 18196 19440
rect 18788 19465 18797 19499
rect 18797 19465 18831 19499
rect 18831 19465 18840 19499
rect 18788 19456 18840 19465
rect 19616 19456 19668 19508
rect 19432 19388 19484 19440
rect 20352 19388 20404 19440
rect 18236 19320 18288 19372
rect 18604 19320 18656 19372
rect 19248 19320 19300 19372
rect 19800 19320 19852 19372
rect 3700 19116 3752 19168
rect 3976 19116 4028 19168
rect 6092 19159 6144 19168
rect 6092 19125 6101 19159
rect 6101 19125 6135 19159
rect 6135 19125 6144 19159
rect 6092 19116 6144 19125
rect 10784 19252 10836 19304
rect 13452 19295 13504 19304
rect 13452 19261 13486 19295
rect 13486 19261 13504 19295
rect 9496 19227 9548 19236
rect 9496 19193 9530 19227
rect 9530 19193 9548 19227
rect 9496 19184 9548 19193
rect 10692 19159 10744 19168
rect 10692 19125 10701 19159
rect 10701 19125 10735 19159
rect 10735 19125 10744 19159
rect 11704 19159 11756 19168
rect 10692 19116 10744 19125
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 12808 19227 12860 19236
rect 12808 19193 12826 19227
rect 12826 19193 12860 19227
rect 13452 19252 13504 19261
rect 13912 19252 13964 19304
rect 14188 19252 14240 19304
rect 15108 19252 15160 19304
rect 12808 19184 12860 19193
rect 13820 19184 13872 19236
rect 14832 19184 14884 19236
rect 13728 19116 13780 19168
rect 13912 19116 13964 19168
rect 16304 19295 16356 19304
rect 16304 19261 16313 19295
rect 16313 19261 16347 19295
rect 16347 19261 16356 19295
rect 16304 19252 16356 19261
rect 16672 19252 16724 19304
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 18144 19252 18196 19304
rect 18972 19295 19024 19304
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 19064 19252 19116 19304
rect 19984 19252 20036 19304
rect 20904 19252 20956 19304
rect 21088 19252 21140 19304
rect 21548 19295 21600 19304
rect 21548 19261 21557 19295
rect 21557 19261 21591 19295
rect 21591 19261 21600 19295
rect 21548 19252 21600 19261
rect 15292 19184 15344 19236
rect 15660 19159 15712 19168
rect 15660 19125 15669 19159
rect 15669 19125 15703 19159
rect 15703 19125 15712 19159
rect 15660 19116 15712 19125
rect 16028 19116 16080 19168
rect 17776 19184 17828 19236
rect 16672 19159 16724 19168
rect 16672 19125 16681 19159
rect 16681 19125 16715 19159
rect 16715 19125 16724 19159
rect 16672 19116 16724 19125
rect 17500 19159 17552 19168
rect 17500 19125 17509 19159
rect 17509 19125 17543 19159
rect 17543 19125 17552 19159
rect 17500 19116 17552 19125
rect 17684 19116 17736 19168
rect 18328 19116 18380 19168
rect 18420 19116 18472 19168
rect 21272 19184 21324 19236
rect 18880 19116 18932 19168
rect 19616 19116 19668 19168
rect 19892 19159 19944 19168
rect 19892 19125 19901 19159
rect 19901 19125 19935 19159
rect 19935 19125 19944 19159
rect 19892 19116 19944 19125
rect 19984 19116 20036 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 20996 19116 21048 19168
rect 22284 19116 22336 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 2504 18955 2556 18964
rect 2504 18921 2513 18955
rect 2513 18921 2547 18955
rect 2547 18921 2556 18955
rect 2504 18912 2556 18921
rect 2872 18912 2924 18964
rect 3148 18912 3200 18964
rect 3608 18912 3660 18964
rect 3884 18912 3936 18964
rect 6092 18912 6144 18964
rect 6460 18955 6512 18964
rect 6460 18921 6469 18955
rect 6469 18921 6503 18955
rect 6503 18921 6512 18955
rect 6460 18912 6512 18921
rect 8576 18912 8628 18964
rect 10692 18912 10744 18964
rect 11796 18912 11848 18964
rect 12440 18912 12492 18964
rect 14740 18912 14792 18964
rect 15936 18912 15988 18964
rect 17592 18912 17644 18964
rect 18144 18912 18196 18964
rect 3332 18844 3384 18896
rect 3700 18844 3752 18896
rect 5724 18844 5776 18896
rect 5908 18844 5960 18896
rect 8852 18844 8904 18896
rect 9588 18844 9640 18896
rect 11060 18844 11112 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 1768 18819 1820 18828
rect 1768 18785 1777 18819
rect 1777 18785 1811 18819
rect 1811 18785 1820 18819
rect 1768 18776 1820 18785
rect 2136 18776 2188 18828
rect 2320 18819 2372 18828
rect 2320 18785 2329 18819
rect 2329 18785 2363 18819
rect 2363 18785 2372 18819
rect 2320 18776 2372 18785
rect 1676 18708 1728 18760
rect 5356 18776 5408 18828
rect 7012 18776 7064 18828
rect 8300 18776 8352 18828
rect 2688 18708 2740 18760
rect 3332 18708 3384 18760
rect 3516 18708 3568 18760
rect 9220 18776 9272 18828
rect 9496 18776 9548 18828
rect 9956 18819 10008 18828
rect 9588 18751 9640 18760
rect 9588 18717 9597 18751
rect 9597 18717 9631 18751
rect 9631 18717 9640 18751
rect 9588 18708 9640 18717
rect 9956 18785 9965 18819
rect 9965 18785 9999 18819
rect 9999 18785 10008 18819
rect 9956 18776 10008 18785
rect 14372 18844 14424 18896
rect 14648 18887 14700 18896
rect 14648 18853 14682 18887
rect 14682 18853 14700 18887
rect 14648 18844 14700 18853
rect 2228 18683 2280 18692
rect 2228 18649 2237 18683
rect 2237 18649 2271 18683
rect 2271 18649 2280 18683
rect 2228 18640 2280 18649
rect 2964 18683 3016 18692
rect 2964 18649 2973 18683
rect 2973 18649 3007 18683
rect 3007 18649 3016 18683
rect 2964 18640 3016 18649
rect 8392 18640 8444 18692
rect 12440 18776 12492 18828
rect 12900 18776 12952 18828
rect 13176 18776 13228 18828
rect 10692 18751 10744 18760
rect 10692 18717 10701 18751
rect 10701 18717 10735 18751
rect 10735 18717 10744 18751
rect 10692 18708 10744 18717
rect 11796 18708 11848 18760
rect 12256 18708 12308 18760
rect 12808 18751 12860 18760
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 13728 18776 13780 18828
rect 16672 18844 16724 18896
rect 18512 18844 18564 18896
rect 18880 18844 18932 18896
rect 19432 18844 19484 18896
rect 19616 18844 19668 18896
rect 19800 18844 19852 18896
rect 15936 18776 15988 18828
rect 16856 18776 16908 18828
rect 17684 18776 17736 18828
rect 18236 18819 18288 18828
rect 18236 18785 18270 18819
rect 18270 18785 18288 18819
rect 18236 18776 18288 18785
rect 18788 18776 18840 18828
rect 20812 18776 20864 18828
rect 21364 18819 21416 18828
rect 21364 18785 21373 18819
rect 21373 18785 21407 18819
rect 21407 18785 21416 18819
rect 21364 18776 21416 18785
rect 21548 18819 21600 18828
rect 21548 18785 21557 18819
rect 21557 18785 21591 18819
rect 21591 18785 21600 18819
rect 21548 18776 21600 18785
rect 2412 18572 2464 18624
rect 3148 18572 3200 18624
rect 3332 18615 3384 18624
rect 3332 18581 3341 18615
rect 3341 18581 3375 18615
rect 3375 18581 3384 18615
rect 3332 18572 3384 18581
rect 4068 18572 4120 18624
rect 8668 18572 8720 18624
rect 9220 18572 9272 18624
rect 9496 18572 9548 18624
rect 14188 18708 14240 18760
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 15844 18751 15896 18760
rect 15844 18717 15853 18751
rect 15853 18717 15887 18751
rect 15887 18717 15896 18751
rect 15844 18708 15896 18717
rect 16948 18708 17000 18760
rect 15752 18615 15804 18624
rect 15752 18581 15761 18615
rect 15761 18581 15795 18615
rect 15795 18581 15804 18615
rect 15752 18572 15804 18581
rect 16580 18572 16632 18624
rect 17316 18572 17368 18624
rect 19616 18572 19668 18624
rect 19800 18572 19852 18624
rect 21088 18615 21140 18624
rect 21088 18581 21097 18615
rect 21097 18581 21131 18615
rect 21131 18581 21140 18615
rect 21088 18572 21140 18581
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 1492 18411 1544 18420
rect 1492 18377 1501 18411
rect 1501 18377 1535 18411
rect 1535 18377 1544 18411
rect 1492 18368 1544 18377
rect 1584 18368 1636 18420
rect 3148 18368 3200 18420
rect 5356 18411 5408 18420
rect 5356 18377 5365 18411
rect 5365 18377 5399 18411
rect 5399 18377 5408 18411
rect 5356 18368 5408 18377
rect 7656 18368 7708 18420
rect 8300 18411 8352 18420
rect 2044 18300 2096 18352
rect 5632 18300 5684 18352
rect 8300 18377 8309 18411
rect 8309 18377 8343 18411
rect 8343 18377 8352 18411
rect 8300 18368 8352 18377
rect 8392 18368 8444 18420
rect 12256 18368 12308 18420
rect 12532 18300 12584 18352
rect 12716 18368 12768 18420
rect 15844 18368 15896 18420
rect 16948 18368 17000 18420
rect 18144 18368 18196 18420
rect 19340 18368 19392 18420
rect 21364 18368 21416 18420
rect 13820 18300 13872 18352
rect 1768 18232 1820 18284
rect 1584 18139 1636 18148
rect 1584 18105 1593 18139
rect 1593 18105 1627 18139
rect 1627 18105 1636 18139
rect 1584 18096 1636 18105
rect 1952 18139 2004 18148
rect 1952 18105 1961 18139
rect 1961 18105 1995 18139
rect 1995 18105 2004 18139
rect 1952 18096 2004 18105
rect 2596 18207 2648 18216
rect 2596 18173 2605 18207
rect 2605 18173 2639 18207
rect 2639 18173 2648 18207
rect 2596 18164 2648 18173
rect 7564 18232 7616 18284
rect 7932 18232 7984 18284
rect 10416 18275 10468 18284
rect 10416 18241 10425 18275
rect 10425 18241 10459 18275
rect 10459 18241 10468 18275
rect 10416 18232 10468 18241
rect 10600 18275 10652 18284
rect 10600 18241 10609 18275
rect 10609 18241 10643 18275
rect 10643 18241 10652 18275
rect 10600 18232 10652 18241
rect 10784 18232 10836 18284
rect 11612 18232 11664 18284
rect 13084 18232 13136 18284
rect 14188 18300 14240 18352
rect 18052 18300 18104 18352
rect 18788 18300 18840 18352
rect 14004 18232 14056 18284
rect 14372 18232 14424 18284
rect 3148 18164 3200 18216
rect 5172 18207 5224 18216
rect 5172 18173 5181 18207
rect 5181 18173 5215 18207
rect 5215 18173 5224 18207
rect 5172 18164 5224 18173
rect 4988 18096 5040 18148
rect 1860 18071 1912 18080
rect 1860 18037 1869 18071
rect 1869 18037 1903 18071
rect 1903 18037 1912 18071
rect 1860 18028 1912 18037
rect 3240 18028 3292 18080
rect 7288 18164 7340 18216
rect 7472 18164 7524 18216
rect 8668 18164 8720 18216
rect 14280 18164 14332 18216
rect 15752 18232 15804 18284
rect 16948 18275 17000 18284
rect 19800 18300 19852 18352
rect 16948 18241 16964 18275
rect 16964 18241 16998 18275
rect 16998 18241 17000 18275
rect 16948 18232 17000 18241
rect 19248 18275 19300 18284
rect 19248 18241 19257 18275
rect 19257 18241 19291 18275
rect 19291 18241 19300 18275
rect 19248 18232 19300 18241
rect 20352 18300 20404 18352
rect 21548 18343 21600 18352
rect 21548 18309 21557 18343
rect 21557 18309 21591 18343
rect 21591 18309 21600 18343
rect 21548 18300 21600 18309
rect 15660 18164 15712 18216
rect 7656 18139 7708 18148
rect 7656 18105 7665 18139
rect 7665 18105 7699 18139
rect 7699 18105 7708 18139
rect 7656 18096 7708 18105
rect 8852 18096 8904 18148
rect 9956 18096 10008 18148
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 8300 18028 8352 18080
rect 8392 18028 8444 18080
rect 10140 18028 10192 18080
rect 10784 18028 10836 18080
rect 13820 18096 13872 18148
rect 14188 18096 14240 18148
rect 14648 18096 14700 18148
rect 14740 18096 14792 18148
rect 18880 18164 18932 18216
rect 12072 18071 12124 18080
rect 12072 18037 12081 18071
rect 12081 18037 12115 18071
rect 12115 18037 12124 18071
rect 12072 18028 12124 18037
rect 12440 18028 12492 18080
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 13452 18028 13504 18080
rect 17316 18096 17368 18148
rect 15844 18028 15896 18080
rect 16120 18028 16172 18080
rect 16488 18071 16540 18080
rect 16488 18037 16497 18071
rect 16497 18037 16531 18071
rect 16531 18037 16540 18071
rect 16488 18028 16540 18037
rect 16580 18028 16632 18080
rect 19892 18164 19944 18216
rect 19984 18207 20036 18216
rect 19984 18173 19993 18207
rect 19993 18173 20027 18207
rect 20027 18173 20036 18207
rect 19984 18164 20036 18173
rect 20352 18207 20404 18216
rect 20352 18173 20361 18207
rect 20361 18173 20395 18207
rect 20395 18173 20404 18207
rect 20628 18207 20680 18216
rect 20352 18164 20404 18173
rect 20628 18173 20637 18207
rect 20637 18173 20671 18207
rect 20671 18173 20680 18207
rect 20628 18164 20680 18173
rect 18420 18071 18472 18080
rect 18420 18037 18429 18071
rect 18429 18037 18463 18071
rect 18463 18037 18472 18071
rect 20444 18096 20496 18148
rect 21180 18139 21232 18148
rect 21180 18105 21189 18139
rect 21189 18105 21223 18139
rect 21223 18105 21232 18139
rect 21180 18096 21232 18105
rect 18420 18028 18472 18037
rect 19432 18028 19484 18080
rect 19984 18028 20036 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 2596 17824 2648 17876
rect 1860 17688 1912 17740
rect 6460 17824 6512 17876
rect 7288 17824 7340 17876
rect 7472 17867 7524 17876
rect 7472 17833 7481 17867
rect 7481 17833 7515 17867
rect 7515 17833 7524 17867
rect 7472 17824 7524 17833
rect 7748 17824 7800 17876
rect 10968 17824 11020 17876
rect 11060 17824 11112 17876
rect 11612 17824 11664 17876
rect 12072 17824 12124 17876
rect 14556 17824 14608 17876
rect 16120 17824 16172 17876
rect 16396 17824 16448 17876
rect 17500 17824 17552 17876
rect 17776 17867 17828 17876
rect 17776 17833 17785 17867
rect 17785 17833 17819 17867
rect 17819 17833 17828 17867
rect 17776 17824 17828 17833
rect 18420 17824 18472 17876
rect 18972 17824 19024 17876
rect 5356 17756 5408 17808
rect 5540 17756 5592 17808
rect 6184 17688 6236 17740
rect 6920 17756 6972 17808
rect 6920 17663 6972 17672
rect 6920 17629 6929 17663
rect 6929 17629 6963 17663
rect 6963 17629 6972 17663
rect 6920 17620 6972 17629
rect 7104 17731 7156 17740
rect 7104 17697 7113 17731
rect 7113 17697 7147 17731
rect 7147 17697 7156 17731
rect 7104 17688 7156 17697
rect 7748 17688 7800 17740
rect 12900 17756 12952 17808
rect 10416 17688 10468 17740
rect 3516 17552 3568 17604
rect 4068 17552 4120 17604
rect 9128 17620 9180 17672
rect 12716 17688 12768 17740
rect 16856 17756 16908 17808
rect 18604 17756 18656 17808
rect 19984 17756 20036 17808
rect 21088 17799 21140 17808
rect 21088 17765 21097 17799
rect 21097 17765 21131 17799
rect 21131 17765 21140 17799
rect 21088 17756 21140 17765
rect 14280 17688 14332 17740
rect 15384 17688 15436 17740
rect 17868 17688 17920 17740
rect 8208 17552 8260 17604
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 3884 17484 3936 17536
rect 6092 17484 6144 17536
rect 6552 17527 6604 17536
rect 6552 17493 6561 17527
rect 6561 17493 6595 17527
rect 6595 17493 6604 17527
rect 6552 17484 6604 17493
rect 8300 17484 8352 17536
rect 10692 17484 10744 17536
rect 11244 17552 11296 17604
rect 14096 17620 14148 17672
rect 11612 17552 11664 17604
rect 14372 17552 14424 17604
rect 14740 17620 14792 17672
rect 15936 17620 15988 17672
rect 16580 17552 16632 17604
rect 17224 17663 17276 17672
rect 17224 17629 17233 17663
rect 17233 17629 17267 17663
rect 17267 17629 17276 17663
rect 17224 17620 17276 17629
rect 17684 17620 17736 17672
rect 19156 17688 19208 17740
rect 19432 17731 19484 17740
rect 19432 17697 19441 17731
rect 19441 17697 19475 17731
rect 19475 17697 19484 17731
rect 19432 17688 19484 17697
rect 17316 17552 17368 17604
rect 16212 17484 16264 17536
rect 16488 17527 16540 17536
rect 16488 17493 16497 17527
rect 16497 17493 16531 17527
rect 16531 17493 16540 17527
rect 16488 17484 16540 17493
rect 16856 17484 16908 17536
rect 18144 17484 18196 17536
rect 20352 17663 20404 17672
rect 20352 17629 20361 17663
rect 20361 17629 20395 17663
rect 20395 17629 20404 17663
rect 20352 17620 20404 17629
rect 20904 17688 20956 17740
rect 21088 17620 21140 17672
rect 20628 17552 20680 17604
rect 21548 17595 21600 17604
rect 21548 17561 21557 17595
rect 21557 17561 21591 17595
rect 21591 17561 21600 17595
rect 21548 17552 21600 17561
rect 19156 17484 19208 17536
rect 20996 17527 21048 17536
rect 20996 17493 21005 17527
rect 21005 17493 21039 17527
rect 21039 17493 21048 17527
rect 20996 17484 21048 17493
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 1952 17280 2004 17332
rect 1584 17212 1636 17264
rect 3884 17280 3936 17332
rect 2872 17144 2924 17196
rect 5172 17280 5224 17332
rect 6920 17280 6972 17332
rect 5356 17255 5408 17264
rect 5356 17221 5365 17255
rect 5365 17221 5399 17255
rect 5399 17221 5408 17255
rect 5356 17212 5408 17221
rect 5816 17212 5868 17264
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6460 17212 6512 17264
rect 6828 17212 6880 17264
rect 8576 17280 8628 17332
rect 10416 17280 10468 17332
rect 10784 17280 10836 17332
rect 11244 17280 11296 17332
rect 13912 17280 13964 17332
rect 14372 17280 14424 17332
rect 15384 17280 15436 17332
rect 16304 17280 16356 17332
rect 17132 17280 17184 17332
rect 17592 17280 17644 17332
rect 19064 17280 19116 17332
rect 20444 17280 20496 17332
rect 6000 17144 6052 17153
rect 3792 17076 3844 17128
rect 3884 17076 3936 17128
rect 1400 17051 1452 17060
rect 1400 17017 1409 17051
rect 1409 17017 1443 17051
rect 1443 17017 1452 17051
rect 1400 17008 1452 17017
rect 1584 17051 1636 17060
rect 1584 17017 1593 17051
rect 1593 17017 1627 17051
rect 1627 17017 1636 17051
rect 1584 17008 1636 17017
rect 2964 17008 3016 17060
rect 4344 17008 4396 17060
rect 5816 17051 5868 17060
rect 5816 17017 5825 17051
rect 5825 17017 5859 17051
rect 5859 17017 5868 17051
rect 5816 17008 5868 17017
rect 3332 16983 3384 16992
rect 3332 16949 3341 16983
rect 3341 16949 3375 16983
rect 3375 16949 3384 16983
rect 3332 16940 3384 16949
rect 4160 16940 4212 16992
rect 5540 16940 5592 16992
rect 6184 17076 6236 17128
rect 8300 17076 8352 17128
rect 10784 17144 10836 17196
rect 13268 17187 13320 17196
rect 13268 17153 13277 17187
rect 13277 17153 13311 17187
rect 13311 17153 13320 17187
rect 13268 17144 13320 17153
rect 13544 17144 13596 17196
rect 7564 17008 7616 17060
rect 9404 17076 9456 17128
rect 11612 17076 11664 17128
rect 9128 17008 9180 17060
rect 9588 17008 9640 17060
rect 12716 17008 12768 17060
rect 9772 16940 9824 16992
rect 9864 16983 9916 16992
rect 9864 16949 9873 16983
rect 9873 16949 9907 16983
rect 9907 16949 9916 16983
rect 9864 16940 9916 16949
rect 10140 16940 10192 16992
rect 17224 17212 17276 17264
rect 17868 17255 17920 17264
rect 17868 17221 17877 17255
rect 17877 17221 17911 17255
rect 17911 17221 17920 17255
rect 17868 17212 17920 17221
rect 18052 17255 18104 17264
rect 18052 17221 18061 17255
rect 18061 17221 18095 17255
rect 18095 17221 18104 17255
rect 18052 17212 18104 17221
rect 18604 17212 18656 17264
rect 15292 17144 15344 17196
rect 16212 17144 16264 17196
rect 16488 17076 16540 17128
rect 16580 17119 16632 17128
rect 16580 17085 16589 17119
rect 16589 17085 16623 17119
rect 16623 17085 16632 17119
rect 16580 17076 16632 17085
rect 18696 17076 18748 17128
rect 18972 17119 19024 17128
rect 18972 17085 18981 17119
rect 18981 17085 19015 17119
rect 19015 17085 19024 17119
rect 18972 17076 19024 17085
rect 20996 17119 21048 17128
rect 17132 17008 17184 17060
rect 13728 16940 13780 16992
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 14372 16983 14424 16992
rect 13912 16940 13964 16949
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 14556 16983 14608 16992
rect 14556 16949 14565 16983
rect 14565 16949 14599 16983
rect 14599 16949 14608 16983
rect 14556 16940 14608 16949
rect 14740 16940 14792 16992
rect 15384 16940 15436 16992
rect 17040 16940 17092 16992
rect 17224 16940 17276 16992
rect 17684 16983 17736 16992
rect 17684 16949 17693 16983
rect 17693 16949 17727 16983
rect 17727 16949 17736 16983
rect 17684 16940 17736 16949
rect 18144 17008 18196 17060
rect 19616 17008 19668 17060
rect 19524 16940 19576 16992
rect 19892 16940 19944 16992
rect 20996 17085 21005 17119
rect 21005 17085 21039 17119
rect 21039 17085 21048 17119
rect 20996 17076 21048 17085
rect 21180 17051 21232 17060
rect 21180 17017 21189 17051
rect 21189 17017 21223 17051
rect 21223 17017 21232 17051
rect 21180 17008 21232 17017
rect 21364 17051 21416 17060
rect 21364 17017 21373 17051
rect 21373 17017 21407 17051
rect 21407 17017 21416 17051
rect 21364 17008 21416 17017
rect 20996 16940 21048 16992
rect 21456 16983 21508 16992
rect 21456 16949 21465 16983
rect 21465 16949 21499 16983
rect 21499 16949 21508 16983
rect 21456 16940 21508 16949
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 2964 16736 3016 16788
rect 3332 16736 3384 16788
rect 5724 16736 5776 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1952 16600 2004 16652
rect 2688 16643 2740 16652
rect 2688 16609 2697 16643
rect 2697 16609 2731 16643
rect 2731 16609 2740 16643
rect 2688 16600 2740 16609
rect 3976 16600 4028 16652
rect 3884 16575 3936 16584
rect 3884 16541 3893 16575
rect 3893 16541 3927 16575
rect 3927 16541 3936 16575
rect 3884 16532 3936 16541
rect 3700 16464 3752 16516
rect 6276 16600 6328 16652
rect 6552 16668 6604 16720
rect 9588 16736 9640 16788
rect 9772 16736 9824 16788
rect 10600 16736 10652 16788
rect 11612 16779 11664 16788
rect 11612 16745 11621 16779
rect 11621 16745 11655 16779
rect 11655 16745 11664 16779
rect 11612 16736 11664 16745
rect 12900 16779 12952 16788
rect 12900 16745 12909 16779
rect 12909 16745 12943 16779
rect 12943 16745 12952 16779
rect 12900 16736 12952 16745
rect 13728 16779 13780 16788
rect 7840 16600 7892 16652
rect 9220 16643 9272 16652
rect 6000 16575 6052 16584
rect 6000 16541 6009 16575
rect 6009 16541 6043 16575
rect 6043 16541 6052 16575
rect 6000 16532 6052 16541
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 8116 16575 8168 16584
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 8208 16575 8260 16584
rect 8208 16541 8217 16575
rect 8217 16541 8251 16575
rect 8251 16541 8260 16575
rect 9220 16609 9229 16643
rect 9229 16609 9263 16643
rect 9263 16609 9272 16643
rect 9220 16600 9272 16609
rect 10140 16600 10192 16652
rect 8208 16532 8260 16541
rect 10968 16668 11020 16720
rect 13728 16745 13737 16779
rect 13737 16745 13771 16779
rect 13771 16745 13780 16779
rect 13728 16736 13780 16745
rect 16580 16736 16632 16788
rect 17040 16736 17092 16788
rect 18696 16779 18748 16788
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11244 16600 11296 16609
rect 10600 16532 10652 16584
rect 10784 16532 10836 16584
rect 11060 16575 11112 16584
rect 11060 16541 11069 16575
rect 11069 16541 11103 16575
rect 11103 16541 11112 16575
rect 11060 16532 11112 16541
rect 13084 16600 13136 16652
rect 17132 16668 17184 16720
rect 18052 16668 18104 16720
rect 15384 16600 15436 16652
rect 17316 16643 17368 16652
rect 17316 16609 17325 16643
rect 17325 16609 17359 16643
rect 17359 16609 17368 16643
rect 17316 16600 17368 16609
rect 18696 16745 18705 16779
rect 18705 16745 18739 16779
rect 18739 16745 18748 16779
rect 18696 16736 18748 16745
rect 19156 16736 19208 16788
rect 19616 16779 19668 16788
rect 19616 16745 19625 16779
rect 19625 16745 19659 16779
rect 19659 16745 19668 16779
rect 19616 16736 19668 16745
rect 20720 16736 20772 16788
rect 21088 16779 21140 16788
rect 21088 16745 21097 16779
rect 21097 16745 21131 16779
rect 21131 16745 21140 16779
rect 21088 16736 21140 16745
rect 18880 16668 18932 16720
rect 7564 16507 7616 16516
rect 7564 16473 7573 16507
rect 7573 16473 7607 16507
rect 7607 16473 7616 16507
rect 7564 16464 7616 16473
rect 7656 16507 7708 16516
rect 7656 16473 7665 16507
rect 7665 16473 7699 16507
rect 7699 16473 7708 16507
rect 7656 16464 7708 16473
rect 7840 16464 7892 16516
rect 8392 16464 8444 16516
rect 10232 16464 10284 16516
rect 13820 16532 13872 16584
rect 13912 16532 13964 16584
rect 15936 16532 15988 16584
rect 17500 16575 17552 16584
rect 17500 16541 17509 16575
rect 17509 16541 17543 16575
rect 17543 16541 17552 16575
rect 17500 16532 17552 16541
rect 2044 16439 2096 16448
rect 2044 16405 2053 16439
rect 2053 16405 2087 16439
rect 2087 16405 2096 16439
rect 2044 16396 2096 16405
rect 5264 16439 5316 16448
rect 5264 16405 5273 16439
rect 5273 16405 5307 16439
rect 5307 16405 5316 16439
rect 5264 16396 5316 16405
rect 5356 16439 5408 16448
rect 5356 16405 5365 16439
rect 5365 16405 5399 16439
rect 5399 16405 5408 16439
rect 5356 16396 5408 16405
rect 8116 16396 8168 16448
rect 8484 16396 8536 16448
rect 9128 16396 9180 16448
rect 9956 16396 10008 16448
rect 14280 16396 14332 16448
rect 20352 16600 20404 16652
rect 20904 16600 20956 16652
rect 21548 16643 21600 16652
rect 21548 16609 21557 16643
rect 21557 16609 21591 16643
rect 21591 16609 21600 16643
rect 21548 16600 21600 16609
rect 19616 16532 19668 16584
rect 20996 16575 21048 16584
rect 20996 16541 21005 16575
rect 21005 16541 21039 16575
rect 21039 16541 21048 16575
rect 20996 16532 21048 16541
rect 15752 16439 15804 16448
rect 15752 16405 15761 16439
rect 15761 16405 15795 16439
rect 15795 16405 15804 16439
rect 15752 16396 15804 16405
rect 17408 16396 17460 16448
rect 21732 16396 21784 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 1584 16192 1636 16244
rect 2872 16192 2924 16244
rect 3976 16192 4028 16244
rect 5816 16235 5868 16244
rect 2044 16124 2096 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 2044 15988 2096 16040
rect 2320 15988 2372 16040
rect 3792 16124 3844 16176
rect 5540 16124 5592 16176
rect 5816 16201 5825 16235
rect 5825 16201 5859 16235
rect 5859 16201 5868 16235
rect 5816 16192 5868 16201
rect 7104 16192 7156 16244
rect 10232 16192 10284 16244
rect 11060 16192 11112 16244
rect 8852 16124 8904 16176
rect 9128 16124 9180 16176
rect 4344 16099 4396 16108
rect 4344 16065 4353 16099
rect 4353 16065 4387 16099
rect 4387 16065 4396 16099
rect 4344 16056 4396 16065
rect 5264 16056 5316 16108
rect 7564 16056 7616 16108
rect 8208 16099 8260 16108
rect 8208 16065 8217 16099
rect 8217 16065 8251 16099
rect 8251 16065 8260 16099
rect 8208 16056 8260 16065
rect 3884 15988 3936 16040
rect 4068 15988 4120 16040
rect 4160 15988 4212 16040
rect 5356 15988 5408 16040
rect 1584 15963 1636 15972
rect 1584 15929 1593 15963
rect 1593 15929 1627 15963
rect 1627 15929 1636 15963
rect 1584 15920 1636 15929
rect 3700 15920 3752 15972
rect 3976 15920 4028 15972
rect 8392 15988 8444 16040
rect 9956 16056 10008 16108
rect 1860 15852 1912 15904
rect 5356 15895 5408 15904
rect 5356 15861 5365 15895
rect 5365 15861 5399 15895
rect 5399 15861 5408 15895
rect 5356 15852 5408 15861
rect 5448 15895 5500 15904
rect 5448 15861 5457 15895
rect 5457 15861 5491 15895
rect 5491 15861 5500 15895
rect 6276 15895 6328 15904
rect 5448 15852 5500 15861
rect 6276 15861 6285 15895
rect 6285 15861 6319 15895
rect 6319 15861 6328 15895
rect 6276 15852 6328 15861
rect 7288 15895 7340 15904
rect 7288 15861 7297 15895
rect 7297 15861 7331 15895
rect 7331 15861 7340 15895
rect 7288 15852 7340 15861
rect 8760 15920 8812 15972
rect 9864 15988 9916 16040
rect 10600 15920 10652 15972
rect 13820 16192 13872 16244
rect 16120 16192 16172 16244
rect 16948 16192 17000 16244
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 14740 16056 14792 16108
rect 16396 16056 16448 16108
rect 13912 15988 13964 16040
rect 15752 15988 15804 16040
rect 16488 15988 16540 16040
rect 8208 15852 8260 15904
rect 13268 15920 13320 15972
rect 15292 15920 15344 15972
rect 15476 15920 15528 15972
rect 17592 16056 17644 16108
rect 20352 16124 20404 16176
rect 20996 16056 21048 16108
rect 19340 15988 19392 16040
rect 17500 15920 17552 15972
rect 15660 15852 15712 15904
rect 17408 15852 17460 15904
rect 17592 15852 17644 15904
rect 19708 15920 19760 15972
rect 20352 15920 20404 15972
rect 21088 15895 21140 15904
rect 21088 15861 21097 15895
rect 21097 15861 21131 15895
rect 21131 15861 21140 15895
rect 21088 15852 21140 15861
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 1584 15648 1636 15700
rect 1952 15648 2004 15700
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 3976 15648 4028 15700
rect 4344 15648 4396 15700
rect 5448 15648 5500 15700
rect 7288 15648 7340 15700
rect 8392 15648 8444 15700
rect 8760 15691 8812 15700
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 8852 15648 8904 15700
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 8208 15580 8260 15632
rect 2136 15444 2188 15496
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 13544 15580 13596 15632
rect 14556 15580 14608 15632
rect 4804 15487 4856 15496
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 5540 15444 5592 15496
rect 5632 15487 5684 15496
rect 5632 15453 5641 15487
rect 5641 15453 5675 15487
rect 5675 15453 5684 15487
rect 5632 15444 5684 15453
rect 6000 15444 6052 15496
rect 8208 15444 8260 15496
rect 8392 15487 8444 15496
rect 8392 15453 8401 15487
rect 8401 15453 8435 15487
rect 8435 15453 8444 15487
rect 8392 15444 8444 15453
rect 7288 15376 7340 15428
rect 8300 15376 8352 15428
rect 9128 15444 9180 15496
rect 10784 15487 10836 15496
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 10784 15444 10836 15453
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 11244 15376 11296 15428
rect 5908 15308 5960 15360
rect 6184 15308 6236 15360
rect 8484 15308 8536 15360
rect 8852 15308 8904 15360
rect 10600 15351 10652 15360
rect 10600 15317 10609 15351
rect 10609 15317 10643 15351
rect 10643 15317 10652 15351
rect 13820 15444 13872 15496
rect 16396 15623 16448 15632
rect 16396 15589 16430 15623
rect 16430 15589 16448 15623
rect 16396 15580 16448 15589
rect 17500 15648 17552 15700
rect 19616 15648 19668 15700
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 20352 15691 20404 15700
rect 20352 15657 20361 15691
rect 20361 15657 20395 15691
rect 20395 15657 20404 15691
rect 20352 15648 20404 15657
rect 20904 15648 20956 15700
rect 15292 15487 15344 15496
rect 13544 15376 13596 15428
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 19340 15512 19392 15564
rect 19432 15512 19484 15564
rect 20352 15512 20404 15564
rect 19064 15487 19116 15496
rect 19064 15453 19073 15487
rect 19073 15453 19107 15487
rect 19107 15453 19116 15487
rect 19708 15487 19760 15496
rect 19064 15444 19116 15453
rect 19708 15453 19717 15487
rect 19717 15453 19751 15487
rect 19751 15453 19760 15487
rect 19708 15444 19760 15453
rect 15384 15376 15436 15428
rect 17960 15376 18012 15428
rect 20628 15512 20680 15564
rect 21548 15555 21600 15564
rect 21548 15521 21557 15555
rect 21557 15521 21591 15555
rect 21591 15521 21600 15555
rect 21548 15512 21600 15521
rect 21456 15444 21508 15496
rect 10600 15308 10652 15317
rect 14464 15308 14516 15360
rect 19432 15351 19484 15360
rect 19432 15317 19441 15351
rect 19441 15317 19475 15351
rect 19475 15317 19484 15351
rect 19432 15308 19484 15317
rect 19616 15308 19668 15360
rect 21824 15308 21876 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 1492 15147 1544 15156
rect 1492 15113 1501 15147
rect 1501 15113 1535 15147
rect 1535 15113 1544 15147
rect 1492 15104 1544 15113
rect 5356 15104 5408 15156
rect 5540 15104 5592 15156
rect 6920 15104 6972 15156
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 9220 15104 9272 15156
rect 11980 15104 12032 15156
rect 12256 15104 12308 15156
rect 15660 15104 15712 15156
rect 16488 15104 16540 15156
rect 17316 15104 17368 15156
rect 18052 15104 18104 15156
rect 19892 15104 19944 15156
rect 21364 15104 21416 15156
rect 2872 14968 2924 15020
rect 4068 14900 4120 14952
rect 5908 14900 5960 14952
rect 3332 14807 3384 14816
rect 3332 14773 3341 14807
rect 3341 14773 3375 14807
rect 3375 14773 3384 14807
rect 3884 14832 3936 14884
rect 9956 15036 10008 15088
rect 15384 15036 15436 15088
rect 6828 14968 6880 15020
rect 8300 14968 8352 15020
rect 8852 14968 8904 15020
rect 10784 14968 10836 15020
rect 11060 14968 11112 15020
rect 11980 14968 12032 15020
rect 7196 14900 7248 14952
rect 8208 14900 8260 14952
rect 8668 14900 8720 14952
rect 9772 14900 9824 14952
rect 3332 14764 3384 14773
rect 5632 14764 5684 14816
rect 6000 14764 6052 14816
rect 6460 14807 6512 14816
rect 6460 14773 6469 14807
rect 6469 14773 6503 14807
rect 6503 14773 6512 14807
rect 6460 14764 6512 14773
rect 7656 14764 7708 14816
rect 7748 14764 7800 14816
rect 8208 14764 8260 14816
rect 8392 14832 8444 14884
rect 9404 14832 9456 14884
rect 12164 14900 12216 14952
rect 12808 14968 12860 15020
rect 14004 14968 14056 15020
rect 15752 14968 15804 15020
rect 17592 15011 17644 15020
rect 17592 14977 17601 15011
rect 17601 14977 17635 15011
rect 17635 14977 17644 15011
rect 17592 14968 17644 14977
rect 17960 14968 18012 15020
rect 14556 14900 14608 14952
rect 19064 14900 19116 14952
rect 10876 14832 10928 14884
rect 14740 14832 14792 14884
rect 15384 14832 15436 14884
rect 19708 14900 19760 14952
rect 20812 15036 20864 15088
rect 21180 15079 21232 15088
rect 21180 15045 21189 15079
rect 21189 15045 21223 15079
rect 21223 15045 21232 15079
rect 21180 15036 21232 15045
rect 10600 14807 10652 14816
rect 10600 14773 10609 14807
rect 10609 14773 10643 14807
rect 10643 14773 10652 14807
rect 10600 14764 10652 14773
rect 10968 14764 11020 14816
rect 11704 14764 11756 14816
rect 13544 14764 13596 14816
rect 15660 14764 15712 14816
rect 16304 14764 16356 14816
rect 17224 14764 17276 14816
rect 17500 14807 17552 14816
rect 17500 14773 17509 14807
rect 17509 14773 17543 14807
rect 17543 14773 17552 14807
rect 17500 14764 17552 14773
rect 18144 14764 18196 14816
rect 18972 14764 19024 14816
rect 19340 14764 19392 14816
rect 19708 14764 19760 14816
rect 19892 14764 19944 14816
rect 21364 14875 21416 14884
rect 21364 14841 21373 14875
rect 21373 14841 21407 14875
rect 21407 14841 21416 14875
rect 21364 14832 21416 14841
rect 21548 14875 21600 14884
rect 21548 14841 21557 14875
rect 21557 14841 21591 14875
rect 21591 14841 21600 14875
rect 21548 14832 21600 14841
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 2136 14603 2188 14612
rect 2136 14569 2145 14603
rect 2145 14569 2179 14603
rect 2179 14569 2188 14603
rect 2136 14560 2188 14569
rect 3608 14560 3660 14612
rect 14280 14560 14332 14612
rect 15752 14603 15804 14612
rect 5540 14492 5592 14544
rect 6552 14492 6604 14544
rect 6736 14492 6788 14544
rect 7472 14492 7524 14544
rect 1584 14467 1636 14476
rect 1584 14433 1593 14467
rect 1593 14433 1627 14467
rect 1627 14433 1636 14467
rect 1584 14424 1636 14433
rect 2136 14424 2188 14476
rect 2596 14467 2648 14476
rect 2596 14433 2605 14467
rect 2605 14433 2639 14467
rect 2639 14433 2648 14467
rect 2596 14424 2648 14433
rect 4988 14467 5040 14476
rect 4988 14433 5017 14467
rect 5017 14433 5040 14467
rect 4988 14424 5040 14433
rect 6828 14424 6880 14476
rect 6920 14424 6972 14476
rect 9772 14492 9824 14544
rect 11152 14492 11204 14544
rect 12808 14492 12860 14544
rect 10968 14424 11020 14476
rect 14004 14492 14056 14544
rect 15476 14492 15528 14544
rect 15752 14569 15761 14603
rect 15761 14569 15795 14603
rect 15795 14569 15804 14603
rect 15752 14560 15804 14569
rect 16304 14603 16356 14612
rect 16304 14569 16313 14603
rect 16313 14569 16347 14603
rect 16347 14569 16356 14603
rect 16304 14560 16356 14569
rect 16672 14560 16724 14612
rect 19340 14560 19392 14612
rect 20628 14560 20680 14612
rect 21272 14560 21324 14612
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 3884 14220 3936 14229
rect 5908 14220 5960 14272
rect 8484 14356 8536 14408
rect 8668 14356 8720 14408
rect 9220 14399 9272 14408
rect 9220 14365 9229 14399
rect 9229 14365 9263 14399
rect 9263 14365 9272 14399
rect 9220 14356 9272 14365
rect 13912 14356 13964 14408
rect 16580 14424 16632 14476
rect 17500 14492 17552 14544
rect 19708 14492 19760 14544
rect 16304 14356 16356 14408
rect 19432 14424 19484 14476
rect 19984 14492 20036 14544
rect 20076 14467 20128 14476
rect 20076 14433 20085 14467
rect 20085 14433 20119 14467
rect 20119 14433 20128 14467
rect 20076 14424 20128 14433
rect 20168 14424 20220 14476
rect 20996 14467 21048 14476
rect 20996 14433 21005 14467
rect 21005 14433 21039 14467
rect 21039 14433 21048 14467
rect 20996 14424 21048 14433
rect 21272 14424 21324 14476
rect 19616 14356 19668 14408
rect 19984 14399 20036 14408
rect 19984 14365 19993 14399
rect 19993 14365 20027 14399
rect 20027 14365 20036 14399
rect 19984 14356 20036 14365
rect 6920 14331 6972 14340
rect 6920 14297 6929 14331
rect 6929 14297 6963 14331
rect 6963 14297 6972 14331
rect 6920 14288 6972 14297
rect 7104 14220 7156 14272
rect 9680 14288 9732 14340
rect 14004 14331 14056 14340
rect 8852 14220 8904 14272
rect 9496 14220 9548 14272
rect 9864 14263 9916 14272
rect 9864 14229 9873 14263
rect 9873 14229 9907 14263
rect 9907 14229 9916 14263
rect 14004 14297 14013 14331
rect 14013 14297 14047 14331
rect 14047 14297 14056 14331
rect 14004 14288 14056 14297
rect 9864 14220 9916 14229
rect 16672 14288 16724 14340
rect 17408 14288 17460 14340
rect 18696 14288 18748 14340
rect 19432 14288 19484 14340
rect 20628 14288 20680 14340
rect 21180 14331 21232 14340
rect 21180 14297 21189 14331
rect 21189 14297 21223 14331
rect 21223 14297 21232 14331
rect 21180 14288 21232 14297
rect 21548 14331 21600 14340
rect 21548 14297 21557 14331
rect 21557 14297 21591 14331
rect 21591 14297 21600 14331
rect 21548 14288 21600 14297
rect 15844 14263 15896 14272
rect 15844 14229 15853 14263
rect 15853 14229 15887 14263
rect 15887 14229 15896 14263
rect 15844 14220 15896 14229
rect 16488 14220 16540 14272
rect 18144 14220 18196 14272
rect 20720 14220 20772 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 2136 14059 2188 14068
rect 2136 14025 2145 14059
rect 2145 14025 2179 14059
rect 2179 14025 2188 14059
rect 2136 14016 2188 14025
rect 1400 13812 1452 13864
rect 1768 13855 1820 13864
rect 1768 13821 1777 13855
rect 1777 13821 1811 13855
rect 1811 13821 1820 13855
rect 1768 13812 1820 13821
rect 2044 13812 2096 13864
rect 2688 14016 2740 14068
rect 4344 14016 4396 14068
rect 4804 14016 4856 14068
rect 8208 14016 8260 14068
rect 3608 13880 3660 13932
rect 3884 13948 3936 14000
rect 3424 13812 3476 13864
rect 4620 13812 4672 13864
rect 4804 13855 4856 13864
rect 4804 13821 4813 13855
rect 4813 13821 4847 13855
rect 4847 13821 4856 13855
rect 4804 13812 4856 13821
rect 1860 13744 1912 13796
rect 2136 13744 2188 13796
rect 6460 13948 6512 14000
rect 7104 13948 7156 14000
rect 6092 13812 6144 13864
rect 1768 13676 1820 13728
rect 4988 13744 5040 13796
rect 5172 13744 5224 13796
rect 6828 13812 6880 13864
rect 8852 13948 8904 14000
rect 9220 13923 9272 13932
rect 4712 13719 4764 13728
rect 4712 13685 4721 13719
rect 4721 13685 4755 13719
rect 4755 13685 4764 13719
rect 4712 13676 4764 13685
rect 8300 13812 8352 13864
rect 8576 13855 8628 13864
rect 8576 13821 8605 13855
rect 8605 13821 8628 13855
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 8576 13812 8628 13821
rect 9128 13812 9180 13864
rect 9588 13812 9640 13864
rect 9864 13880 9916 13932
rect 11796 14016 11848 14068
rect 13544 14059 13596 14068
rect 13544 14025 13553 14059
rect 13553 14025 13587 14059
rect 13587 14025 13596 14059
rect 13544 14016 13596 14025
rect 14740 14016 14792 14068
rect 11060 13880 11112 13932
rect 11152 13855 11204 13864
rect 11152 13821 11161 13855
rect 11161 13821 11195 13855
rect 11195 13821 11204 13855
rect 11152 13812 11204 13821
rect 12808 13880 12860 13932
rect 12992 13880 13044 13932
rect 13544 13880 13596 13932
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 16304 13923 16356 13932
rect 16304 13889 16313 13923
rect 16313 13889 16347 13923
rect 16347 13889 16356 13923
rect 16304 13880 16356 13889
rect 12256 13744 12308 13796
rect 12624 13812 12676 13864
rect 15200 13812 15252 13864
rect 15844 13812 15896 13864
rect 16120 13812 16172 13864
rect 12992 13744 13044 13796
rect 15660 13744 15712 13796
rect 16580 13787 16632 13796
rect 16580 13753 16589 13787
rect 16589 13753 16623 13787
rect 16623 13753 16632 13787
rect 16580 13744 16632 13753
rect 17592 13744 17644 13796
rect 19340 13812 19392 13864
rect 19616 13855 19668 13864
rect 19616 13821 19634 13855
rect 19634 13821 19668 13855
rect 20352 13880 20404 13932
rect 21180 13880 21232 13932
rect 19616 13812 19668 13821
rect 8668 13676 8720 13728
rect 9496 13719 9548 13728
rect 9496 13685 9505 13719
rect 9505 13685 9539 13719
rect 9539 13685 9548 13719
rect 9496 13676 9548 13685
rect 10968 13676 11020 13728
rect 11796 13676 11848 13728
rect 13084 13676 13136 13728
rect 13452 13676 13504 13728
rect 15200 13676 15252 13728
rect 16488 13676 16540 13728
rect 19064 13676 19116 13728
rect 20444 13812 20496 13864
rect 20720 13744 20772 13796
rect 20352 13719 20404 13728
rect 20352 13685 20361 13719
rect 20361 13685 20395 13719
rect 20395 13685 20404 13719
rect 20352 13676 20404 13685
rect 20628 13676 20680 13728
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 4712 13472 4764 13524
rect 7564 13472 7616 13524
rect 7748 13515 7800 13524
rect 7748 13481 7757 13515
rect 7757 13481 7791 13515
rect 7791 13481 7800 13515
rect 7748 13472 7800 13481
rect 8484 13472 8536 13524
rect 1492 13447 1544 13456
rect 1492 13413 1501 13447
rect 1501 13413 1535 13447
rect 1535 13413 1544 13447
rect 1492 13404 1544 13413
rect 1768 13336 1820 13388
rect 2964 13336 3016 13388
rect 4988 13379 5040 13388
rect 4988 13345 4997 13379
rect 4997 13345 5031 13379
rect 5031 13345 5040 13379
rect 4988 13336 5040 13345
rect 5080 13379 5132 13388
rect 5080 13345 5089 13379
rect 5089 13345 5123 13379
rect 5123 13345 5132 13379
rect 5080 13336 5132 13345
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 5816 13336 5868 13388
rect 7564 13336 7616 13388
rect 3608 13132 3660 13184
rect 6920 13268 6972 13320
rect 8576 13268 8628 13320
rect 9588 13311 9640 13320
rect 9588 13277 9597 13311
rect 9597 13277 9631 13311
rect 9631 13277 9640 13311
rect 9588 13268 9640 13277
rect 10784 13336 10836 13388
rect 13360 13336 13412 13388
rect 13084 13268 13136 13320
rect 13636 13268 13688 13320
rect 15476 13404 15528 13456
rect 15752 13404 15804 13456
rect 19616 13472 19668 13524
rect 20076 13472 20128 13524
rect 20628 13515 20680 13524
rect 20628 13481 20637 13515
rect 20637 13481 20671 13515
rect 20671 13481 20680 13515
rect 20628 13472 20680 13481
rect 21364 13472 21416 13524
rect 7840 13132 7892 13184
rect 14096 13200 14148 13252
rect 14556 13243 14608 13252
rect 14556 13209 14565 13243
rect 14565 13209 14599 13243
rect 14599 13209 14608 13243
rect 14556 13200 14608 13209
rect 10876 13132 10928 13184
rect 11060 13132 11112 13184
rect 11796 13132 11848 13184
rect 12992 13132 13044 13184
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 18972 13336 19024 13388
rect 20904 13336 20956 13388
rect 21548 13379 21600 13388
rect 21548 13345 21557 13379
rect 21557 13345 21591 13379
rect 21591 13345 21600 13379
rect 21548 13336 21600 13345
rect 20444 13268 20496 13320
rect 14924 13132 14976 13184
rect 16856 13132 16908 13184
rect 19616 13200 19668 13252
rect 20168 13200 20220 13252
rect 21088 13200 21140 13252
rect 21548 13132 21600 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 2136 12928 2188 12980
rect 2596 12928 2648 12980
rect 2780 12928 2832 12980
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 3792 12971 3844 12980
rect 3792 12937 3801 12971
rect 3801 12937 3835 12971
rect 3835 12937 3844 12971
rect 3792 12928 3844 12937
rect 7564 12971 7616 12980
rect 7564 12937 7573 12971
rect 7573 12937 7607 12971
rect 7607 12937 7616 12971
rect 7564 12928 7616 12937
rect 12992 12928 13044 12980
rect 13636 12971 13688 12980
rect 13636 12937 13645 12971
rect 13645 12937 13679 12971
rect 13679 12937 13688 12971
rect 13636 12928 13688 12937
rect 14372 12928 14424 12980
rect 14740 12928 14792 12980
rect 19616 12928 19668 12980
rect 19984 12928 20036 12980
rect 20536 12928 20588 12980
rect 1400 12860 1452 12912
rect 1952 12792 2004 12844
rect 2136 12792 2188 12844
rect 2412 12792 2464 12844
rect 9588 12860 9640 12912
rect 5356 12835 5408 12844
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 6920 12835 6972 12844
rect 6920 12801 6929 12835
rect 6929 12801 6963 12835
rect 6963 12801 6972 12835
rect 6920 12792 6972 12801
rect 9772 12792 9824 12844
rect 11612 12792 11664 12844
rect 13360 12860 13412 12912
rect 16948 12903 17000 12912
rect 16948 12869 16957 12903
rect 16957 12869 16991 12903
rect 16991 12869 17000 12903
rect 16948 12860 17000 12869
rect 18328 12860 18380 12912
rect 20628 12860 20680 12912
rect 14372 12792 14424 12844
rect 14924 12792 14976 12844
rect 15292 12792 15344 12844
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 2964 12724 3016 12776
rect 3608 12724 3660 12776
rect 3056 12656 3108 12708
rect 5448 12656 5500 12708
rect 2780 12588 2832 12640
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 5080 12631 5132 12640
rect 5080 12597 5089 12631
rect 5089 12597 5123 12631
rect 5123 12597 5132 12631
rect 5080 12588 5132 12597
rect 6552 12588 6604 12640
rect 8760 12724 8812 12776
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 11796 12724 11848 12776
rect 8300 12656 8352 12708
rect 16856 12724 16908 12776
rect 17040 12724 17092 12776
rect 18420 12724 18472 12776
rect 9496 12588 9548 12640
rect 9680 12631 9732 12640
rect 9680 12597 9689 12631
rect 9689 12597 9723 12631
rect 9723 12597 9732 12631
rect 10140 12631 10192 12640
rect 9680 12588 9732 12597
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 14280 12656 14332 12708
rect 20444 12792 20496 12844
rect 20904 12792 20956 12844
rect 21456 12767 21508 12776
rect 21456 12733 21465 12767
rect 21465 12733 21499 12767
rect 21499 12733 21508 12767
rect 21456 12724 21508 12733
rect 20444 12656 20496 12708
rect 14004 12631 14056 12640
rect 14004 12597 14013 12631
rect 14013 12597 14047 12631
rect 14047 12597 14056 12631
rect 14004 12588 14056 12597
rect 15752 12631 15804 12640
rect 15752 12597 15761 12631
rect 15761 12597 15795 12631
rect 15795 12597 15804 12631
rect 15752 12588 15804 12597
rect 18604 12588 18656 12640
rect 18788 12631 18840 12640
rect 18788 12597 18797 12631
rect 18797 12597 18831 12631
rect 18831 12597 18840 12631
rect 18788 12588 18840 12597
rect 18880 12631 18932 12640
rect 18880 12597 18889 12631
rect 18889 12597 18923 12631
rect 18923 12597 18932 12631
rect 18880 12588 18932 12597
rect 19616 12588 19668 12640
rect 20812 12588 20864 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 2136 12384 2188 12436
rect 2320 12384 2372 12436
rect 2872 12384 2924 12436
rect 3424 12384 3476 12436
rect 4712 12384 4764 12436
rect 9772 12384 9824 12436
rect 10048 12384 10100 12436
rect 11612 12384 11664 12436
rect 13820 12384 13872 12436
rect 14004 12384 14056 12436
rect 18788 12384 18840 12436
rect 19156 12384 19208 12436
rect 19616 12384 19668 12436
rect 1676 12316 1728 12368
rect 11060 12316 11112 12368
rect 2688 12291 2740 12300
rect 2688 12257 2706 12291
rect 2706 12257 2740 12291
rect 2688 12248 2740 12257
rect 2872 12248 2924 12300
rect 4344 12291 4396 12300
rect 4344 12257 4353 12291
rect 4353 12257 4387 12291
rect 4387 12257 4396 12291
rect 4344 12248 4396 12257
rect 5172 12291 5224 12300
rect 5172 12257 5206 12291
rect 5206 12257 5224 12291
rect 5172 12248 5224 12257
rect 3976 12180 4028 12232
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 4712 12180 4764 12232
rect 10048 12248 10100 12300
rect 11704 12291 11756 12300
rect 11704 12257 11713 12291
rect 11713 12257 11747 12291
rect 11747 12257 11756 12291
rect 11704 12248 11756 12257
rect 6460 12180 6512 12232
rect 9312 12180 9364 12232
rect 9588 12180 9640 12232
rect 10876 12180 10928 12232
rect 11612 12180 11664 12232
rect 18604 12316 18656 12368
rect 18696 12316 18748 12368
rect 15108 12248 15160 12300
rect 16120 12248 16172 12300
rect 17868 12248 17920 12300
rect 18052 12291 18104 12300
rect 18052 12257 18061 12291
rect 18061 12257 18095 12291
rect 18095 12257 18104 12291
rect 18052 12248 18104 12257
rect 7932 12112 7984 12164
rect 9220 12087 9272 12096
rect 9220 12053 9229 12087
rect 9229 12053 9263 12087
rect 9263 12053 9272 12087
rect 9220 12044 9272 12053
rect 10784 12044 10836 12096
rect 12072 12044 12124 12096
rect 12440 12044 12492 12096
rect 13820 12180 13872 12232
rect 15292 12180 15344 12232
rect 16764 12180 16816 12232
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 18144 12223 18196 12232
rect 18144 12189 18153 12223
rect 18153 12189 18187 12223
rect 18187 12189 18196 12223
rect 18144 12180 18196 12189
rect 18420 12180 18472 12232
rect 18696 12180 18748 12232
rect 19156 12223 19208 12232
rect 19156 12189 19165 12223
rect 19165 12189 19199 12223
rect 19199 12189 19208 12223
rect 19156 12180 19208 12189
rect 19984 12316 20036 12368
rect 20352 12384 20404 12436
rect 20628 12316 20680 12368
rect 20720 12316 20772 12368
rect 20352 12248 20404 12300
rect 21180 12291 21232 12300
rect 21180 12257 21189 12291
rect 21189 12257 21223 12291
rect 21223 12257 21232 12291
rect 21180 12248 21232 12257
rect 21456 12291 21508 12300
rect 21456 12257 21465 12291
rect 21465 12257 21499 12291
rect 21499 12257 21508 12291
rect 21456 12248 21508 12257
rect 13728 12112 13780 12164
rect 19708 12112 19760 12164
rect 13820 12044 13872 12096
rect 14372 12044 14424 12096
rect 15844 12044 15896 12096
rect 16028 12087 16080 12096
rect 16028 12053 16037 12087
rect 16037 12053 16071 12087
rect 16071 12053 16080 12087
rect 16028 12044 16080 12053
rect 16120 12087 16172 12096
rect 16120 12053 16129 12087
rect 16129 12053 16163 12087
rect 16163 12053 16172 12087
rect 16120 12044 16172 12053
rect 19064 12044 19116 12096
rect 20352 12044 20404 12096
rect 20536 12112 20588 12164
rect 21456 12044 21508 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 2688 11840 2740 11892
rect 4896 11840 4948 11892
rect 5448 11840 5500 11892
rect 6000 11840 6052 11892
rect 6276 11840 6328 11892
rect 6552 11883 6604 11892
rect 6552 11849 6561 11883
rect 6561 11849 6595 11883
rect 6595 11849 6604 11883
rect 6552 11840 6604 11849
rect 8392 11840 8444 11892
rect 13452 11840 13504 11892
rect 14096 11883 14148 11892
rect 14096 11849 14105 11883
rect 14105 11849 14139 11883
rect 14139 11849 14148 11883
rect 14096 11840 14148 11849
rect 15476 11840 15528 11892
rect 15844 11840 15896 11892
rect 3056 11815 3108 11824
rect 3056 11781 3065 11815
rect 3065 11781 3099 11815
rect 3099 11781 3108 11815
rect 3056 11772 3108 11781
rect 5172 11772 5224 11824
rect 5356 11815 5408 11824
rect 5356 11781 5365 11815
rect 5365 11781 5399 11815
rect 5399 11781 5408 11815
rect 5356 11772 5408 11781
rect 3516 11704 3568 11756
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 4988 11704 5040 11756
rect 6644 11772 6696 11824
rect 7748 11772 7800 11824
rect 6552 11704 6604 11756
rect 7380 11704 7432 11756
rect 7932 11747 7984 11756
rect 7932 11713 7941 11747
rect 7941 11713 7975 11747
rect 7975 11713 7984 11747
rect 7932 11704 7984 11713
rect 8208 11704 8260 11756
rect 2872 11636 2924 11688
rect 3240 11636 3292 11688
rect 9220 11704 9272 11756
rect 9680 11704 9732 11756
rect 10692 11747 10744 11756
rect 10692 11713 10701 11747
rect 10701 11713 10735 11747
rect 10735 11713 10744 11747
rect 10692 11704 10744 11713
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 11980 11747 12032 11756
rect 10784 11704 10836 11713
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 8484 11679 8536 11688
rect 2412 11568 2464 11620
rect 8484 11645 8493 11679
rect 8493 11645 8527 11679
rect 8527 11645 8536 11679
rect 8484 11636 8536 11645
rect 10508 11636 10560 11688
rect 11704 11636 11756 11688
rect 4436 11568 4488 11620
rect 1400 11543 1452 11552
rect 1400 11509 1409 11543
rect 1409 11509 1443 11543
rect 1443 11509 1452 11543
rect 1400 11500 1452 11509
rect 5448 11543 5500 11552
rect 5448 11509 5457 11543
rect 5457 11509 5491 11543
rect 5491 11509 5500 11543
rect 5816 11543 5868 11552
rect 5448 11500 5500 11509
rect 5816 11509 5825 11543
rect 5825 11509 5859 11543
rect 5859 11509 5868 11543
rect 5816 11500 5868 11509
rect 6920 11543 6972 11552
rect 6920 11509 6929 11543
rect 6929 11509 6963 11543
rect 6963 11509 6972 11543
rect 6920 11500 6972 11509
rect 12440 11568 12492 11620
rect 13820 11636 13872 11688
rect 16028 11772 16080 11824
rect 16764 11840 16816 11892
rect 18604 11840 18656 11892
rect 19524 11840 19576 11892
rect 20996 11840 21048 11892
rect 21732 11840 21784 11892
rect 18512 11772 18564 11824
rect 19064 11772 19116 11824
rect 20904 11772 20956 11824
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 13084 11568 13136 11620
rect 14280 11568 14332 11620
rect 15752 11636 15804 11688
rect 16764 11636 16816 11688
rect 16948 11679 17000 11688
rect 16948 11645 16957 11679
rect 16957 11645 16991 11679
rect 16991 11645 17000 11679
rect 16948 11636 17000 11645
rect 20996 11679 21048 11688
rect 20996 11645 21005 11679
rect 21005 11645 21039 11679
rect 21039 11645 21048 11679
rect 20996 11636 21048 11645
rect 21456 11679 21508 11688
rect 21456 11645 21465 11679
rect 21465 11645 21499 11679
rect 21499 11645 21508 11679
rect 21456 11636 21508 11645
rect 11244 11543 11296 11552
rect 11244 11509 11253 11543
rect 11253 11509 11287 11543
rect 11287 11509 11296 11543
rect 11244 11500 11296 11509
rect 12164 11543 12216 11552
rect 12164 11509 12173 11543
rect 12173 11509 12207 11543
rect 12207 11509 12216 11543
rect 12164 11500 12216 11509
rect 12532 11500 12584 11552
rect 17040 11500 17092 11552
rect 17868 11568 17920 11620
rect 18788 11568 18840 11620
rect 20168 11568 20220 11620
rect 21548 11568 21600 11620
rect 18052 11500 18104 11552
rect 19064 11543 19116 11552
rect 19064 11509 19073 11543
rect 19073 11509 19107 11543
rect 19107 11509 19116 11543
rect 19064 11500 19116 11509
rect 19340 11500 19392 11552
rect 20076 11500 20128 11552
rect 21456 11500 21508 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 1676 11296 1728 11348
rect 1952 11339 2004 11348
rect 1952 11305 1961 11339
rect 1961 11305 1995 11339
rect 1995 11305 2004 11339
rect 1952 11296 2004 11305
rect 4344 11296 4396 11348
rect 5080 11296 5132 11348
rect 5724 11296 5776 11348
rect 6920 11296 6972 11348
rect 8392 11296 8444 11348
rect 9680 11339 9732 11348
rect 9680 11305 9689 11339
rect 9689 11305 9723 11339
rect 9723 11305 9732 11339
rect 9680 11296 9732 11305
rect 10600 11296 10652 11348
rect 3148 11228 3200 11280
rect 5448 11228 5500 11280
rect 7472 11228 7524 11280
rect 1492 11203 1544 11212
rect 1492 11169 1501 11203
rect 1501 11169 1535 11203
rect 1535 11169 1544 11203
rect 1492 11160 1544 11169
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 2872 11160 2924 11212
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 5908 11160 5960 11212
rect 3332 11135 3384 11144
rect 2412 11024 2464 11076
rect 3332 11101 3341 11135
rect 3341 11101 3375 11135
rect 3375 11101 3384 11135
rect 3332 11092 3384 11101
rect 3516 11135 3568 11144
rect 3516 11101 3525 11135
rect 3525 11101 3559 11135
rect 3559 11101 3568 11135
rect 3516 11092 3568 11101
rect 4252 11135 4304 11144
rect 2964 11024 3016 11076
rect 4252 11101 4261 11135
rect 4261 11101 4295 11135
rect 4295 11101 4304 11135
rect 4252 11092 4304 11101
rect 4436 11092 4488 11144
rect 5448 11135 5500 11144
rect 5448 11101 5457 11135
rect 5457 11101 5491 11135
rect 5491 11101 5500 11135
rect 6552 11160 6604 11212
rect 7840 11160 7892 11212
rect 8944 11228 8996 11280
rect 9404 11228 9456 11280
rect 11796 11296 11848 11348
rect 12164 11296 12216 11348
rect 13544 11339 13596 11348
rect 13544 11305 13553 11339
rect 13553 11305 13587 11339
rect 13587 11305 13596 11339
rect 13544 11296 13596 11305
rect 11244 11228 11296 11280
rect 15384 11296 15436 11348
rect 13820 11228 13872 11280
rect 15016 11228 15068 11280
rect 16856 11296 16908 11348
rect 17040 11339 17092 11348
rect 17040 11305 17049 11339
rect 17049 11305 17083 11339
rect 17083 11305 17092 11339
rect 17040 11296 17092 11305
rect 10692 11160 10744 11212
rect 13912 11203 13964 11212
rect 5448 11092 5500 11101
rect 5356 11024 5408 11076
rect 5540 11024 5592 11076
rect 6644 11092 6696 11144
rect 8208 11092 8260 11144
rect 9496 11092 9548 11144
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 12440 11092 12492 11144
rect 13912 11169 13921 11203
rect 13921 11169 13955 11203
rect 13955 11169 13964 11203
rect 13912 11160 13964 11169
rect 14004 11160 14056 11212
rect 14280 11092 14332 11144
rect 14556 11160 14608 11212
rect 18880 11296 18932 11348
rect 19064 11296 19116 11348
rect 19708 11296 19760 11348
rect 19156 11228 19208 11280
rect 19248 11228 19300 11280
rect 19524 11228 19576 11280
rect 20536 11228 20588 11280
rect 21640 11228 21692 11280
rect 14832 11092 14884 11144
rect 8760 11024 8812 11076
rect 4160 10956 4212 11008
rect 6644 10999 6696 11008
rect 6644 10965 6653 10999
rect 6653 10965 6687 10999
rect 6687 10965 6696 10999
rect 6644 10956 6696 10965
rect 9588 10956 9640 11008
rect 11152 10956 11204 11008
rect 12348 11024 12400 11076
rect 17868 11160 17920 11212
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 12440 10956 12492 11008
rect 12900 10956 12952 11008
rect 13820 10956 13872 11008
rect 14832 10999 14884 11008
rect 14832 10965 14841 10999
rect 14841 10965 14875 10999
rect 14875 10965 14884 10999
rect 14832 10956 14884 10965
rect 16856 11092 16908 11144
rect 17592 11092 17644 11144
rect 17776 11092 17828 11144
rect 20352 11160 20404 11212
rect 21548 11160 21600 11212
rect 18696 11067 18748 11076
rect 18696 11033 18705 11067
rect 18705 11033 18739 11067
rect 18739 11033 18748 11067
rect 18696 11024 18748 11033
rect 19984 11092 20036 11144
rect 20720 11092 20772 11144
rect 16764 10956 16816 11008
rect 17132 10999 17184 11008
rect 17132 10965 17141 10999
rect 17141 10965 17175 10999
rect 17175 10965 17184 10999
rect 17132 10956 17184 10965
rect 17592 10956 17644 11008
rect 18880 10956 18932 11008
rect 20904 11024 20956 11076
rect 21916 11024 21968 11076
rect 19708 10956 19760 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 3332 10752 3384 10804
rect 4252 10795 4304 10804
rect 4252 10761 4261 10795
rect 4261 10761 4295 10795
rect 4295 10761 4304 10795
rect 4252 10752 4304 10761
rect 4344 10752 4396 10804
rect 5724 10752 5776 10804
rect 7012 10752 7064 10804
rect 8300 10752 8352 10804
rect 9128 10752 9180 10804
rect 3148 10727 3200 10736
rect 3148 10693 3157 10727
rect 3157 10693 3191 10727
rect 3191 10693 3200 10727
rect 3148 10684 3200 10693
rect 1492 10616 1544 10668
rect 2412 10616 2464 10668
rect 2872 10659 2924 10668
rect 2872 10625 2881 10659
rect 2881 10625 2915 10659
rect 2915 10625 2924 10659
rect 2872 10616 2924 10625
rect 1400 10480 1452 10532
rect 1676 10523 1728 10532
rect 1676 10489 1685 10523
rect 1685 10489 1719 10523
rect 1719 10489 1728 10523
rect 1676 10480 1728 10489
rect 4712 10548 4764 10600
rect 5448 10616 5500 10668
rect 7104 10616 7156 10668
rect 11152 10752 11204 10804
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 11980 10752 12032 10804
rect 10140 10684 10192 10736
rect 10416 10684 10468 10736
rect 5540 10548 5592 10600
rect 7748 10548 7800 10600
rect 8760 10548 8812 10600
rect 4160 10480 4212 10532
rect 4804 10523 4856 10532
rect 4804 10489 4813 10523
rect 4813 10489 4847 10523
rect 4847 10489 4856 10523
rect 4804 10480 4856 10489
rect 7380 10480 7432 10532
rect 9496 10548 9548 10600
rect 9404 10480 9456 10532
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 17224 10752 17276 10804
rect 18144 10752 18196 10804
rect 18972 10752 19024 10804
rect 19064 10752 19116 10804
rect 20168 10795 20220 10804
rect 13084 10684 13136 10736
rect 19708 10684 19760 10736
rect 14280 10659 14332 10668
rect 10600 10616 10652 10625
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 12348 10548 12400 10600
rect 12440 10548 12492 10600
rect 13084 10591 13136 10600
rect 13084 10557 13093 10591
rect 13093 10557 13127 10591
rect 13127 10557 13136 10591
rect 13084 10548 13136 10557
rect 14004 10548 14056 10600
rect 15476 10616 15528 10668
rect 15844 10616 15896 10668
rect 16396 10616 16448 10668
rect 17040 10659 17092 10668
rect 14832 10548 14884 10600
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 17224 10659 17276 10668
rect 17224 10625 17233 10659
rect 17233 10625 17267 10659
rect 17267 10625 17276 10659
rect 17224 10616 17276 10625
rect 18880 10616 18932 10668
rect 19156 10659 19208 10668
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 2320 10455 2372 10464
rect 2320 10421 2329 10455
rect 2329 10421 2363 10455
rect 2363 10421 2372 10455
rect 2320 10412 2372 10421
rect 3792 10455 3844 10464
rect 3792 10421 3801 10455
rect 3801 10421 3835 10455
rect 3835 10421 3844 10455
rect 3792 10412 3844 10421
rect 4896 10412 4948 10464
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 5632 10455 5684 10464
rect 5632 10421 5641 10455
rect 5641 10421 5675 10455
rect 5675 10421 5684 10455
rect 6460 10455 6512 10464
rect 5632 10412 5684 10421
rect 6460 10421 6469 10455
rect 6469 10421 6503 10455
rect 6503 10421 6512 10455
rect 6460 10412 6512 10421
rect 7472 10455 7524 10464
rect 7472 10421 7481 10455
rect 7481 10421 7515 10455
rect 7515 10421 7524 10455
rect 7472 10412 7524 10421
rect 9128 10412 9180 10464
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 9496 10455 9548 10464
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 9956 10412 10008 10464
rect 12900 10480 12952 10532
rect 13268 10480 13320 10532
rect 15476 10480 15528 10532
rect 15936 10480 15988 10532
rect 16948 10480 17000 10532
rect 17132 10548 17184 10600
rect 19340 10548 19392 10600
rect 19524 10548 19576 10600
rect 19616 10591 19668 10600
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 20168 10761 20177 10795
rect 20177 10761 20211 10795
rect 20211 10761 20220 10795
rect 20168 10752 20220 10761
rect 20996 10795 21048 10804
rect 20996 10761 21005 10795
rect 21005 10761 21039 10795
rect 21039 10761 21048 10795
rect 20996 10752 21048 10761
rect 21180 10684 21232 10736
rect 20720 10659 20772 10668
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 20628 10548 20680 10600
rect 20904 10548 20956 10600
rect 21456 10523 21508 10532
rect 21456 10489 21465 10523
rect 21465 10489 21499 10523
rect 21499 10489 21508 10523
rect 21456 10480 21508 10489
rect 12072 10412 12124 10464
rect 13544 10412 13596 10464
rect 13912 10412 13964 10464
rect 14096 10455 14148 10464
rect 14096 10421 14105 10455
rect 14105 10421 14139 10455
rect 14139 10421 14148 10455
rect 14096 10412 14148 10421
rect 14280 10412 14332 10464
rect 15292 10455 15344 10464
rect 15292 10421 15301 10455
rect 15301 10421 15335 10455
rect 15335 10421 15344 10455
rect 15292 10412 15344 10421
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 15752 10412 15804 10421
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 16764 10455 16816 10464
rect 16764 10421 16773 10455
rect 16773 10421 16807 10455
rect 16807 10421 16816 10455
rect 16764 10412 16816 10421
rect 17132 10412 17184 10464
rect 19708 10455 19760 10464
rect 19708 10421 19717 10455
rect 19717 10421 19751 10455
rect 19751 10421 19760 10455
rect 19708 10412 19760 10421
rect 20168 10412 20220 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 1584 10208 1636 10260
rect 2228 10251 2280 10260
rect 2228 10217 2237 10251
rect 2237 10217 2271 10251
rect 2271 10217 2280 10251
rect 2228 10208 2280 10217
rect 3792 10208 3844 10260
rect 5448 10251 5500 10260
rect 5448 10217 5457 10251
rect 5457 10217 5491 10251
rect 5491 10217 5500 10251
rect 5448 10208 5500 10217
rect 8392 10208 8444 10260
rect 9128 10251 9180 10260
rect 9128 10217 9137 10251
rect 9137 10217 9171 10251
rect 9171 10217 9180 10251
rect 9128 10208 9180 10217
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 9588 10251 9640 10260
rect 9588 10217 9597 10251
rect 9597 10217 9631 10251
rect 9631 10217 9640 10251
rect 9588 10208 9640 10217
rect 5540 10140 5592 10192
rect 6644 10140 6696 10192
rect 1492 10115 1544 10124
rect 1492 10081 1501 10115
rect 1501 10081 1535 10115
rect 1535 10081 1544 10115
rect 1492 10072 1544 10081
rect 1952 10115 2004 10124
rect 1952 10081 1961 10115
rect 1961 10081 1995 10115
rect 1995 10081 2004 10115
rect 1952 10072 2004 10081
rect 2044 10115 2096 10124
rect 2044 10081 2053 10115
rect 2053 10081 2087 10115
rect 2087 10081 2096 10115
rect 2044 10072 2096 10081
rect 4804 10072 4856 10124
rect 11704 10140 11756 10192
rect 12532 10208 12584 10260
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 14280 10208 14332 10260
rect 14372 10208 14424 10260
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 5724 10004 5776 10056
rect 8668 10072 8720 10124
rect 12072 10115 12124 10124
rect 12072 10081 12081 10115
rect 12081 10081 12115 10115
rect 12115 10081 12124 10115
rect 12072 10072 12124 10081
rect 12900 10115 12952 10124
rect 12900 10081 12909 10115
rect 12909 10081 12943 10115
rect 12943 10081 12952 10115
rect 12900 10072 12952 10081
rect 1860 9868 1912 9920
rect 7104 9868 7156 9920
rect 8760 10004 8812 10056
rect 9312 10004 9364 10056
rect 9588 9868 9640 9920
rect 9680 9868 9732 9920
rect 12440 10004 12492 10056
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 15752 10140 15804 10192
rect 15936 10208 15988 10260
rect 17592 10251 17644 10260
rect 17132 10140 17184 10192
rect 17592 10217 17601 10251
rect 17601 10217 17635 10251
rect 17635 10217 17644 10251
rect 17592 10208 17644 10217
rect 19616 10251 19668 10260
rect 19616 10217 19625 10251
rect 19625 10217 19659 10251
rect 19659 10217 19668 10251
rect 19616 10208 19668 10217
rect 19340 10140 19392 10192
rect 14188 10072 14240 10124
rect 13544 10004 13596 10056
rect 14372 10004 14424 10056
rect 12992 9936 13044 9988
rect 15568 10072 15620 10124
rect 15844 10115 15896 10124
rect 15844 10081 15862 10115
rect 15862 10081 15896 10115
rect 15844 10072 15896 10081
rect 17224 10072 17276 10124
rect 21272 10208 21324 10260
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 20812 10115 20864 10124
rect 20812 10081 20821 10115
rect 20821 10081 20855 10115
rect 20855 10081 20864 10115
rect 20812 10072 20864 10081
rect 21456 10115 21508 10124
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 19340 10004 19392 10056
rect 20444 10004 20496 10056
rect 13084 9868 13136 9920
rect 20904 9936 20956 9988
rect 21548 9936 21600 9988
rect 18144 9868 18196 9920
rect 20536 9911 20588 9920
rect 20536 9877 20545 9911
rect 20545 9877 20579 9911
rect 20579 9877 20588 9911
rect 20536 9868 20588 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 1952 9664 2004 9716
rect 2136 9639 2188 9648
rect 2136 9605 2145 9639
rect 2145 9605 2179 9639
rect 2179 9605 2188 9639
rect 2136 9596 2188 9605
rect 2320 9596 2372 9648
rect 2780 9528 2832 9580
rect 1584 9460 1636 9512
rect 2596 9503 2648 9512
rect 2596 9469 2605 9503
rect 2605 9469 2639 9503
rect 2639 9469 2648 9503
rect 2596 9460 2648 9469
rect 3148 9503 3200 9512
rect 1492 9435 1544 9444
rect 1492 9401 1501 9435
rect 1501 9401 1535 9435
rect 1535 9401 1544 9435
rect 1492 9392 1544 9401
rect 1860 9435 1912 9444
rect 1860 9401 1869 9435
rect 1869 9401 1903 9435
rect 1903 9401 1912 9435
rect 1860 9392 1912 9401
rect 2872 9324 2924 9376
rect 3148 9469 3157 9503
rect 3157 9469 3191 9503
rect 3191 9469 3200 9503
rect 3148 9460 3200 9469
rect 4344 9664 4396 9716
rect 4528 9571 4580 9580
rect 4528 9537 4537 9571
rect 4537 9537 4571 9571
rect 4571 9537 4580 9571
rect 4988 9664 5040 9716
rect 5632 9596 5684 9648
rect 7472 9664 7524 9716
rect 12532 9664 12584 9716
rect 13176 9664 13228 9716
rect 15108 9664 15160 9716
rect 15292 9664 15344 9716
rect 15568 9664 15620 9716
rect 4528 9528 4580 9537
rect 6736 9596 6788 9648
rect 5908 9460 5960 9512
rect 6184 9528 6236 9580
rect 6368 9528 6420 9580
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 8392 9503 8444 9512
rect 8392 9469 8401 9503
rect 8401 9469 8435 9503
rect 8435 9469 8444 9503
rect 8392 9460 8444 9469
rect 4252 9392 4304 9444
rect 4712 9392 4764 9444
rect 7196 9392 7248 9444
rect 7564 9367 7616 9376
rect 7564 9333 7573 9367
rect 7573 9333 7607 9367
rect 7607 9333 7616 9367
rect 7564 9324 7616 9333
rect 9404 9596 9456 9648
rect 11244 9596 11296 9648
rect 15844 9596 15896 9648
rect 16672 9639 16724 9648
rect 16672 9605 16681 9639
rect 16681 9605 16715 9639
rect 16715 9605 16724 9639
rect 16672 9596 16724 9605
rect 16948 9639 17000 9648
rect 16948 9605 16957 9639
rect 16957 9605 16991 9639
rect 16991 9605 17000 9639
rect 16948 9596 17000 9605
rect 9680 9528 9732 9580
rect 10140 9503 10192 9512
rect 10140 9469 10149 9503
rect 10149 9469 10183 9503
rect 10183 9469 10192 9503
rect 10140 9460 10192 9469
rect 13084 9528 13136 9580
rect 13268 9528 13320 9580
rect 15476 9528 15528 9580
rect 12164 9435 12216 9444
rect 12164 9401 12198 9435
rect 12198 9401 12216 9435
rect 12164 9392 12216 9401
rect 12624 9392 12676 9444
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 12808 9324 12860 9376
rect 16396 9460 16448 9512
rect 16672 9460 16724 9512
rect 19432 9664 19484 9716
rect 20812 9664 20864 9716
rect 21088 9596 21140 9648
rect 21364 9639 21416 9648
rect 21364 9605 21373 9639
rect 21373 9605 21407 9639
rect 21407 9605 21416 9639
rect 21364 9596 21416 9605
rect 20720 9571 20772 9580
rect 20720 9537 20729 9571
rect 20729 9537 20763 9571
rect 20763 9537 20772 9571
rect 20720 9528 20772 9537
rect 21180 9503 21232 9512
rect 21180 9469 21189 9503
rect 21189 9469 21223 9503
rect 21223 9469 21232 9503
rect 21180 9460 21232 9469
rect 21548 9503 21600 9512
rect 21548 9469 21557 9503
rect 21557 9469 21591 9503
rect 21591 9469 21600 9503
rect 21548 9460 21600 9469
rect 14556 9392 14608 9444
rect 15384 9324 15436 9376
rect 16304 9324 16356 9376
rect 17592 9392 17644 9444
rect 19432 9435 19484 9444
rect 18144 9324 18196 9376
rect 18236 9324 18288 9376
rect 19432 9401 19472 9435
rect 19472 9401 19484 9435
rect 19432 9392 19484 9401
rect 20444 9392 20496 9444
rect 19616 9324 19668 9376
rect 20076 9324 20128 9376
rect 20536 9367 20588 9376
rect 20536 9333 20545 9367
rect 20545 9333 20579 9367
rect 20579 9333 20588 9367
rect 20536 9324 20588 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 2596 9120 2648 9172
rect 4712 9120 4764 9172
rect 5356 9120 5408 9172
rect 6184 9163 6236 9172
rect 6184 9129 6193 9163
rect 6193 9129 6227 9163
rect 6227 9129 6236 9163
rect 6184 9120 6236 9129
rect 9772 9163 9824 9172
rect 9772 9129 9781 9163
rect 9781 9129 9815 9163
rect 9815 9129 9824 9163
rect 9772 9120 9824 9129
rect 1952 9027 2004 9036
rect 1952 8993 1986 9027
rect 1986 8993 2004 9027
rect 1952 8984 2004 8993
rect 2412 8984 2464 9036
rect 3240 8916 3292 8968
rect 3148 8848 3200 8900
rect 5908 9052 5960 9104
rect 7196 9052 7248 9104
rect 5448 8984 5500 9036
rect 5724 8984 5776 9036
rect 8208 8984 8260 9036
rect 8392 9027 8444 9036
rect 8392 8993 8401 9027
rect 8401 8993 8435 9027
rect 8435 8993 8444 9027
rect 8392 8984 8444 8993
rect 8576 9052 8628 9104
rect 9036 9052 9088 9104
rect 11888 9120 11940 9172
rect 12900 9120 12952 9172
rect 13452 9120 13504 9172
rect 14556 9120 14608 9172
rect 15936 9120 15988 9172
rect 16212 9120 16264 9172
rect 16304 9120 16356 9172
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 12716 8984 12768 9036
rect 18236 9052 18288 9104
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 6092 8916 6144 8968
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 8484 8959 8536 8968
rect 8484 8925 8493 8959
rect 8493 8925 8527 8959
rect 8527 8925 8536 8959
rect 8484 8916 8536 8925
rect 8576 8959 8628 8968
rect 8576 8925 8585 8959
rect 8585 8925 8619 8959
rect 8619 8925 8628 8959
rect 8576 8916 8628 8925
rect 8760 8916 8812 8968
rect 11336 8959 11388 8968
rect 8668 8848 8720 8900
rect 2780 8780 2832 8832
rect 3424 8780 3476 8832
rect 5816 8780 5868 8832
rect 8208 8780 8260 8832
rect 8392 8780 8444 8832
rect 9404 8848 9456 8900
rect 9680 8848 9732 8900
rect 11336 8925 11345 8959
rect 11345 8925 11379 8959
rect 11379 8925 11388 8959
rect 11336 8916 11388 8925
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 15476 8959 15528 8968
rect 9036 8780 9088 8832
rect 9772 8780 9824 8832
rect 12164 8780 12216 8832
rect 15476 8925 15485 8959
rect 15485 8925 15519 8959
rect 15519 8925 15528 8959
rect 15476 8916 15528 8925
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 14648 8780 14700 8832
rect 16304 8823 16356 8832
rect 16304 8789 16313 8823
rect 16313 8789 16347 8823
rect 16347 8789 16356 8823
rect 16304 8780 16356 8789
rect 16580 8823 16632 8832
rect 16580 8789 16589 8823
rect 16589 8789 16623 8823
rect 16623 8789 16632 8823
rect 17132 8984 17184 9036
rect 17592 9027 17644 9036
rect 17592 8993 17601 9027
rect 17601 8993 17635 9027
rect 17635 8993 17644 9027
rect 17592 8984 17644 8993
rect 18144 8984 18196 9036
rect 19432 9120 19484 9172
rect 18420 9052 18472 9104
rect 19524 9052 19576 9104
rect 19432 8984 19484 9036
rect 20168 9120 20220 9172
rect 20536 9120 20588 9172
rect 21088 9120 21140 9172
rect 19892 9095 19944 9104
rect 19892 9061 19901 9095
rect 19901 9061 19935 9095
rect 19935 9061 19944 9095
rect 19892 9052 19944 9061
rect 21456 9027 21508 9036
rect 21456 8993 21465 9027
rect 21465 8993 21499 9027
rect 21499 8993 21508 9027
rect 21456 8984 21508 8993
rect 19892 8916 19944 8968
rect 20352 8916 20404 8968
rect 20720 8959 20772 8968
rect 20720 8925 20729 8959
rect 20729 8925 20763 8959
rect 20763 8925 20772 8959
rect 20720 8916 20772 8925
rect 18604 8848 18656 8900
rect 20904 8848 20956 8900
rect 16580 8780 16632 8789
rect 18880 8780 18932 8832
rect 20168 8823 20220 8832
rect 20168 8789 20177 8823
rect 20177 8789 20211 8823
rect 20211 8789 20220 8823
rect 20168 8780 20220 8789
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 2872 8576 2924 8628
rect 1952 8440 2004 8492
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 5448 8619 5500 8628
rect 3240 8551 3292 8560
rect 3240 8517 3249 8551
rect 3249 8517 3283 8551
rect 3283 8517 3292 8551
rect 3240 8508 3292 8517
rect 3516 8440 3568 8492
rect 4252 8508 4304 8560
rect 4988 8508 5040 8560
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 5540 8576 5592 8628
rect 5724 8508 5776 8560
rect 6184 8576 6236 8628
rect 8576 8576 8628 8628
rect 8668 8576 8720 8628
rect 12532 8576 12584 8628
rect 12716 8576 12768 8628
rect 16120 8576 16172 8628
rect 19340 8619 19392 8628
rect 19340 8585 19349 8619
rect 19349 8585 19383 8619
rect 19383 8585 19392 8619
rect 19340 8576 19392 8585
rect 19984 8576 20036 8628
rect 20996 8619 21048 8628
rect 20996 8585 21005 8619
rect 21005 8585 21039 8619
rect 21039 8585 21048 8619
rect 20996 8576 21048 8585
rect 21732 8576 21784 8628
rect 8760 8508 8812 8560
rect 9772 8508 9824 8560
rect 16304 8508 16356 8560
rect 18144 8508 18196 8560
rect 5080 8372 5132 8424
rect 5540 8440 5592 8492
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 11244 8440 11296 8492
rect 16580 8440 16632 8492
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 20352 8440 20404 8492
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 6092 8372 6144 8424
rect 6184 8372 6236 8424
rect 6460 8372 6512 8424
rect 7380 8372 7432 8424
rect 9680 8372 9732 8424
rect 9772 8415 9824 8424
rect 9772 8381 9781 8415
rect 9781 8381 9815 8415
rect 9815 8381 9824 8415
rect 9772 8372 9824 8381
rect 3148 8304 3200 8356
rect 1400 8279 1452 8288
rect 1400 8245 1409 8279
rect 1409 8245 1443 8279
rect 1443 8245 1452 8279
rect 1400 8236 1452 8245
rect 2688 8236 2740 8288
rect 5632 8304 5684 8356
rect 6828 8347 6880 8356
rect 6828 8313 6840 8347
rect 6840 8313 6880 8347
rect 6828 8304 6880 8313
rect 7012 8304 7064 8356
rect 14096 8304 14148 8356
rect 16856 8304 16908 8356
rect 17684 8304 17736 8356
rect 21088 8347 21140 8356
rect 21088 8313 21097 8347
rect 21097 8313 21131 8347
rect 21131 8313 21140 8347
rect 21088 8304 21140 8313
rect 21456 8347 21508 8356
rect 21456 8313 21465 8347
rect 21465 8313 21499 8347
rect 21499 8313 21508 8347
rect 21456 8304 21508 8313
rect 4896 8236 4948 8288
rect 5080 8279 5132 8288
rect 5080 8245 5089 8279
rect 5089 8245 5123 8279
rect 5123 8245 5132 8279
rect 5908 8279 5960 8288
rect 5080 8236 5132 8245
rect 5908 8245 5917 8279
rect 5917 8245 5951 8279
rect 5951 8245 5960 8279
rect 5908 8236 5960 8245
rect 18972 8279 19024 8288
rect 18972 8245 18981 8279
rect 18981 8245 19015 8279
rect 19015 8245 19024 8279
rect 18972 8236 19024 8245
rect 19984 8236 20036 8288
rect 20536 8279 20588 8288
rect 20536 8245 20545 8279
rect 20545 8245 20579 8279
rect 20579 8245 20588 8279
rect 20536 8236 20588 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 1952 8032 2004 8084
rect 1400 7964 1452 8016
rect 15200 8032 15252 8084
rect 18052 8032 18104 8084
rect 18972 8032 19024 8084
rect 19708 8075 19760 8084
rect 19708 8041 19717 8075
rect 19717 8041 19751 8075
rect 19751 8041 19760 8075
rect 19708 8032 19760 8041
rect 20168 8075 20220 8084
rect 20168 8041 20177 8075
rect 20177 8041 20211 8075
rect 20211 8041 20220 8075
rect 20168 8032 20220 8041
rect 20260 8032 20312 8084
rect 21824 8032 21876 8084
rect 3424 7964 3476 8016
rect 1768 7939 1820 7948
rect 1768 7905 1777 7939
rect 1777 7905 1811 7939
rect 1811 7905 1820 7939
rect 1768 7896 1820 7905
rect 3516 7896 3568 7948
rect 3884 7896 3936 7948
rect 5540 7964 5592 8016
rect 6092 7964 6144 8016
rect 8208 7964 8260 8016
rect 8852 7964 8904 8016
rect 20076 8007 20128 8016
rect 20076 7973 20085 8007
rect 20085 7973 20119 8007
rect 20119 7973 20128 8007
rect 20076 7964 20128 7973
rect 20352 7964 20404 8016
rect 20812 7896 20864 7948
rect 21180 7939 21232 7948
rect 21180 7905 21189 7939
rect 21189 7905 21223 7939
rect 21223 7905 21232 7939
rect 21180 7896 21232 7905
rect 21456 7939 21508 7948
rect 21456 7905 21465 7939
rect 21465 7905 21499 7939
rect 21499 7905 21508 7939
rect 21456 7896 21508 7905
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 6184 7871 6236 7880
rect 3056 7692 3108 7744
rect 3148 7692 3200 7744
rect 6184 7837 6193 7871
rect 6193 7837 6227 7871
rect 6227 7837 6236 7871
rect 6184 7828 6236 7837
rect 7380 7828 7432 7880
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 17960 7828 18012 7880
rect 18144 7828 18196 7880
rect 20444 7828 20496 7880
rect 6092 7803 6144 7812
rect 6092 7769 6101 7803
rect 6101 7769 6135 7803
rect 6135 7769 6144 7803
rect 6092 7760 6144 7769
rect 7656 7803 7708 7812
rect 7656 7769 7665 7803
rect 7665 7769 7699 7803
rect 7699 7769 7708 7803
rect 7656 7760 7708 7769
rect 12256 7760 12308 7812
rect 4988 7692 5040 7744
rect 6828 7692 6880 7744
rect 8852 7692 8904 7744
rect 21088 7692 21140 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 1768 7488 1820 7540
rect 14740 7488 14792 7540
rect 16856 7488 16908 7540
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 2872 7463 2924 7472
rect 2872 7429 2881 7463
rect 2881 7429 2915 7463
rect 2915 7429 2924 7463
rect 2872 7420 2924 7429
rect 4896 7463 4948 7472
rect 4896 7429 4905 7463
rect 4905 7429 4939 7463
rect 4939 7429 4948 7463
rect 4896 7420 4948 7429
rect 4988 7420 5040 7472
rect 7380 7463 7432 7472
rect 7380 7429 7389 7463
rect 7389 7429 7423 7463
rect 7423 7429 7432 7463
rect 7380 7420 7432 7429
rect 1492 7352 1544 7404
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 5540 7352 5592 7404
rect 9588 7352 9640 7404
rect 5264 7284 5316 7336
rect 19340 7327 19392 7336
rect 19340 7293 19349 7327
rect 19349 7293 19383 7327
rect 19383 7293 19392 7327
rect 19340 7284 19392 7293
rect 1400 7216 1452 7268
rect 4160 7216 4212 7268
rect 4804 7216 4856 7268
rect 8576 7216 8628 7268
rect 20996 7284 21048 7336
rect 19800 7216 19852 7268
rect 4252 7148 4304 7200
rect 4988 7148 5040 7200
rect 5448 7148 5500 7200
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 20720 7191 20772 7200
rect 20720 7157 20729 7191
rect 20729 7157 20763 7191
rect 20763 7157 20772 7191
rect 20720 7148 20772 7157
rect 21180 7191 21232 7200
rect 21180 7157 21189 7191
rect 21189 7157 21223 7191
rect 21223 7157 21232 7191
rect 21180 7148 21232 7157
rect 21272 7191 21324 7200
rect 21272 7157 21281 7191
rect 21281 7157 21315 7191
rect 21315 7157 21324 7191
rect 21272 7148 21324 7157
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 1400 6944 1452 6996
rect 1676 6944 1728 6996
rect 5724 6944 5776 6996
rect 20996 6987 21048 6996
rect 20996 6953 21005 6987
rect 21005 6953 21039 6987
rect 21039 6953 21048 6987
rect 20996 6944 21048 6953
rect 1492 6851 1544 6860
rect 1492 6817 1501 6851
rect 1501 6817 1535 6851
rect 1535 6817 1544 6851
rect 1492 6808 1544 6817
rect 2964 6851 3016 6860
rect 2964 6817 2982 6851
rect 2982 6817 3016 6851
rect 2964 6808 3016 6817
rect 3424 6808 3476 6860
rect 19340 6808 19392 6860
rect 19616 6851 19668 6860
rect 19616 6817 19625 6851
rect 19625 6817 19659 6851
rect 19659 6817 19668 6851
rect 19616 6808 19668 6817
rect 20720 6808 20772 6860
rect 21456 6851 21508 6860
rect 21456 6817 21465 6851
rect 21465 6817 21499 6851
rect 21499 6817 21508 6851
rect 21456 6808 21508 6817
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 5540 6740 5592 6792
rect 5080 6672 5132 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 3700 6604 3752 6656
rect 11796 6604 11848 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 1584 6400 1636 6452
rect 10508 6400 10560 6452
rect 21088 6332 21140 6384
rect 21180 6264 21232 6316
rect 1492 6171 1544 6180
rect 1492 6137 1501 6171
rect 1501 6137 1535 6171
rect 1535 6137 1544 6171
rect 1492 6128 1544 6137
rect 14648 6128 14700 6180
rect 21456 6171 21508 6180
rect 21456 6137 21465 6171
rect 21465 6137 21499 6171
rect 21499 6137 21508 6171
rect 21456 6128 21508 6137
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 1400 5856 1452 5908
rect 21272 5856 21324 5908
rect 9220 5788 9272 5840
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 20168 5720 20220 5772
rect 21548 5763 21600 5772
rect 21548 5729 21557 5763
rect 21557 5729 21591 5763
rect 21591 5729 21600 5763
rect 21548 5720 21600 5729
rect 21364 5652 21416 5704
rect 20720 5584 20772 5636
rect 20168 5559 20220 5568
rect 20168 5525 20177 5559
rect 20177 5525 20211 5559
rect 20211 5525 20220 5559
rect 20168 5516 20220 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 6276 5244 6328 5296
rect 20904 5244 20956 5296
rect 1492 5151 1544 5160
rect 1492 5117 1501 5151
rect 1501 5117 1535 5151
rect 1535 5117 1544 5151
rect 1492 5108 1544 5117
rect 21456 5151 21508 5160
rect 21456 5117 21465 5151
rect 21465 5117 21499 5151
rect 21499 5117 21508 5151
rect 21456 5108 21508 5117
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 3332 4768 3384 4820
rect 21364 4811 21416 4820
rect 21364 4777 21373 4811
rect 21373 4777 21407 4811
rect 21407 4777 21416 4811
rect 21364 4768 21416 4777
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 1676 4675 1728 4684
rect 1676 4641 1685 4675
rect 1685 4641 1719 4675
rect 1719 4641 1728 4675
rect 1676 4632 1728 4641
rect 21272 4675 21324 4684
rect 21272 4641 21281 4675
rect 21281 4641 21315 4675
rect 21315 4641 21324 4675
rect 21272 4632 21324 4641
rect 21548 4675 21600 4684
rect 21548 4641 21557 4675
rect 21557 4641 21591 4675
rect 21591 4641 21600 4675
rect 21548 4632 21600 4641
rect 20168 4564 20220 4616
rect 6368 4496 6420 4548
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 5356 4224 5408 4276
rect 1400 4063 1452 4072
rect 1400 4029 1409 4063
rect 1409 4029 1443 4063
rect 1443 4029 1452 4063
rect 1400 4020 1452 4029
rect 21548 4063 21600 4072
rect 21548 4029 21557 4063
rect 21557 4029 21591 4063
rect 21591 4029 21600 4063
rect 21548 4020 21600 4029
rect 19892 3884 19944 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 4344 3680 4396 3732
rect 21640 3680 21692 3732
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 21548 3587 21600 3596
rect 21548 3553 21557 3587
rect 21557 3553 21591 3587
rect 21591 3553 21600 3587
rect 21548 3544 21600 3553
rect 21456 3476 21508 3528
rect 1492 3408 1544 3460
rect 1952 3408 2004 3460
rect 19984 3408 20036 3460
rect 20996 3408 21048 3460
rect 1768 3340 1820 3392
rect 20628 3383 20680 3392
rect 20628 3349 20637 3383
rect 20637 3349 20671 3383
rect 20671 3349 20680 3383
rect 20628 3340 20680 3349
rect 21548 3340 21600 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 4252 3136 4304 3188
rect 5172 3136 5224 3188
rect 6736 3136 6788 3188
rect 20444 3136 20496 3188
rect 20996 3136 21048 3188
rect 4988 3068 5040 3120
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 1676 2975 1728 2984
rect 1676 2941 1685 2975
rect 1685 2941 1719 2975
rect 1719 2941 1728 2975
rect 1676 2932 1728 2941
rect 1952 2975 2004 2984
rect 1952 2941 1961 2975
rect 1961 2941 1995 2975
rect 1995 2941 2004 2975
rect 1952 2932 2004 2941
rect 5908 3000 5960 3052
rect 20628 3000 20680 3052
rect 4988 2975 5040 2984
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 11520 2932 11572 2984
rect 20536 2932 20588 2984
rect 20812 2932 20864 2984
rect 21272 2975 21324 2984
rect 21272 2941 21281 2975
rect 21281 2941 21315 2975
rect 21315 2941 21324 2975
rect 21272 2932 21324 2941
rect 21548 2975 21600 2984
rect 21548 2941 21557 2975
rect 21557 2941 21591 2975
rect 21591 2941 21600 2975
rect 21548 2932 21600 2941
rect 2872 2864 2924 2916
rect 5448 2864 5500 2916
rect 15568 2907 15620 2916
rect 15568 2873 15577 2907
rect 15577 2873 15611 2907
rect 15611 2873 15620 2907
rect 15568 2864 15620 2873
rect 20628 2864 20680 2916
rect 2780 2796 2832 2848
rect 18144 2796 18196 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 2044 2592 2096 2644
rect 2688 2592 2740 2644
rect 2964 2635 3016 2644
rect 2964 2601 2973 2635
rect 2973 2601 3007 2635
rect 3007 2601 3016 2635
rect 2964 2592 3016 2601
rect 5172 2592 5224 2644
rect 11520 2635 11572 2644
rect 11520 2601 11529 2635
rect 11529 2601 11563 2635
rect 11563 2601 11572 2635
rect 11520 2592 11572 2601
rect 15568 2592 15620 2644
rect 19432 2592 19484 2644
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 2780 2524 2832 2576
rect 7104 2567 7156 2576
rect 7104 2533 7113 2567
rect 7113 2533 7147 2567
rect 7147 2533 7156 2567
rect 7104 2524 7156 2533
rect 17960 2524 18012 2576
rect 21916 2592 21968 2644
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 2412 2456 2464 2508
rect 3516 2499 3568 2508
rect 3516 2465 3525 2499
rect 3525 2465 3559 2499
rect 3559 2465 3568 2499
rect 3516 2456 3568 2465
rect 11704 2499 11756 2508
rect 11704 2465 11713 2499
rect 11713 2465 11747 2499
rect 11747 2465 11756 2499
rect 11704 2456 11756 2465
rect 16120 2456 16172 2508
rect 20352 2499 20404 2508
rect 20352 2465 20361 2499
rect 20361 2465 20395 2499
rect 20395 2465 20404 2499
rect 20352 2456 20404 2465
rect 20628 2499 20680 2508
rect 20628 2465 20637 2499
rect 20637 2465 20671 2499
rect 20671 2465 20680 2499
rect 20628 2456 20680 2465
rect 20720 2456 20772 2508
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 21456 2499 21508 2508
rect 21456 2465 21465 2499
rect 21465 2465 21499 2499
rect 21499 2465 21508 2499
rect 21456 2456 21508 2465
rect 4988 2388 5040 2440
rect 6920 2363 6972 2372
rect 6920 2329 6929 2363
rect 6929 2329 6963 2363
rect 6963 2329 6972 2363
rect 6920 2320 6972 2329
rect 2872 2252 2924 2304
rect 16120 2252 16172 2304
rect 20444 2252 20496 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 1584 2048 1636 2100
rect 4160 2048 4212 2100
<< metal2 >>
rect 202 22200 258 23000
rect 570 22200 626 23000
rect 1030 22200 1086 23000
rect 1398 22200 1454 23000
rect 1858 22200 1914 23000
rect 2318 22200 2374 23000
rect 2686 22200 2742 23000
rect 3146 22200 3202 23000
rect 3330 22264 3386 22273
rect 216 19854 244 22200
rect 584 20330 612 22200
rect 1044 20398 1072 22200
rect 1412 20806 1440 22200
rect 1872 20874 1900 22200
rect 1860 20868 1912 20874
rect 1860 20810 1912 20816
rect 1400 20800 1452 20806
rect 1400 20742 1452 20748
rect 1858 20768 1914 20777
rect 1858 20703 1914 20712
rect 1492 20528 1544 20534
rect 1492 20470 1544 20476
rect 1032 20392 1084 20398
rect 1032 20334 1084 20340
rect 1504 20330 1532 20470
rect 572 20324 624 20330
rect 572 20266 624 20272
rect 1492 20324 1544 20330
rect 1492 20266 1544 20272
rect 1872 20058 1900 20703
rect 2134 20360 2190 20369
rect 2134 20295 2136 20304
rect 2188 20295 2190 20304
rect 2136 20266 2188 20272
rect 2228 20256 2280 20262
rect 2228 20198 2280 20204
rect 1860 20052 1912 20058
rect 1860 19994 1912 20000
rect 2044 19984 2096 19990
rect 2044 19926 2096 19932
rect 1584 19916 1636 19922
rect 1584 19858 1636 19864
rect 1952 19916 2004 19922
rect 1952 19858 2004 19864
rect 204 19848 256 19854
rect 204 19790 256 19796
rect 1398 19816 1454 19825
rect 1398 19751 1400 19760
rect 1452 19751 1454 19760
rect 1400 19722 1452 19728
rect 1596 19446 1624 19858
rect 1768 19780 1820 19786
rect 1768 19722 1820 19728
rect 1584 19440 1636 19446
rect 1398 19408 1454 19417
rect 1584 19382 1636 19388
rect 1398 19343 1454 19352
rect 1412 19310 1440 19343
rect 1780 19310 1808 19722
rect 1964 19514 1992 19858
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 2056 19360 2084 19926
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2148 19378 2176 19858
rect 2240 19394 2268 20198
rect 2332 20074 2360 22200
rect 2700 20942 2728 22200
rect 2962 21720 3018 21729
rect 2962 21655 3018 21664
rect 2778 21312 2834 21321
rect 2778 21247 2834 21256
rect 2688 20936 2740 20942
rect 2688 20878 2740 20884
rect 2792 20602 2820 21247
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2594 20496 2650 20505
rect 2594 20431 2596 20440
rect 2648 20431 2650 20440
rect 2778 20496 2834 20505
rect 2778 20431 2780 20440
rect 2596 20402 2648 20408
rect 2832 20431 2834 20440
rect 2780 20402 2832 20408
rect 2502 20360 2558 20369
rect 2502 20295 2504 20304
rect 2556 20295 2558 20304
rect 2504 20266 2556 20272
rect 2332 20046 2544 20074
rect 2516 19990 2544 20046
rect 2504 19984 2556 19990
rect 2504 19926 2556 19932
rect 2688 19848 2740 19854
rect 2594 19816 2650 19825
rect 2688 19790 2740 19796
rect 2594 19751 2596 19760
rect 2648 19751 2650 19760
rect 2596 19722 2648 19728
rect 2700 19446 2728 19790
rect 2884 19768 2912 20742
rect 2976 20602 3004 21655
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 3056 20324 3108 20330
rect 3056 20266 3108 20272
rect 2964 19780 3016 19786
rect 2884 19740 2964 19768
rect 2964 19722 3016 19728
rect 2780 19712 2832 19718
rect 2976 19689 3004 19722
rect 2780 19654 2832 19660
rect 2962 19680 3018 19689
rect 2688 19440 2740 19446
rect 1872 19332 2084 19360
rect 2136 19372 2188 19378
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1768 19304 1820 19310
rect 1768 19246 1820 19252
rect 1398 18864 1454 18873
rect 1398 18799 1400 18808
rect 1452 18799 1454 18808
rect 1584 18828 1636 18834
rect 1400 18770 1452 18776
rect 1584 18770 1636 18776
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1490 18456 1546 18465
rect 1596 18426 1624 18770
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1490 18391 1492 18400
rect 1544 18391 1546 18400
rect 1584 18420 1636 18426
rect 1492 18362 1544 18368
rect 1584 18362 1636 18368
rect 1584 18148 1636 18154
rect 1584 18090 1636 18096
rect 1492 17536 1544 17542
rect 1490 17504 1492 17513
rect 1544 17504 1546 17513
rect 1490 17439 1546 17448
rect 1596 17270 1624 18090
rect 1584 17264 1636 17270
rect 1584 17206 1636 17212
rect 1398 17096 1454 17105
rect 1398 17031 1400 17040
rect 1452 17031 1454 17040
rect 1584 17060 1636 17066
rect 1400 17002 1452 17008
rect 1584 17002 1636 17008
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1412 16561 1440 16594
rect 1398 16552 1454 16561
rect 1398 16487 1454 16496
rect 1596 16250 1624 17002
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1398 16144 1454 16153
rect 1398 16079 1400 16088
rect 1452 16079 1454 16088
rect 1400 16050 1452 16056
rect 1584 15972 1636 15978
rect 1584 15914 1636 15920
rect 1596 15706 1624 15914
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1398 15600 1454 15609
rect 1398 15535 1400 15544
rect 1452 15535 1454 15544
rect 1400 15506 1452 15512
rect 1490 15192 1546 15201
rect 1490 15127 1492 15136
rect 1544 15127 1546 15136
rect 1492 15098 1544 15104
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1492 14272 1544 14278
rect 1490 14240 1492 14249
rect 1544 14240 1546 14249
rect 1490 14175 1546 14184
rect 1400 13864 1452 13870
rect 1320 13812 1400 13818
rect 1320 13806 1452 13812
rect 1320 13790 1440 13806
rect 1320 13705 1348 13790
rect 1306 13696 1362 13705
rect 1306 13631 1362 13640
rect 1320 12889 1348 13631
rect 1492 13456 1544 13462
rect 1492 13398 1544 13404
rect 1398 13288 1454 13297
rect 1398 13223 1454 13232
rect 1412 12918 1440 13223
rect 1400 12912 1452 12918
rect 1306 12880 1362 12889
rect 1400 12854 1452 12860
rect 1306 12815 1362 12824
rect 1412 12782 1440 12854
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1504 12209 1532 13398
rect 1490 12200 1546 12209
rect 1490 12135 1546 12144
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 10538 1440 11494
rect 1504 11218 1532 12038
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1504 10985 1532 11154
rect 1490 10976 1546 10985
rect 1490 10911 1546 10920
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1400 10532 1452 10538
rect 1400 10474 1452 10480
rect 1412 10441 1440 10474
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 1504 10130 1532 10610
rect 1596 10266 1624 14418
rect 1688 12434 1716 18702
rect 1780 18290 1808 18770
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1872 18170 1900 19332
rect 2240 19366 2636 19394
rect 2688 19382 2740 19388
rect 2136 19314 2188 19320
rect 2412 19304 2464 19310
rect 1950 19272 2006 19281
rect 2412 19246 2464 19252
rect 1950 19207 2006 19216
rect 2044 19236 2096 19242
rect 1964 19174 1992 19207
rect 2044 19178 2096 19184
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 2056 18358 2084 19178
rect 2136 18828 2188 18834
rect 2136 18770 2188 18776
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2044 18352 2096 18358
rect 2044 18294 2096 18300
rect 1780 18142 1900 18170
rect 1952 18148 2004 18154
rect 1780 13954 1808 18142
rect 1952 18090 2004 18096
rect 1860 18080 1912 18086
rect 1858 18048 1860 18057
rect 1912 18048 1914 18057
rect 1858 17983 1914 17992
rect 1860 17740 1912 17746
rect 1860 17682 1912 17688
rect 1872 15910 1900 17682
rect 1964 17338 1992 18090
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1860 15904 1912 15910
rect 1860 15846 1912 15852
rect 1964 15706 1992 16594
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 2056 16182 2084 16390
rect 2044 16176 2096 16182
rect 2044 16118 2096 16124
rect 2056 16046 2084 16118
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2148 15586 2176 18770
rect 2226 18728 2282 18737
rect 2226 18663 2228 18672
rect 2280 18663 2282 18672
rect 2228 18634 2280 18640
rect 2332 16130 2360 18770
rect 2424 18630 2452 19246
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2516 18873 2544 18906
rect 2502 18864 2558 18873
rect 2502 18799 2558 18808
rect 2412 18624 2464 18630
rect 2412 18566 2464 18572
rect 2608 18306 2636 19366
rect 2688 19304 2740 19310
rect 2688 19246 2740 19252
rect 2700 18766 2728 19246
rect 2792 18816 2820 19654
rect 2962 19615 3018 19624
rect 3068 19514 3096 20266
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2870 19000 2926 19009
rect 2870 18935 2872 18944
rect 2924 18935 2926 18944
rect 2872 18906 2924 18912
rect 2792 18788 2912 18816
rect 2688 18760 2740 18766
rect 2688 18702 2740 18708
rect 2608 18278 2728 18306
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 2608 17882 2636 18158
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2700 16658 2728 18278
rect 2884 17354 2912 18788
rect 2976 18698 3004 19110
rect 2964 18692 3016 18698
rect 2964 18634 3016 18640
rect 2884 17326 3004 17354
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 2884 16250 2912 17138
rect 2976 17066 3004 17326
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2976 16794 3004 17002
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 1964 15558 2176 15586
rect 2240 16102 2360 16130
rect 1858 14648 1914 14657
rect 1858 14583 1860 14592
rect 1912 14583 1914 14592
rect 1860 14554 1912 14560
rect 1780 13926 1900 13954
rect 1768 13864 1820 13870
rect 1766 13832 1768 13841
rect 1820 13832 1822 13841
rect 1872 13802 1900 13926
rect 1766 13767 1822 13776
rect 1860 13796 1912 13802
rect 1860 13738 1912 13744
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1780 13394 1808 13670
rect 1964 13512 1992 15558
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 2148 14618 2176 15438
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 2148 14074 2176 14418
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1872 13484 1992 13512
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1780 12594 1808 13330
rect 1872 12730 1900 13484
rect 1950 12880 2006 12889
rect 1950 12815 1952 12824
rect 2004 12815 2006 12824
rect 1952 12786 2004 12792
rect 1872 12702 1992 12730
rect 1780 12566 1900 12594
rect 1688 12406 1808 12434
rect 1676 12368 1728 12374
rect 1676 12310 1728 12316
rect 1688 11354 1716 12310
rect 1780 11506 1808 12406
rect 1872 12345 1900 12566
rect 1858 12336 1914 12345
rect 1858 12271 1914 12280
rect 1780 11478 1900 11506
rect 1766 11384 1822 11393
rect 1676 11348 1728 11354
rect 1766 11319 1822 11328
rect 1676 11290 1728 11296
rect 1780 11218 1808 11319
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1674 10568 1730 10577
rect 1674 10503 1676 10512
rect 1728 10503 1730 10512
rect 1676 10474 1728 10480
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1504 10033 1532 10066
rect 1490 10024 1546 10033
rect 1872 10010 1900 11478
rect 1964 11354 1992 12702
rect 2056 11540 2084 13806
rect 2136 13796 2188 13802
rect 2136 13738 2188 13744
rect 2148 12986 2176 13738
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 2148 12442 2176 12786
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2056 11512 2176 11540
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1490 9959 1546 9968
rect 1688 9982 1900 10010
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1504 9081 1532 9386
rect 1596 9178 1624 9454
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1490 9072 1546 9081
rect 1490 9007 1546 9016
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 8129 1440 8230
rect 1398 8120 1454 8129
rect 1398 8055 1454 8064
rect 1412 8022 1440 8055
rect 1400 8016 1452 8022
rect 1400 7958 1452 7964
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1400 7268 1452 7274
rect 1400 7210 1452 7216
rect 1412 7177 1440 7210
rect 1398 7168 1454 7177
rect 1398 7103 1454 7112
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1412 5914 1440 6938
rect 1504 6866 1532 7346
rect 1688 7002 1716 9982
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1872 9450 1900 9862
rect 1964 9722 1992 10066
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 2056 9489 2084 10066
rect 2148 9654 2176 11512
rect 2240 10266 2268 16102
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2332 15706 2360 15982
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2884 15026 2912 16186
rect 3068 15858 3096 19246
rect 3160 18970 3188 22200
rect 3330 22199 3386 22208
rect 3606 22200 3662 23000
rect 3882 22672 3938 22681
rect 3882 22607 3938 22616
rect 3344 20602 3372 22199
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 3424 20868 3476 20874
rect 3424 20810 3476 20816
rect 3332 20596 3384 20602
rect 3332 20538 3384 20544
rect 3238 20360 3294 20369
rect 3238 20295 3294 20304
rect 3332 20324 3384 20330
rect 3252 19514 3280 20295
rect 3332 20266 3384 20272
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3160 18426 3188 18566
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3146 18320 3202 18329
rect 3146 18255 3202 18264
rect 3160 18222 3188 18255
rect 3148 18216 3200 18222
rect 3148 18158 3200 18164
rect 3252 18086 3280 19314
rect 3344 18902 3372 20266
rect 3436 19961 3464 20810
rect 3422 19952 3478 19961
rect 3528 19922 3556 20878
rect 3620 20262 3648 22200
rect 3792 20596 3844 20602
rect 3792 20538 3844 20544
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3422 19887 3424 19896
rect 3476 19887 3478 19896
rect 3516 19916 3568 19922
rect 3424 19858 3476 19864
rect 3516 19858 3568 19864
rect 3424 19780 3476 19786
rect 3424 19722 3476 19728
rect 3436 19514 3464 19722
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3712 19378 3740 20266
rect 3804 19786 3832 20538
rect 3896 20534 3924 22607
rect 3974 22200 4030 23000
rect 4434 22200 4490 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6090 22200 6146 23000
rect 6550 22200 6606 23000
rect 7010 22200 7066 23000
rect 7378 22200 7434 23000
rect 7838 22200 7894 23000
rect 8206 22200 8262 23000
rect 8666 22200 8722 23000
rect 9126 22200 9182 23000
rect 9494 22200 9550 23000
rect 9954 22200 10010 23000
rect 10414 22200 10470 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12070 22200 12126 23000
rect 12530 22200 12586 23000
rect 12898 22200 12954 23000
rect 13358 22200 13414 23000
rect 13818 22200 13874 23000
rect 14186 22200 14242 23000
rect 14646 22200 14702 23000
rect 15106 22200 15162 23000
rect 15474 22200 15530 23000
rect 15934 22200 15990 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17590 22200 17646 23000
rect 18050 22200 18106 23000
rect 18510 22200 18566 23000
rect 18878 22200 18934 23000
rect 18970 22672 19026 22681
rect 18970 22607 19026 22616
rect 3884 20528 3936 20534
rect 3884 20470 3936 20476
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 3792 19780 3844 19786
rect 3792 19722 3844 19728
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3608 19304 3660 19310
rect 3608 19246 3660 19252
rect 3332 18896 3384 18902
rect 3332 18838 3384 18844
rect 3528 18766 3556 19246
rect 3620 18970 3648 19246
rect 3700 19168 3752 19174
rect 3700 19110 3752 19116
rect 3608 18964 3660 18970
rect 3608 18906 3660 18912
rect 3712 18902 3740 19110
rect 3700 18896 3752 18902
rect 3700 18838 3752 18844
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3344 18630 3372 18702
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3344 16794 3372 16934
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3068 15830 3188 15858
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2596 14476 2648 14482
rect 2596 14418 2648 14424
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2332 12442 2360 13262
rect 2608 12986 2636 14418
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2700 13705 2728 14010
rect 2686 13696 2742 13705
rect 2686 13631 2742 13640
rect 2964 13388 3016 13394
rect 2964 13330 3016 13336
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2424 11626 2452 12786
rect 2792 12646 2820 12922
rect 2976 12889 3004 13330
rect 2962 12880 3018 12889
rect 2962 12815 3018 12824
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2884 12306 2912 12378
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 2700 11898 2728 12242
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2884 11694 2912 12242
rect 2872 11688 2924 11694
rect 2792 11648 2872 11676
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2424 11082 2452 11562
rect 2412 11076 2464 11082
rect 2412 11018 2464 11024
rect 2424 10674 2452 11018
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2332 9654 2360 10406
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2042 9480 2098 9489
rect 1860 9444 1912 9450
rect 2042 9415 2098 9424
rect 1860 9386 1912 9392
rect 1872 8673 1900 9386
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1858 8664 1914 8673
rect 1858 8599 1914 8608
rect 1964 8498 1992 8978
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1964 8090 1992 8434
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1780 7721 1808 7890
rect 1766 7712 1822 7721
rect 1766 7647 1822 7656
rect 1780 7546 1808 7647
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1504 6769 1532 6802
rect 1490 6760 1546 6769
rect 1490 6695 1546 6704
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 6458 1624 6598
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1490 6216 1546 6225
rect 1490 6151 1492 6160
rect 1544 6151 1546 6160
rect 1492 6122 1544 6128
rect 1400 5908 1452 5914
rect 1400 5850 1452 5856
rect 1398 5808 1454 5817
rect 1398 5743 1400 5752
rect 1452 5743 1454 5752
rect 1400 5714 1452 5720
rect 1490 5264 1546 5273
rect 1490 5199 1546 5208
rect 1504 5166 1532 5199
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1674 4856 1730 4865
rect 1674 4791 1730 4800
rect 1688 4690 1716 4791
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1412 4457 1440 4626
rect 1398 4448 1454 4457
rect 1398 4383 1454 4392
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 1412 3913 1440 4014
rect 1398 3904 1454 3913
rect 1398 3839 1454 3848
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1412 3505 1440 3538
rect 1398 3496 1454 3505
rect 1398 3431 1454 3440
rect 1492 3460 1544 3466
rect 1492 3402 1544 3408
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1400 2984 1452 2990
rect 1398 2952 1400 2961
rect 1452 2952 1454 2961
rect 1398 2887 1454 2896
rect 1398 2544 1454 2553
rect 1504 2530 1532 3402
rect 1768 3392 1820 3398
rect 1688 3340 1768 3346
rect 1688 3334 1820 3340
rect 1688 3318 1808 3334
rect 1688 2990 1716 3318
rect 1964 2990 1992 3402
rect 1676 2984 1728 2990
rect 1676 2926 1728 2932
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 1454 2502 1532 2530
rect 1398 2479 1400 2488
rect 1452 2479 1454 2488
rect 1400 2450 1452 2456
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1596 2106 1624 2246
rect 1584 2100 1636 2106
rect 1584 2042 1636 2048
rect 1688 1057 1716 2926
rect 1964 1601 1992 2926
rect 2044 2644 2096 2650
rect 2332 2632 2360 9590
rect 2792 9586 2820 11648
rect 2872 11630 2924 11636
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2884 10674 2912 11154
rect 2976 11082 3004 12718
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 3068 11830 3096 12650
rect 3056 11824 3108 11830
rect 3056 11766 3108 11772
rect 3160 11370 3188 15830
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3252 11694 3280 12582
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3068 11342 3188 11370
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2608 9178 2636 9454
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2424 8634 2452 8978
rect 2792 8838 2820 9522
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2884 8945 2912 9318
rect 2870 8936 2926 8945
rect 2870 8871 2926 8880
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2700 2650 2728 8230
rect 2792 8129 2820 8434
rect 2778 8120 2834 8129
rect 2778 8055 2834 8064
rect 2884 7478 2912 8570
rect 3068 7750 3096 11342
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3344 11234 3372 14758
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3436 12442 3464 13806
rect 3528 12986 3556 17546
rect 3804 17134 3832 19722
rect 3896 18970 3924 20334
rect 3988 19310 4016 22200
rect 4448 20890 4476 22200
rect 4356 20862 4476 20890
rect 4356 20534 4384 20862
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4816 20534 4844 22200
rect 5276 20534 5304 22200
rect 4344 20528 4396 20534
rect 4344 20470 4396 20476
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5736 20398 5764 22200
rect 6104 20398 6132 22200
rect 6564 20398 6592 22200
rect 6736 20528 6788 20534
rect 6736 20470 6788 20476
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 6092 20392 6144 20398
rect 6092 20334 6144 20340
rect 6552 20392 6604 20398
rect 6552 20334 6604 20340
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 4080 20058 4108 20266
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4172 19961 4200 19994
rect 4158 19952 4214 19961
rect 4264 19922 4292 20198
rect 4158 19887 4214 19896
rect 4252 19916 4304 19922
rect 4252 19858 4304 19864
rect 4068 19780 4120 19786
rect 4068 19722 4120 19728
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 4080 19446 4108 19722
rect 4264 19689 4292 19722
rect 4908 19718 4936 20266
rect 4896 19712 4948 19718
rect 4250 19680 4306 19689
rect 4896 19654 4948 19660
rect 4250 19615 4306 19624
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4068 19440 4120 19446
rect 4068 19382 4120 19388
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 19174 4016 19246
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 4080 17649 4108 18566
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4066 17640 4122 17649
rect 4066 17575 4068 17584
rect 4120 17575 4122 17584
rect 4068 17546 4120 17552
rect 3884 17536 3936 17542
rect 4080 17515 4108 17546
rect 3884 17478 3936 17484
rect 3896 17338 3924 17478
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3896 16590 3924 17070
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3712 15978 3740 16458
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3620 13938 3648 14554
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3620 12782 3648 13126
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3160 10742 3188 11222
rect 3344 11206 3464 11234
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3344 10810 3372 11086
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3148 10736 3200 10742
rect 3148 10678 3200 10684
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3160 8906 3188 9454
rect 3240 8968 3292 8974
rect 3436 8922 3464 11206
rect 3528 11150 3556 11698
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3240 8910 3292 8916
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3252 8566 3280 8910
rect 3344 8894 3464 8922
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3160 7750 3188 8298
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2096 2604 2360 2632
rect 2688 2644 2740 2650
rect 2044 2586 2096 2592
rect 2688 2586 2740 2592
rect 2792 2582 2820 2790
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 2424 2394 2452 2450
rect 2332 2366 2452 2394
rect 1950 1592 2006 1601
rect 1950 1527 2006 1536
rect 1674 1048 1730 1057
rect 1674 983 1730 992
rect 2332 800 2360 2366
rect 2318 0 2374 800
rect 2792 649 2820 2518
rect 2884 2310 2912 2858
rect 2976 2650 3004 6802
rect 3344 4826 3372 8894
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3436 8022 3464 8774
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3424 8016 3476 8022
rect 3424 7958 3476 7964
rect 3436 7886 3464 7958
rect 3528 7954 3556 8434
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3436 6866 3464 7822
rect 3528 7410 3556 7890
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3712 6662 3740 15914
rect 3804 12986 3832 16118
rect 3896 16046 3924 16526
rect 3988 16250 4016 16594
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 4172 16046 4200 16934
rect 4356 16114 4384 17002
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4160 16040 4212 16046
rect 4160 15982 4212 15988
rect 3976 15972 4028 15978
rect 3976 15914 4028 15920
rect 3988 15706 4016 15914
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 4080 14958 4108 15982
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3896 14278 3924 14826
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3896 14006 3924 14214
rect 4356 14074 4384 15642
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4816 14074 4844 15438
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4632 13530 4660 13806
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 13530 4752 13670
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 12442 4752 12582
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4344 12300 4396 12306
rect 3988 12238 4016 12269
rect 4344 12242 4396 12248
rect 3976 12232 4028 12238
rect 3974 12200 3976 12209
rect 4028 12200 4030 12209
rect 3974 12135 4030 12144
rect 3988 11762 4016 12135
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 4356 11354 4384 12242
rect 4712 12232 4764 12238
rect 4710 12200 4712 12209
rect 4764 12200 4766 12209
rect 4710 12135 4766 12144
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4436 11620 4488 11626
rect 4436 11562 4488 11568
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4172 10656 4200 10950
rect 4264 10810 4292 11086
rect 4356 10810 4384 11154
rect 4448 11150 4476 11562
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4172 10628 4292 10656
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3804 10266 3832 10406
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3884 7948 3936 7954
rect 3884 7890 3936 7896
rect 3896 7410 3924 7890
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 4172 7274 4200 10474
rect 4264 9450 4292 10628
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4724 10418 4752 10542
rect 4816 10538 4844 13806
rect 4908 12073 4936 19654
rect 4988 18148 5040 18154
rect 4988 18090 5040 18096
rect 5000 15858 5028 18090
rect 5092 15994 5120 20334
rect 6104 20058 6132 20334
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6092 20052 6144 20058
rect 6092 19994 6144 20000
rect 6288 19718 6316 20198
rect 6276 19712 6328 19718
rect 6276 19654 6328 19660
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5356 18828 5408 18834
rect 5356 18770 5408 18776
rect 5368 18426 5396 18770
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 5184 17338 5212 18158
rect 5356 17808 5408 17814
rect 5460 17796 5488 19450
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 5908 19236 5960 19242
rect 5908 19178 5960 19184
rect 5920 18902 5948 19178
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 6104 18970 6132 19110
rect 6472 18970 6500 19246
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 5632 18352 5684 18358
rect 5632 18294 5684 18300
rect 5540 17808 5592 17814
rect 5460 17768 5540 17796
rect 5356 17750 5408 17756
rect 5540 17750 5592 17756
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5368 17270 5396 17750
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5276 16114 5304 16390
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5368 16046 5396 16390
rect 5552 16182 5580 16934
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 5356 16040 5408 16046
rect 5092 15966 5304 15994
rect 5356 15982 5408 15988
rect 5000 15830 5120 15858
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 5000 13802 5028 14418
rect 4988 13796 5040 13802
rect 4988 13738 5040 13744
rect 5092 13394 5120 15830
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5080 13388 5132 13394
rect 5080 13330 5132 13336
rect 4894 12064 4950 12073
rect 4894 11999 4950 12008
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4908 10470 4936 11834
rect 5000 11762 5028 13330
rect 5184 13326 5212 13738
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 11234 5028 11698
rect 5092 11354 5120 12582
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 5184 11830 5212 12242
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 5276 11608 5304 15966
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5368 15162 5396 15846
rect 5460 15706 5488 15846
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5644 15586 5672 18294
rect 5736 16794 5764 18838
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 5816 17264 5868 17270
rect 5868 17212 6040 17218
rect 5816 17206 6040 17212
rect 5828 17202 6040 17206
rect 5828 17196 6052 17202
rect 5828 17190 6000 17196
rect 6000 17138 6052 17144
rect 5816 17060 5868 17066
rect 5816 17002 5868 17008
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5828 16250 5856 17002
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5644 15558 5764 15586
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5552 15162 5580 15438
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5552 14550 5580 15098
rect 5644 14822 5672 15438
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5368 11830 5396 12786
rect 5736 12753 5764 15558
rect 6012 15502 6040 16526
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 5920 14958 5948 15302
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5920 14278 5948 14894
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5722 12744 5778 12753
rect 5448 12708 5500 12714
rect 5722 12679 5778 12688
rect 5448 12650 5500 12656
rect 5460 11898 5488 12650
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5184 11580 5304 11608
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5000 11206 5120 11234
rect 4896 10464 4948 10470
rect 4724 10390 4844 10418
rect 4896 10406 4948 10412
rect 4816 10130 4844 10390
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 4356 9353 4384 9658
rect 4526 9616 4582 9625
rect 4526 9551 4528 9560
rect 4580 9551 4582 9560
rect 4528 9522 4580 9528
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4342 9344 4398 9353
rect 4342 9279 4398 9288
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2778 640 2834 649
rect 2778 575 2834 584
rect 2884 241 2912 2246
rect 3528 2009 3556 2450
rect 4172 2106 4200 7210
rect 4264 7206 4292 8502
rect 4356 7886 4384 9279
rect 4724 9178 4752 9386
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4264 3194 4292 7142
rect 4356 3738 4384 7822
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4816 7274 4844 10066
rect 4908 8537 4936 10406
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9722 5028 9998
rect 4988 9716 5040 9722
rect 4988 9658 5040 9664
rect 5000 8566 5028 9658
rect 4988 8560 5040 8566
rect 4894 8528 4950 8537
rect 4988 8502 5040 8508
rect 4894 8463 4950 8472
rect 5092 8430 5120 11206
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 4908 7478 4936 8230
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 5000 7478 5028 7686
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 5000 3126 5028 7142
rect 5092 6730 5120 8230
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 5184 3194 5212 11580
rect 5262 11520 5318 11529
rect 5262 11455 5318 11464
rect 5276 7449 5304 11455
rect 5368 11082 5396 11766
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11286 5488 11494
rect 5736 11354 5764 12679
rect 5828 11558 5856 13330
rect 6012 11898 6040 14758
rect 6104 13870 6132 17478
rect 6196 17134 6224 17682
rect 6472 17270 6500 17818
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6460 17264 6512 17270
rect 6460 17206 6512 17212
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6196 16590 6224 17070
rect 6564 16726 6592 17478
rect 6552 16720 6604 16726
rect 6552 16662 6604 16668
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6196 15366 6224 16526
rect 6288 15910 6316 16594
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6288 14056 6316 15846
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6196 14028 6316 14056
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5460 10674 5488 11086
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 10266 5488 10610
rect 5552 10606 5580 11018
rect 5736 10810 5764 11290
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5540 10600 5592 10606
rect 5592 10548 5764 10554
rect 5540 10542 5764 10548
rect 5552 10526 5764 10542
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5552 10198 5580 10406
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5644 9654 5672 10406
rect 5736 10062 5764 10526
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5632 9648 5684 9654
rect 5736 9625 5764 9998
rect 5632 9590 5684 9596
rect 5722 9616 5778 9625
rect 5722 9551 5778 9560
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5262 7440 5318 7449
rect 5262 7375 5318 7384
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5000 2446 5028 2926
rect 5276 2774 5304 7278
rect 5368 6798 5396 9114
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5460 8634 5488 8978
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5446 8528 5502 8537
rect 5552 8498 5580 8570
rect 5446 8463 5502 8472
rect 5540 8492 5592 8498
rect 5460 7206 5488 8463
rect 5540 8434 5592 8440
rect 5552 8022 5580 8434
rect 5644 8362 5672 8910
rect 5736 8566 5764 8978
rect 5828 8922 5856 11494
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5920 9518 5948 11154
rect 6196 9586 6224 14028
rect 6472 14006 6500 14758
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6564 13546 6592 14486
rect 6656 13716 6684 20198
rect 6748 14550 6776 20470
rect 7024 20398 7052 22200
rect 7392 20398 7420 22200
rect 7472 20528 7524 20534
rect 7472 20470 7524 20476
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6932 19904 6960 20198
rect 7024 20058 7052 20334
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 6932 19876 7144 19904
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 6932 17814 6960 19722
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6932 17338 6960 17614
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6828 17264 6880 17270
rect 6880 17212 6960 17218
rect 6828 17206 6960 17212
rect 6840 17190 6960 17206
rect 6932 15162 6960 17190
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6840 14482 6868 14962
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6840 13870 6868 14418
rect 6932 14346 6960 14418
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6656 13688 6868 13716
rect 6564 13518 6776 13546
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6460 12232 6512 12238
rect 6458 12200 6460 12209
rect 6512 12200 6514 12209
rect 6458 12135 6514 12144
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5920 9110 5948 9454
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 6092 8968 6144 8974
rect 5828 8894 5948 8922
rect 6092 8910 6144 8916
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5828 8498 5856 8774
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5920 8294 5948 8894
rect 6104 8430 6132 8910
rect 6196 8634 6224 9114
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5552 7410 5580 7958
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5446 7032 5502 7041
rect 5446 6967 5502 6976
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 4282 5396 6734
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5460 2922 5488 6967
rect 5552 6798 5580 7346
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5736 7002 5764 7142
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5920 3058 5948 8230
rect 6104 8022 6132 8366
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6104 7818 6132 7958
rect 6196 7886 6224 8366
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 6288 5302 6316 11834
rect 6472 10470 6500 12135
rect 6564 11898 6592 12582
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6564 11218 6592 11698
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6656 11150 6684 11766
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6380 4554 6408 9522
rect 6472 8430 6500 10406
rect 6656 10198 6684 10950
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6748 9654 6776 13518
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6840 8514 6868 13688
rect 6932 13326 6960 14282
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 6932 12850 6960 13262
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11354 6960 11494
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7024 10810 7052 18770
rect 7116 17921 7144 19876
rect 7102 17912 7158 17921
rect 7102 17847 7158 17856
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 7116 16250 7144 17682
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7208 14958 7236 20198
rect 7484 18306 7512 20470
rect 7852 20398 7880 22200
rect 8220 20398 8248 22200
rect 8680 20398 8708 22200
rect 9140 20398 9168 22200
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 8220 20058 8248 20334
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8680 19990 8708 20334
rect 8760 20256 8812 20262
rect 9036 20256 9088 20262
rect 8760 20198 8812 20204
rect 8956 20216 9036 20244
rect 8668 19984 8720 19990
rect 8668 19926 8720 19932
rect 8772 19922 8800 20198
rect 8852 19984 8904 19990
rect 8852 19926 8904 19932
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8760 19916 8812 19922
rect 8760 19858 8812 19864
rect 8116 19440 8168 19446
rect 8116 19382 8168 19388
rect 7748 19372 7800 19378
rect 7748 19314 7800 19320
rect 8128 19334 8156 19382
rect 7654 19000 7710 19009
rect 7654 18935 7710 18944
rect 7668 18426 7696 18935
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7392 18278 7512 18306
rect 7564 18284 7616 18290
rect 7288 18216 7340 18222
rect 7286 18184 7288 18193
rect 7340 18184 7342 18193
rect 7286 18119 7342 18128
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7300 17882 7328 18022
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7300 15706 7328 15846
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7116 14006 7144 14214
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7300 11370 7328 15370
rect 7392 11762 7420 18278
rect 7564 18226 7616 18232
rect 7472 18216 7524 18222
rect 7472 18158 7524 18164
rect 7484 17882 7512 18158
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7470 17776 7526 17785
rect 7470 17711 7526 17720
rect 7484 14550 7512 17711
rect 7576 17066 7604 18226
rect 7656 18148 7708 18154
rect 7656 18090 7708 18096
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7576 16522 7604 17002
rect 7668 16522 7696 18090
rect 7760 17882 7788 19314
rect 8128 19306 8524 19334
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8312 18426 8340 18770
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8404 18426 8432 18634
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 7930 18320 7986 18329
rect 7930 18255 7932 18264
rect 7984 18255 7986 18264
rect 7932 18226 7984 18232
rect 8390 18184 8446 18193
rect 8390 18119 8446 18128
rect 8404 18086 8432 18119
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7760 16640 7788 17682
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7840 16652 7892 16658
rect 7760 16612 7840 16640
rect 7840 16594 7892 16600
rect 8220 16590 8248 17546
rect 8312 17542 8340 18022
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 7656 16516 7708 16522
rect 7656 16458 7708 16464
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 7576 16114 7604 16458
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7852 15994 7880 16458
rect 8128 16454 8156 16526
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8220 16114 8248 16526
rect 8312 16130 8340 17070
rect 8404 16522 8432 18022
rect 8496 17320 8524 19306
rect 8588 18970 8616 19858
rect 8864 19718 8892 19926
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8852 18896 8904 18902
rect 8852 18838 8904 18844
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8680 18222 8708 18566
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8864 18154 8892 18838
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8576 17332 8628 17338
rect 8496 17292 8576 17320
rect 8392 16516 8444 16522
rect 8392 16458 8444 16464
rect 8496 16454 8524 17292
rect 8576 17274 8628 17280
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8852 16176 8904 16182
rect 8208 16108 8260 16114
rect 8312 16102 8616 16130
rect 8852 16118 8904 16124
rect 8208 16050 8260 16056
rect 7576 15966 7880 15994
rect 8220 15994 8248 16050
rect 8392 16040 8444 16046
rect 8220 15966 8340 15994
rect 8392 15982 8444 15988
rect 7472 14544 7524 14550
rect 7472 14486 7524 14492
rect 7576 13530 7604 15966
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8220 15638 8248 15846
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8220 15314 8248 15438
rect 8312 15434 8340 15966
rect 8404 15706 8432 15982
rect 8392 15700 8444 15706
rect 8444 15660 8524 15688
rect 8392 15642 8444 15648
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8220 15286 8340 15314
rect 8312 15162 8340 15286
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8206 15056 8262 15065
rect 8206 14991 8262 15000
rect 8300 15020 8352 15026
rect 8220 14958 8248 14991
rect 8300 14962 8352 14968
rect 8208 14952 8260 14958
rect 7654 14920 7710 14929
rect 8208 14894 8260 14900
rect 7654 14855 7710 14864
rect 7668 14822 7696 14855
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 7760 13530 7788 14758
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 8220 14074 8248 14758
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8312 13870 8340 14962
rect 8404 14890 8432 15438
rect 8496 15366 8524 15660
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7564 13524 7616 13530
rect 7748 13524 7800 13530
rect 7616 13484 7696 13512
rect 7564 13466 7616 13472
rect 7564 13388 7616 13394
rect 7668 13376 7696 13484
rect 7748 13466 7800 13472
rect 7668 13348 7788 13376
rect 7564 13330 7616 13336
rect 7576 12986 7604 13330
rect 7760 13274 7788 13348
rect 7760 13246 7880 13274
rect 7852 13190 7880 13246
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 8312 12714 8340 13806
rect 8496 13530 8524 14350
rect 8588 13954 8616 16102
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8772 15706 8800 15914
rect 8864 15706 8892 16118
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8864 15026 8892 15302
rect 8852 15020 8904 15026
rect 8772 14980 8852 15008
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8680 14414 8708 14894
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8588 13926 8708 13954
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7300 11342 7512 11370
rect 7484 11286 7512 11342
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7760 11234 7788 11766
rect 7944 11762 7972 12106
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7760 11218 7880 11234
rect 7760 11212 7892 11218
rect 7760 11206 7840 11212
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7116 9926 7144 10610
rect 7760 10606 7788 11206
rect 7840 11154 7892 11160
rect 8220 11150 8248 11698
rect 8404 11354 8432 11834
rect 8496 11694 8524 13466
rect 8588 13326 8616 13806
rect 8680 13734 8708 13926
rect 8772 13852 8800 14980
rect 8852 14962 8904 14968
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 14006 8892 14214
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8772 13824 8892 13852
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8772 11082 8800 12718
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7010 8936 7066 8945
rect 7010 8871 7066 8880
rect 6748 8486 6868 8514
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6748 3194 6776 8486
rect 7024 8362 7052 8871
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 6840 7750 6868 8298
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 5184 2746 5304 2774
rect 5184 2650 5212 2746
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 7116 2582 7144 9862
rect 7392 9586 7420 10474
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 9722 7512 10406
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7472 9716 7524 9722
rect 8312 9674 8340 10746
rect 8772 10606 8800 11018
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 7472 9658 7524 9664
rect 8220 9646 8340 9674
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 9110 7236 9386
rect 7564 9376 7616 9382
rect 7562 9344 7564 9353
rect 7616 9344 7618 9353
rect 7562 9279 7618 9288
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 8220 9042 8248 9646
rect 8404 9518 8432 10202
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8680 9586 8708 10066
rect 8772 10062 8800 10542
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8576 9104 8628 9110
rect 8496 9052 8576 9058
rect 8496 9046 8628 9052
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8496 9030 8616 9046
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7392 8430 7420 8910
rect 8404 8838 8432 8978
rect 8496 8974 8524 9030
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7654 8120 7710 8129
rect 7886 8112 8182 8132
rect 7654 8055 7710 8064
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7478 7420 7822
rect 7668 7818 7696 8055
rect 8220 8022 8248 8774
rect 8588 8634 8616 8910
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8680 8634 8708 8842
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 8588 7274 8616 8570
rect 8772 8566 8800 8910
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 8864 8022 8892 13824
rect 8956 11286 8984 20216
rect 9036 20198 9088 20204
rect 9036 19916 9088 19922
rect 9036 19858 9088 19864
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 9048 9110 9076 19858
rect 9140 19786 9168 20334
rect 9416 20058 9444 20538
rect 9508 20398 9536 22200
rect 9968 20602 9996 22200
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 10048 20528 10100 20534
rect 10100 20488 10364 20516
rect 10048 20470 10100 20476
rect 9864 20460 9916 20466
rect 9864 20402 9916 20408
rect 9496 20392 9548 20398
rect 9548 20352 9628 20380
rect 9496 20334 9548 20340
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9312 19984 9364 19990
rect 9312 19926 9364 19932
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9140 17678 9168 19246
rect 9232 18834 9260 19858
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9232 18630 9260 18770
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9140 17066 9168 17614
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9140 16454 9168 17002
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9128 16448 9180 16454
rect 9128 16390 9180 16396
rect 9140 16182 9168 16390
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 9140 15502 9168 16118
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 13870 9168 15438
rect 9232 15162 9260 16594
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9232 13938 9260 14350
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9218 13832 9274 13841
rect 9218 13767 9274 13776
rect 9232 12434 9260 13767
rect 9140 12406 9260 12434
rect 9140 10810 9168 12406
rect 9324 12238 9352 19926
rect 9416 17134 9444 19994
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9508 19514 9536 19722
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9508 19242 9536 19450
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9508 18834 9536 19178
rect 9600 18902 9628 20352
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9588 18896 9640 18902
rect 9588 18838 9640 18844
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9508 16674 9536 18566
rect 9600 18057 9628 18702
rect 9586 18048 9642 18057
rect 9586 17983 9642 17992
rect 9588 17060 9640 17066
rect 9588 17002 9640 17008
rect 9600 16794 9628 17002
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9508 16646 9628 16674
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9232 11762 9260 12038
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9416 11370 9444 14826
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 13734 9536 14214
rect 9600 13977 9628 16646
rect 9692 14804 9720 20198
rect 9876 17082 9904 20402
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 9968 20058 9996 20198
rect 9956 20052 10008 20058
rect 9956 19994 10008 20000
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9968 18834 9996 19654
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9968 17377 9996 18090
rect 9954 17368 10010 17377
rect 9954 17303 10010 17312
rect 9876 17054 9996 17082
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9784 16794 9812 16934
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9876 16046 9904 16934
rect 9968 16561 9996 17054
rect 9954 16552 10010 16561
rect 9954 16487 10010 16496
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 16114 9996 16390
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9864 16040 9916 16046
rect 9864 15982 9916 15988
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9772 14952 9824 14958
rect 9770 14920 9772 14929
rect 9824 14920 9826 14929
rect 9770 14855 9826 14864
rect 9692 14776 9812 14804
rect 9784 14550 9812 14776
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9678 14376 9734 14385
rect 9678 14311 9680 14320
rect 9732 14311 9734 14320
rect 9680 14282 9732 14288
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9586 13968 9642 13977
rect 9876 13938 9904 14214
rect 9586 13903 9642 13912
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9600 13326 9628 13806
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9600 12918 9628 13262
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9232 11342 9444 11370
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9140 10713 9168 10746
rect 9126 10704 9182 10713
rect 9126 10639 9182 10648
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 10266 9168 10406
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 9048 8838 9076 9046
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8864 7750 8892 7958
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 9232 5846 9260 11342
rect 9404 11280 9456 11286
rect 9404 11222 9456 11228
rect 9416 10538 9444 11222
rect 9508 11150 9536 12582
rect 9588 12232 9640 12238
rect 9588 12174 9640 12180
rect 9600 11370 9628 12174
rect 9692 11762 9720 12582
rect 9784 12442 9812 12786
rect 9772 12436 9824 12442
rect 9968 12434 9996 15030
rect 10060 12782 10088 20198
rect 10138 18320 10194 18329
rect 10138 18255 10194 18264
rect 10152 18086 10180 18255
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16658 10180 16934
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10138 16552 10194 16561
rect 10138 16487 10194 16496
rect 10232 16516 10284 16522
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 10152 12646 10180 16487
rect 10232 16458 10284 16464
rect 10244 16250 10272 16458
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 9772 12378 9824 12384
rect 9876 12406 9996 12434
rect 10048 12436 10100 12442
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9600 11354 9720 11370
rect 9600 11348 9732 11354
rect 9600 11342 9680 11348
rect 9680 11290 9732 11296
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9508 10606 9536 11086
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9324 10062 9352 10406
rect 9508 10266 9536 10406
rect 9600 10266 9628 10950
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9416 8906 9444 9590
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9600 8242 9628 9862
rect 9692 9586 9720 9862
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9692 8906 9720 9522
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9784 9178 9812 9318
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9876 8945 9904 12406
rect 10048 12378 10100 12384
rect 10060 12306 10088 12378
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9956 10464 10008 10470
rect 10152 10452 10180 10678
rect 10008 10424 10180 10452
rect 9956 10406 10008 10412
rect 10336 9674 10364 20488
rect 10428 20398 10456 22200
rect 10796 20398 10824 22200
rect 11256 20398 11284 22200
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 10416 20392 10468 20398
rect 10416 20334 10468 20340
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 11244 20392 11296 20398
rect 11244 20334 11296 20340
rect 11716 20380 11744 22200
rect 11980 20596 12032 20602
rect 11980 20538 12032 20544
rect 11796 20392 11848 20398
rect 11716 20352 11796 20380
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10428 17746 10456 18226
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10428 10742 10456 17274
rect 10520 11694 10548 20198
rect 10600 19984 10652 19990
rect 10600 19926 10652 19932
rect 10612 19514 10640 19926
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10704 19258 10732 19858
rect 10796 19310 10824 20334
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10612 19230 10732 19258
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10612 18748 10640 19230
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10704 18970 10732 19110
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10692 18760 10744 18766
rect 10612 18720 10692 18748
rect 10692 18702 10744 18708
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10612 16794 10640 18226
rect 10704 17542 10732 18702
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 10796 18086 10824 18226
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10690 17368 10746 17377
rect 10796 17338 10824 18022
rect 10690 17303 10746 17312
rect 10784 17332 10836 17338
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10600 16584 10652 16590
rect 10598 16552 10600 16561
rect 10652 16552 10654 16561
rect 10598 16487 10654 16496
rect 10600 15972 10652 15978
rect 10600 15914 10652 15920
rect 10612 15366 10640 15914
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10704 14906 10732 17303
rect 10784 17274 10836 17280
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10796 16590 10824 17138
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 10796 15502 10824 16526
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10796 15026 10824 15438
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10704 14878 10824 14906
rect 10888 14890 10916 19994
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 11072 17882 11100 18838
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10980 16726 11008 17818
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11072 16250 11100 16526
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10612 11540 10640 14758
rect 10796 13394 10824 14878
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10980 14822 11008 15438
rect 11072 15026 11100 15506
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11164 14906 11192 20198
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11256 19378 11284 19790
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11716 19514 11744 20352
rect 11796 20334 11848 20340
rect 11992 20330 12020 20538
rect 12084 20398 12112 22200
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12256 20528 12308 20534
rect 12256 20470 12308 20476
rect 12072 20392 12124 20398
rect 12072 20334 12124 20340
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11716 19174 11744 19314
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11808 18970 11836 19790
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11612 18284 11664 18290
rect 11612 18226 11664 18232
rect 11624 17882 11652 18226
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11610 17640 11666 17649
rect 11244 17604 11296 17610
rect 11610 17575 11612 17584
rect 11244 17546 11296 17552
rect 11664 17575 11666 17584
rect 11612 17546 11664 17552
rect 11256 17338 11284 17546
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11624 16794 11652 17070
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11256 15434 11284 16594
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11164 14878 11284 14906
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 11152 14544 11204 14550
rect 11152 14486 11204 14492
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10980 13734 11008 14418
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 11072 13190 11100 13874
rect 11164 13870 11192 14486
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10888 12889 10916 13126
rect 10874 12880 10930 12889
rect 10874 12815 10930 12824
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10796 11762 10824 12038
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10520 11512 10640 11540
rect 10520 11257 10548 11512
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10506 11248 10562 11257
rect 10506 11183 10562 11192
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10244 9646 10364 9674
rect 10140 9512 10192 9518
rect 10244 9500 10272 9646
rect 10192 9472 10272 9500
rect 10140 9454 10192 9460
rect 9862 8936 9918 8945
rect 9680 8900 9732 8906
rect 9862 8871 9918 8880
rect 9680 8842 9732 8848
rect 9692 8430 9720 8842
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8566 9812 8774
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9784 8242 9812 8366
rect 9600 8214 9812 8242
rect 9600 7410 9628 8214
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 10520 6458 10548 11183
rect 10612 10674 10640 11290
rect 10704 11218 10732 11698
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10784 11144 10836 11150
rect 10888 11132 10916 12174
rect 11072 11665 11100 12310
rect 11058 11656 11114 11665
rect 11256 11642 11284 14878
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11624 12442 11652 12786
rect 11612 12436 11664 12442
rect 11716 12434 11744 14758
rect 11808 14074 11836 18702
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11808 13734 11836 14010
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11808 12782 11836 13126
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11716 12406 11836 12434
rect 11612 12378 11664 12384
rect 11624 12238 11652 12378
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11716 11694 11744 12242
rect 11704 11688 11756 11694
rect 11256 11614 11376 11642
rect 11704 11630 11756 11636
rect 11058 11591 11114 11600
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11256 11286 11284 11494
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 10836 11104 10916 11132
rect 10784 11086 10836 11092
rect 11152 11008 11204 11014
rect 11348 10996 11376 11614
rect 11808 11354 11836 12406
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11152 10950 11204 10956
rect 11256 10968 11376 10996
rect 11164 10810 11192 10950
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 11256 9654 11284 10968
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11716 10198 11744 10746
rect 11704 10192 11756 10198
rect 11704 10134 11756 10140
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10796 8945 10824 8978
rect 10782 8936 10838 8945
rect 10782 8871 10838 8880
rect 11256 8498 11284 9590
rect 11336 8968 11388 8974
rect 11334 8936 11336 8945
rect 11388 8936 11390 8945
rect 11334 8871 11390 8880
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11808 6662 11836 11290
rect 11900 9178 11928 20198
rect 12084 19446 12112 20334
rect 12072 19440 12124 19446
rect 12072 19382 12124 19388
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 12084 17882 12112 18022
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11992 15162 12020 15438
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11978 15056 12034 15065
rect 12176 15042 12204 20470
rect 12268 18766 12296 20470
rect 12544 20398 12572 22200
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12348 20256 12400 20262
rect 12348 20198 12400 20204
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12268 18193 12296 18362
rect 12254 18184 12310 18193
rect 12254 18119 12310 18128
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 11978 14991 11980 15000
rect 12032 14991 12034 15000
rect 12084 15014 12204 15042
rect 11980 14962 12032 14968
rect 12084 12102 12112 15014
rect 12164 14952 12216 14958
rect 12164 14894 12216 14900
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11992 10810 12020 11698
rect 12176 11642 12204 14894
rect 12268 13802 12296 15098
rect 12360 14226 12388 20198
rect 12440 19984 12492 19990
rect 12440 19926 12492 19932
rect 12452 18970 12480 19926
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12452 18193 12480 18770
rect 12532 18352 12584 18358
rect 12530 18320 12532 18329
rect 12584 18320 12586 18329
rect 12530 18255 12586 18264
rect 12438 18184 12494 18193
rect 12438 18119 12494 18128
rect 12452 18086 12480 18119
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12636 14385 12664 20198
rect 12728 20058 12756 20334
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12820 19922 12848 20470
rect 12912 20398 12940 22200
rect 13372 20602 13400 22200
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13728 20528 13780 20534
rect 13832 20516 13860 22200
rect 14200 20534 14228 22200
rect 14660 20534 14688 22200
rect 13780 20488 13860 20516
rect 14188 20528 14240 20534
rect 13728 20470 13780 20476
rect 14188 20470 14240 20476
rect 14648 20528 14700 20534
rect 15120 20516 15148 22200
rect 15488 20534 15516 22200
rect 15948 20602 15976 22200
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15200 20528 15252 20534
rect 15120 20488 15200 20516
rect 14648 20470 14700 20476
rect 15200 20470 15252 20476
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 16316 20466 16344 22200
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16776 20398 16804 22200
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12820 19394 12848 19858
rect 12912 19514 12940 20334
rect 14004 20324 14056 20330
rect 14004 20266 14056 20272
rect 14280 20324 14332 20330
rect 14832 20324 14884 20330
rect 14280 20266 14332 20272
rect 14384 20284 14832 20312
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12728 19366 12848 19394
rect 12728 18426 12756 19366
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12820 18766 12848 19178
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12912 17814 12940 18770
rect 12900 17808 12952 17814
rect 12900 17750 12952 17756
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12728 17066 12756 17682
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12912 16794 12940 17750
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12820 14550 12848 14962
rect 12808 14544 12860 14550
rect 12808 14486 12860 14492
rect 12622 14376 12678 14385
rect 12622 14311 12678 14320
rect 12360 14198 12480 14226
rect 12256 13796 12308 13802
rect 12256 13738 12308 13744
rect 12452 13002 12480 14198
rect 12636 13870 12664 14311
rect 12820 13938 12848 14486
rect 13004 13938 13032 19654
rect 13372 19334 13400 19790
rect 13372 19310 13492 19334
rect 13372 19306 13504 19310
rect 13452 19304 13504 19306
rect 13452 19246 13504 19252
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 13188 18306 13216 18770
rect 13096 18290 13216 18306
rect 13084 18284 13216 18290
rect 13136 18278 13216 18284
rect 13450 18320 13506 18329
rect 13450 18255 13506 18264
rect 13084 18226 13136 18232
rect 13464 18086 13492 18255
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13280 16674 13308 17138
rect 13096 16658 13308 16674
rect 13084 16652 13308 16658
rect 13136 16646 13308 16652
rect 13084 16594 13136 16600
rect 13280 15978 13308 16646
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 13372 15858 13400 18022
rect 13556 17202 13584 19790
rect 13648 18136 13676 19858
rect 14016 19802 14044 20266
rect 14096 20256 14148 20262
rect 14148 20216 14228 20244
rect 14096 20198 14148 20204
rect 14200 20058 14228 20216
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14016 19774 14136 19802
rect 14108 19718 14136 19774
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14016 19394 14044 19654
rect 14016 19366 14228 19394
rect 14200 19310 14228 19366
rect 13912 19304 13964 19310
rect 14188 19304 14240 19310
rect 13964 19252 14044 19258
rect 13912 19246 14044 19252
rect 14188 19246 14240 19252
rect 13820 19236 13872 19242
rect 13924 19230 14044 19246
rect 13820 19178 13872 19184
rect 13728 19168 13780 19174
rect 13728 19110 13780 19116
rect 13740 18834 13768 19110
rect 13728 18828 13780 18834
rect 13728 18770 13780 18776
rect 13832 18358 13860 19178
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13820 18148 13872 18154
rect 13648 18108 13820 18136
rect 13820 18090 13872 18096
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 16794 13768 16934
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13832 16674 13860 18090
rect 13924 17338 13952 19110
rect 14016 18290 14044 19230
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14200 18358 14228 18702
rect 14188 18352 14240 18358
rect 14188 18294 14240 18300
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14016 17218 14044 18226
rect 14200 18154 14228 18294
rect 14292 18222 14320 20266
rect 14384 18902 14412 20284
rect 14832 20266 14884 20272
rect 15476 20324 15528 20330
rect 15476 20266 15528 20272
rect 15844 20324 15896 20330
rect 15844 20266 15896 20272
rect 15936 20324 15988 20330
rect 15936 20266 15988 20272
rect 16212 20324 16264 20330
rect 16212 20266 16264 20272
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 14740 19916 14792 19922
rect 14740 19858 14792 19864
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14372 18896 14424 18902
rect 14372 18838 14424 18844
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14384 18290 14412 18702
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 14568 17882 14596 19722
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14660 18902 14688 19382
rect 14752 18970 14780 19858
rect 14844 19786 14872 19858
rect 14832 19780 14884 19786
rect 14832 19722 14884 19728
rect 14924 19712 14976 19718
rect 14830 19680 14886 19689
rect 14924 19654 14976 19660
rect 15108 19712 15160 19718
rect 15108 19654 15160 19660
rect 14830 19615 14886 19624
rect 14844 19242 14872 19615
rect 14936 19446 14964 19654
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 15120 19310 15148 19654
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 14832 19236 14884 19242
rect 15212 19224 15240 19994
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15292 19712 15344 19718
rect 15396 19689 15424 19858
rect 15292 19654 15344 19660
rect 15382 19680 15438 19689
rect 15304 19514 15332 19654
rect 15382 19615 15438 19624
rect 15488 19514 15516 20266
rect 15856 20058 15884 20266
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15292 19236 15344 19242
rect 15212 19196 15292 19224
rect 14832 19178 14884 19184
rect 15292 19178 15344 19184
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 14740 18964 14792 18970
rect 14740 18906 14792 18912
rect 14648 18896 14700 18902
rect 14648 18838 14700 18844
rect 14646 18320 14702 18329
rect 14646 18255 14702 18264
rect 14660 18154 14688 18255
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 13924 17190 14044 17218
rect 13924 16998 13952 17190
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13280 15830 13400 15858
rect 13740 16646 13860 16674
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12992 13932 13044 13938
rect 12992 13874 13044 13880
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12992 13796 13044 13802
rect 12992 13738 13044 13744
rect 13004 13190 13032 13738
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 13096 13326 13124 13670
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 12360 12974 12480 13002
rect 13004 12986 13032 13126
rect 12992 12980 13044 12986
rect 12360 12968 12388 12974
rect 12268 12940 12388 12968
rect 12268 12434 12296 12940
rect 12992 12922 13044 12928
rect 13280 12434 13308 15830
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 13556 15434 13584 15574
rect 13544 15428 13596 15434
rect 13544 15370 13596 15376
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14074 13584 14758
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13452 13728 13504 13734
rect 13452 13670 13504 13676
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13372 12918 13400 13330
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13464 12434 13492 13670
rect 12268 12406 12388 12434
rect 12176 11614 12296 11642
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12176 11354 12204 11494
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 12084 10130 12112 10406
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 12176 8838 12204 9386
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12268 7818 12296 11614
rect 12360 11082 12388 12406
rect 13188 12406 13308 12434
rect 13372 12406 13492 12434
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11626 12480 12038
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12452 11014 12480 11086
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10606 12480 10950
rect 12348 10600 12400 10606
rect 12346 10568 12348 10577
rect 12440 10600 12492 10606
rect 12400 10568 12402 10577
rect 12440 10542 12492 10548
rect 12346 10503 12402 10512
rect 12452 10062 12480 10542
rect 12544 10266 12572 11494
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12912 10538 12940 10950
rect 13096 10742 13124 11562
rect 13084 10736 13136 10742
rect 13084 10678 13136 10684
rect 13096 10606 13124 10678
rect 13084 10600 13136 10606
rect 12990 10568 13046 10577
rect 12900 10532 12952 10538
rect 13084 10542 13136 10548
rect 12990 10503 13046 10512
rect 12900 10474 12952 10480
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12544 8634 12572 9658
rect 12636 9450 12664 9998
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12820 9382 12848 9998
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12912 9178 12940 10066
rect 13004 9994 13032 10503
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13096 9926 13124 10542
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 9586 13124 9862
rect 13188 9722 13216 12406
rect 13372 11778 13400 12406
rect 13556 11914 13584 13874
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13648 12986 13676 13262
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13740 12753 13768 16646
rect 13924 16590 13952 16934
rect 13820 16584 13872 16590
rect 13820 16526 13872 16532
rect 13912 16584 13964 16590
rect 13912 16526 13964 16532
rect 13832 16250 13860 16526
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13832 15502 13860 16186
rect 13924 16046 13952 16526
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13924 14414 13952 15982
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14016 14550 14044 14962
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 14016 14346 14044 14486
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 14108 14226 14136 17614
rect 14292 16454 14320 17682
rect 14372 17604 14424 17610
rect 14372 17546 14424 17552
rect 14384 17338 14412 17546
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 13924 14198 14136 14226
rect 13726 12744 13782 12753
rect 13726 12679 13782 12688
rect 13740 12170 13768 12679
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13832 12238 13860 12378
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13464 11898 13584 11914
rect 13452 11892 13584 11898
rect 13504 11886 13584 11892
rect 13452 11834 13504 11840
rect 13372 11750 13492 11778
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13280 10266 13308 10474
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12728 8634 12756 8978
rect 13280 8974 13308 9522
rect 13464 9178 13492 11750
rect 13556 11354 13584 11886
rect 13832 11694 13860 12038
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13832 11014 13860 11222
rect 13924 11218 13952 14198
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14016 12442 14044 12582
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14108 11898 14136 13194
rect 14292 12714 14320 14554
rect 14384 12986 14412 16934
rect 14568 15638 14596 16934
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 14186 12608 14242 12617
rect 14186 12543 14242 12552
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13924 10470 13952 11154
rect 14016 10606 14044 11154
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 13556 10062 13584 10406
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 14108 8362 14136 10406
rect 14200 10130 14228 12543
rect 14384 12102 14412 12786
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14280 11620 14332 11626
rect 14280 11562 14332 11568
rect 14292 11150 14320 11562
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14292 10674 14320 11086
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 14292 10266 14320 10406
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14384 10062 14412 10202
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14476 8820 14504 15302
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14568 13258 14596 14894
rect 14660 13410 14688 18090
rect 14752 17678 14780 18090
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 15396 17338 15424 17682
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14752 16114 14780 16934
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 15304 15978 15332 17138
rect 15396 16998 15424 17274
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15304 15502 15332 15914
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15396 15434 15424 16594
rect 15474 16552 15530 16561
rect 15474 16487 15530 16496
rect 15488 15978 15516 16487
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15384 15428 15436 15434
rect 15384 15370 15436 15376
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15396 14890 15424 15030
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 15384 14884 15436 14890
rect 15384 14826 15436 14832
rect 14752 14074 14780 14826
rect 15580 14770 15608 19790
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15672 18222 15700 19110
rect 15948 18970 15976 20266
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16040 19174 16068 20198
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16132 19446 16160 19858
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 16224 18873 16252 20266
rect 16684 20097 16712 20266
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16670 20088 16726 20097
rect 16670 20023 16726 20032
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16210 18864 16266 18873
rect 15936 18828 15988 18834
rect 16210 18799 16266 18808
rect 15936 18770 15988 18776
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15764 18290 15792 18566
rect 15856 18426 15884 18702
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 15844 18080 15896 18086
rect 15948 18068 15976 18770
rect 15896 18040 15976 18068
rect 15844 18022 15896 18028
rect 15948 17678 15976 18040
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16132 17882 16160 18022
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16224 17202 16252 17478
rect 16316 17338 16344 19246
rect 16408 17882 16436 19858
rect 16500 19666 16528 19858
rect 16776 19825 16804 20198
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16762 19816 16818 19825
rect 16672 19780 16724 19786
rect 16762 19751 16818 19760
rect 16672 19722 16724 19728
rect 16500 19638 16620 19666
rect 16592 18630 16620 19638
rect 16684 19310 16712 19722
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16684 18902 16712 19110
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16684 18465 16712 18838
rect 16868 18834 16896 19994
rect 17236 19990 17264 22200
rect 17604 19990 17632 22200
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17972 20602 18000 20742
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17224 19984 17276 19990
rect 17224 19926 17276 19932
rect 17592 19984 17644 19990
rect 17592 19926 17644 19932
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17144 19718 17172 19790
rect 17696 19718 17724 20266
rect 18064 19990 18092 22200
rect 18524 21298 18552 22200
rect 18524 21270 18644 21298
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 18052 19984 18104 19990
rect 18052 19926 18104 19932
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17144 19514 17172 19654
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17972 19394 18000 19858
rect 18052 19780 18104 19786
rect 18052 19722 18104 19728
rect 17604 19366 18000 19394
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 16948 18760 17000 18766
rect 16762 18728 16818 18737
rect 16948 18702 17000 18708
rect 16762 18663 16818 18672
rect 16670 18456 16726 18465
rect 16670 18391 16726 18400
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16500 17542 16528 18022
rect 16592 17610 16620 18022
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15752 16448 15804 16454
rect 15948 16402 15976 16526
rect 15804 16396 15976 16402
rect 15752 16390 15976 16396
rect 15764 16374 15976 16390
rect 15764 16046 15792 16374
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15162 15700 15846
rect 16132 15502 16160 16186
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16408 15638 16436 16050
rect 16500 16046 16528 17070
rect 16592 16794 16620 17070
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 16396 15632 16448 15638
rect 16396 15574 16448 15580
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16500 15162 16528 15982
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15396 14742 15608 14770
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15212 13734 15240 13806
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14660 13382 14872 13410
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14568 11218 14596 13194
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14568 9178 14596 9386
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14648 8832 14700 8838
rect 14476 8792 14648 8820
rect 14648 8774 14700 8780
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 14660 6186 14688 8774
rect 14752 7546 14780 12922
rect 14844 12753 14872 13382
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14936 12850 14964 13126
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14830 12744 14886 12753
rect 14830 12679 14886 12688
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15120 11801 15148 12242
rect 15106 11792 15162 11801
rect 15106 11727 15162 11736
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15016 11280 15068 11286
rect 15016 11222 15068 11228
rect 15028 11150 15056 11222
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 14844 11014 14872 11086
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14844 10606 14872 10950
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15106 9888 15162 9897
rect 15106 9823 15162 9832
rect 15120 9722 15148 9823
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15212 8090 15240 13670
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15304 12238 15332 12786
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15396 11665 15424 14742
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15488 14056 15516 14486
rect 15488 14028 15608 14056
rect 15580 13938 15608 14028
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15672 13802 15700 14758
rect 15764 14618 15792 14962
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 16316 14618 16344 14758
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 15764 13462 15792 14554
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15856 13870 15884 14214
rect 16316 13938 16344 14350
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15488 11898 15516 13398
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15764 11694 15792 12582
rect 16132 12434 16160 13806
rect 16500 13734 16528 14214
rect 16592 13802 16620 14418
rect 16684 14346 16712 14554
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16776 12434 16804 18663
rect 16960 18426 16988 18702
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16960 18290 16988 18362
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 16868 17542 16896 17750
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16868 13190 16896 17478
rect 16960 16250 16988 18226
rect 17144 17338 17172 19246
rect 17500 19168 17552 19174
rect 17500 19110 17552 19116
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17328 18154 17356 18566
rect 17316 18148 17368 18154
rect 17316 18090 17368 18096
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 17236 17270 17264 17614
rect 17328 17610 17356 18090
rect 17512 17882 17540 19110
rect 17604 18970 17632 19366
rect 18064 19310 18092 19722
rect 18156 19446 18184 20266
rect 18432 19700 18460 20334
rect 18616 20330 18644 21270
rect 18892 20602 18920 22200
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 18984 20330 19012 22607
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 19798 22264 19854 22273
rect 19352 20466 19380 22200
rect 19720 21842 19748 22200
rect 19798 22199 19854 22208
rect 20166 22200 20222 23000
rect 20626 22200 20682 23000
rect 20994 22200 21050 23000
rect 21454 22200 21510 23000
rect 21914 22200 21970 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 19628 21814 19748 21842
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19628 20398 19656 21814
rect 19706 21720 19762 21729
rect 19706 21655 19762 21664
rect 19720 20534 19748 21655
rect 19708 20528 19760 20534
rect 19708 20470 19760 20476
rect 19616 20392 19668 20398
rect 19616 20334 19668 20340
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 18604 20324 18656 20330
rect 18604 20266 18656 20272
rect 18972 20324 19024 20330
rect 18972 20266 19024 20272
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 18696 20256 18748 20262
rect 18748 20216 18828 20244
rect 18696 20198 18748 20204
rect 18800 20058 18828 20216
rect 19062 20088 19118 20097
rect 18788 20052 18840 20058
rect 19168 20058 19196 20266
rect 19248 20256 19300 20262
rect 19300 20216 19380 20244
rect 19248 20198 19300 20204
rect 19062 20023 19118 20032
rect 19156 20052 19208 20058
rect 18788 19994 18840 20000
rect 19076 19990 19104 20023
rect 19156 19994 19208 20000
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 18892 19718 18920 19858
rect 18788 19712 18840 19718
rect 18432 19672 18644 19700
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18616 19496 18644 19672
rect 18788 19654 18840 19660
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18800 19514 18828 19654
rect 18340 19468 18644 19496
rect 18788 19508 18840 19514
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17696 18834 17724 19110
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17788 17882 17816 19178
rect 18156 18970 18184 19246
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18248 18834 18276 19314
rect 18340 19174 18368 19468
rect 18788 19450 18840 19456
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18236 18828 18288 18834
rect 18236 18770 18288 18776
rect 18248 18714 18276 18770
rect 18432 18737 18460 19110
rect 18510 19000 18566 19009
rect 18510 18935 18566 18944
rect 18524 18902 18552 18935
rect 18512 18896 18564 18902
rect 18512 18838 18564 18844
rect 18156 18686 18276 18714
rect 18418 18728 18474 18737
rect 18050 18592 18106 18601
rect 18050 18527 18106 18536
rect 18064 18358 18092 18527
rect 18156 18426 18184 18686
rect 18418 18663 18474 18672
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18144 18420 18196 18426
rect 18144 18362 18196 18368
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17316 17604 17368 17610
rect 17316 17546 17368 17552
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17052 16794 17080 16934
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 17144 16726 17172 17002
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17132 16720 17184 16726
rect 17132 16662 17184 16668
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17236 14822 17264 16934
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17328 15162 17356 16594
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17420 15910 17448 16390
rect 17512 15978 17540 16526
rect 17604 16114 17632 17274
rect 17696 16998 17724 17614
rect 17880 17270 17908 17682
rect 18064 17270 18092 18294
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18432 17882 18460 18022
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 18616 17814 18644 19314
rect 18972 19304 19024 19310
rect 18694 19272 18750 19281
rect 18972 19246 19024 19252
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 18694 19207 18750 19216
rect 18604 17808 18656 17814
rect 18604 17750 18656 17756
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17592 16108 17644 16114
rect 17592 16050 17644 16056
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17420 14346 17448 15846
rect 17512 15706 17540 15914
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17604 15026 17632 15846
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17512 14550 17540 14758
rect 17500 14544 17552 14550
rect 17500 14486 17552 14492
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17604 13326 17632 13738
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 16856 13184 16908 13190
rect 16856 13126 16908 13132
rect 16868 12782 16896 13126
rect 16948 12912 17000 12918
rect 17880 12889 17908 17206
rect 18156 17066 18184 17478
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18708 17354 18736 19207
rect 18880 19168 18932 19174
rect 18878 19136 18880 19145
rect 18932 19136 18934 19145
rect 18878 19071 18934 19080
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18800 18358 18828 18770
rect 18788 18352 18840 18358
rect 18788 18294 18840 18300
rect 18892 18222 18920 18838
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18616 17326 18736 17354
rect 18616 17270 18644 17326
rect 18604 17264 18656 17270
rect 18604 17206 18656 17212
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17972 15026 18000 15370
rect 18064 15162 18092 16662
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 18156 14906 18184 17002
rect 18708 16794 18736 17070
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18892 16726 18920 18158
rect 18984 17882 19012 19246
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 19076 17338 19104 19246
rect 19168 17746 19196 19858
rect 19260 19378 19288 19858
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19246 19136 19302 19145
rect 19246 19071 19302 19080
rect 19260 18290 19288 19071
rect 19352 18426 19380 20216
rect 19444 20058 19472 20266
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19444 18902 19472 19382
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19536 18306 19564 19654
rect 19628 19514 19656 19858
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19616 19168 19668 19174
rect 19614 19136 19616 19145
rect 19668 19136 19670 19145
rect 19614 19071 19670 19080
rect 19616 18896 19668 18902
rect 19616 18838 19668 18844
rect 19628 18630 19656 18838
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19248 18284 19300 18290
rect 19536 18278 19656 18306
rect 19248 18226 19300 18232
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19444 17746 19472 18022
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19156 17536 19208 17542
rect 19156 17478 19208 17484
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18880 16720 18932 16726
rect 18880 16662 18932 16668
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 17972 14878 18184 14906
rect 16948 12854 17000 12860
rect 17866 12880 17922 12889
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 16132 12406 16436 12434
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16132 12102 16160 12242
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15856 11898 15884 12038
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 16040 11830 16068 12038
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 15752 11688 15804 11694
rect 15382 11656 15438 11665
rect 15752 11630 15804 11636
rect 15382 11591 15438 11600
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15304 9722 15332 10406
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15396 9382 15424 11290
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15488 10538 15516 10610
rect 15476 10532 15528 10538
rect 15476 10474 15528 10480
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 10198 15792 10406
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15856 10130 15884 10610
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 15948 10266 15976 10474
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15580 9722 15608 10066
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15856 9654 15884 10066
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15488 8974 15516 9522
rect 15948 9178 15976 10202
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 16132 8634 16160 12038
rect 16408 10674 16436 12406
rect 16684 12406 16804 12434
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 9178 16252 10406
rect 16408 9518 16436 10610
rect 16684 10033 16712 12406
rect 16960 12238 16988 12854
rect 17866 12815 17922 12824
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16776 11898 16804 12174
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 17052 11778 17080 12718
rect 17868 12300 17920 12306
rect 17972 12288 18000 14878
rect 18984 14822 19012 17070
rect 19168 16794 19196 17478
rect 19628 17218 19656 18278
rect 19536 17190 19656 17218
rect 19536 16998 19564 17190
rect 19616 17060 19668 17066
rect 19616 17002 19668 17008
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19628 16794 19656 17002
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19628 16590 19656 16730
rect 19616 16584 19668 16590
rect 19616 16526 19668 16532
rect 19720 16402 19748 20334
rect 19812 20262 19840 22199
rect 20180 20602 20208 22200
rect 20442 21312 20498 21321
rect 20442 21247 20498 21256
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 20456 20534 20484 21247
rect 20534 20768 20590 20777
rect 20534 20703 20590 20712
rect 20548 20602 20576 20703
rect 20536 20596 20588 20602
rect 20536 20538 20588 20544
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 20444 20324 20496 20330
rect 20444 20266 20496 20272
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 20456 20058 20484 20266
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20640 19990 20668 22200
rect 21008 20482 21036 22200
rect 21468 20806 21496 22200
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 20916 20454 21036 20482
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19812 18902 19840 19314
rect 19996 19310 20024 19858
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 19800 18896 19852 18902
rect 19800 18838 19852 18844
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19812 18358 19840 18566
rect 19800 18352 19852 18358
rect 19800 18294 19852 18300
rect 19536 16374 19748 16402
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19352 15570 19380 15982
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19076 14958 19104 15438
rect 19064 14952 19116 14958
rect 19352 14906 19380 15506
rect 19444 15366 19472 15506
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19064 14894 19116 14900
rect 19168 14878 19380 14906
rect 18144 14816 18196 14822
rect 18144 14758 18196 14764
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18156 14278 18184 14758
rect 18696 14340 18748 14346
rect 19168 14328 19196 14878
rect 19340 14816 19392 14822
rect 19260 14764 19340 14770
rect 19260 14758 19392 14764
rect 19260 14742 19380 14758
rect 19260 14328 19288 14742
rect 19444 14634 19472 15302
rect 19352 14618 19472 14634
rect 19340 14612 19472 14618
rect 19392 14606 19472 14612
rect 19340 14554 19392 14560
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19444 14346 19472 14418
rect 18696 14282 18748 14288
rect 19076 14300 19196 14328
rect 19252 14300 19288 14328
rect 19432 14340 19484 14346
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18328 12912 18380 12918
rect 18326 12880 18328 12889
rect 18380 12880 18382 12889
rect 18326 12815 18382 12824
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 17920 12260 18000 12288
rect 18052 12300 18104 12306
rect 17868 12242 17920 12248
rect 18052 12242 18104 12248
rect 16960 11750 17080 11778
rect 17958 11792 18014 11801
rect 16960 11694 16988 11750
rect 17958 11727 18014 11736
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 17774 11656 17830 11665
rect 16776 11014 16804 11630
rect 17774 11591 17830 11600
rect 17868 11620 17920 11626
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17052 11354 17080 11494
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16868 11150 16896 11290
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16776 10470 16804 10950
rect 17052 10674 17080 11290
rect 17788 11150 17816 11591
rect 17868 11562 17920 11568
rect 17880 11218 17908 11562
rect 17972 11336 18000 11727
rect 18064 11558 18092 12242
rect 18432 12238 18460 12718
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18616 12374 18644 12582
rect 18708 12481 18736 14282
rect 19076 13734 19104 14300
rect 19252 14090 19280 14300
rect 19432 14282 19484 14288
rect 19252 14062 19288 14090
rect 19064 13728 19116 13734
rect 19064 13670 19116 13676
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18788 12640 18840 12646
rect 18788 12582 18840 12588
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18694 12472 18750 12481
rect 18800 12442 18828 12582
rect 18694 12407 18750 12416
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18696 12368 18748 12374
rect 18892 12322 18920 12582
rect 18984 12434 19012 13330
rect 19156 12436 19208 12442
rect 18984 12406 19104 12434
rect 18748 12316 18828 12322
rect 18696 12310 18828 12316
rect 18708 12294 18828 12310
rect 18892 12294 19012 12322
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18420 12232 18472 12238
rect 18696 12232 18748 12238
rect 18472 12180 18644 12186
rect 18420 12174 18644 12180
rect 18696 12174 18748 12180
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17972 11308 18092 11336
rect 17958 11248 18014 11257
rect 17868 11212 17920 11218
rect 17958 11183 17960 11192
rect 17868 11154 17920 11160
rect 18012 11183 18014 11192
rect 17960 11154 18012 11160
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17880 11098 17908 11154
rect 17604 11014 17632 11086
rect 17880 11070 18000 11098
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 17144 10606 17172 10950
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17236 10674 17264 10746
rect 17224 10668 17276 10674
rect 17224 10610 17276 10616
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16670 10024 16726 10033
rect 16670 9959 16726 9968
rect 16684 9654 16712 9959
rect 16960 9654 16988 10474
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 17144 10198 17172 10406
rect 17604 10266 17632 10950
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 16684 9518 16712 9590
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 9178 16344 9318
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 17144 9042 17172 10134
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9897 17264 10066
rect 17222 9888 17278 9897
rect 17222 9823 17278 9832
rect 17592 9444 17644 9450
rect 17592 9386 17644 9392
rect 17604 9042 17632 9386
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16316 8566 16344 8774
rect 16304 8560 16356 8566
rect 16304 8502 16356 8508
rect 16592 8498 16620 8774
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16868 8362 16896 8910
rect 17144 8498 17172 8978
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 16856 8356 16908 8362
rect 16856 8298 16908 8304
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 16868 7546 16896 8298
rect 17696 7886 17724 8298
rect 17972 7886 18000 11070
rect 18064 8090 18092 11308
rect 18156 10810 18184 12174
rect 18432 12158 18644 12174
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18616 11898 18644 12158
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18524 11529 18552 11766
rect 18510 11520 18566 11529
rect 18510 11455 18566 11464
rect 18708 11082 18736 12174
rect 18800 11626 18828 12294
rect 18878 12200 18934 12209
rect 18878 12135 18934 12144
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18892 11354 18920 12135
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18144 10804 18196 10810
rect 18144 10746 18196 10752
rect 18892 10674 18920 10950
rect 18984 10810 19012 12294
rect 19076 12102 19104 12406
rect 19156 12378 19208 12384
rect 19168 12345 19196 12378
rect 19154 12336 19210 12345
rect 19154 12271 19210 12280
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19064 11824 19116 11830
rect 19168 11812 19196 12174
rect 19116 11784 19196 11812
rect 19064 11766 19116 11772
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11354 19104 11494
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19168 11286 19196 11784
rect 19260 11744 19288 14062
rect 19338 13968 19394 13977
rect 19338 13903 19394 13912
rect 19352 13870 19380 13903
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 19430 12744 19486 12753
rect 19430 12679 19486 12688
rect 19252 11716 19288 11744
rect 19252 11642 19280 11716
rect 19252 11614 19288 11642
rect 19260 11286 19288 11614
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 19076 10713 19104 10746
rect 19062 10704 19118 10713
rect 18880 10668 18932 10674
rect 19168 10674 19196 11222
rect 19062 10639 19118 10648
rect 19156 10668 19208 10674
rect 18880 10610 18932 10616
rect 19156 10610 19208 10616
rect 19352 10606 19380 11494
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19340 10192 19392 10198
rect 19338 10160 19340 10169
rect 19392 10160 19394 10169
rect 19338 10095 19394 10104
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9382 18184 9862
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 9110 18276 9318
rect 18236 9104 18288 9110
rect 18420 9104 18472 9110
rect 18288 9052 18420 9058
rect 18236 9046 18472 9052
rect 18144 9036 18196 9042
rect 18248 9030 18460 9046
rect 18144 8978 18196 8984
rect 18156 8566 18184 8978
rect 18602 8936 18658 8945
rect 18602 8871 18604 8880
rect 18656 8871 18658 8880
rect 18604 8842 18656 8848
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18892 8498 18920 8774
rect 19352 8634 19380 9998
rect 19444 9722 19472 12679
rect 19536 11898 19564 16374
rect 19708 15972 19760 15978
rect 19708 15914 19760 15920
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19628 15366 19656 15642
rect 19720 15502 19748 15914
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19720 14822 19748 14894
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19708 14544 19760 14550
rect 19708 14486 19760 14492
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19628 13870 19656 14350
rect 19616 13864 19668 13870
rect 19616 13806 19668 13812
rect 19628 13530 19656 13806
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19614 13288 19670 13297
rect 19614 13223 19616 13232
rect 19668 13223 19670 13232
rect 19616 13194 19668 13200
rect 19616 12980 19668 12986
rect 19616 12922 19668 12928
rect 19628 12646 19656 12922
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19616 12436 19668 12442
rect 19720 12434 19748 14486
rect 19668 12406 19748 12434
rect 19616 12378 19668 12384
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19522 11792 19578 11801
rect 19522 11727 19578 11736
rect 19536 11286 19564 11727
rect 19720 11354 19748 12106
rect 19708 11348 19760 11354
rect 19708 11290 19760 11296
rect 19524 11280 19576 11286
rect 19524 11222 19576 11228
rect 19708 11008 19760 11014
rect 19708 10950 19760 10956
rect 19720 10742 19748 10950
rect 19708 10736 19760 10742
rect 19708 10678 19760 10684
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19444 9178 19472 9386
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19536 9110 19564 10542
rect 19628 10266 19656 10542
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19524 9104 19576 9110
rect 19524 9046 19576 9052
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18984 8090 19012 8230
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 11532 2650 11560 2926
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 15580 2650 15608 2858
rect 18064 2774 18092 8026
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18156 2854 18184 7822
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19352 6866 19380 7278
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 17972 2746 18092 2774
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 17972 2582 18000 2746
rect 19444 2650 19472 8978
rect 19628 6866 19656 9318
rect 19720 8090 19748 10406
rect 19708 8084 19760 8090
rect 19708 8026 19760 8032
rect 19812 7274 19840 18294
rect 19904 18222 19932 19110
rect 19996 18222 20024 19110
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19996 17814 20024 18022
rect 19984 17808 20036 17814
rect 19984 17750 20036 17756
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19904 15706 19932 16934
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19904 15162 19932 15642
rect 19892 15156 19944 15162
rect 19892 15098 19944 15104
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19904 9110 19932 14758
rect 19996 14550 20024 17750
rect 19984 14544 20036 14550
rect 19984 14486 20036 14492
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 19996 12986 20024 14350
rect 20088 13530 20116 14418
rect 20076 13524 20128 13530
rect 20076 13466 20128 13472
rect 20180 13258 20208 14418
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19984 12368 20036 12374
rect 19982 12336 19984 12345
rect 20036 12336 20038 12345
rect 19982 12271 20038 12280
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19996 11150 20024 11698
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20076 11552 20128 11558
rect 20074 11520 20076 11529
rect 20128 11520 20130 11529
rect 20074 11455 20130 11464
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 20180 10810 20208 11562
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19892 9104 19944 9110
rect 19892 9046 19944 9052
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19800 7268 19852 7274
rect 19800 7210 19852 7216
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19904 3942 19932 8910
rect 19996 8634 20024 10066
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19982 8528 20038 8537
rect 19982 8463 20038 8472
rect 19996 8294 20024 8463
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19996 3466 20024 8230
rect 20088 8022 20116 9318
rect 20180 9178 20208 10406
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20180 8090 20208 8774
rect 20272 8090 20300 19654
rect 20364 19446 20392 19858
rect 20352 19440 20404 19446
rect 20352 19382 20404 19388
rect 20732 19281 20760 20334
rect 20916 19990 20944 20454
rect 21178 20360 21234 20369
rect 20996 20324 21048 20330
rect 21178 20295 21180 20304
rect 20996 20266 21048 20272
rect 21232 20295 21234 20304
rect 21180 20266 21232 20272
rect 20904 19984 20956 19990
rect 20904 19926 20956 19932
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20718 19272 20774 19281
rect 20718 19207 20774 19216
rect 20720 19168 20772 19174
rect 20534 19136 20590 19145
rect 20720 19110 20772 19116
rect 20534 19071 20590 19080
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20364 18222 20392 18294
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20444 18148 20496 18154
rect 20444 18090 20496 18096
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20364 16658 20392 17614
rect 20456 17338 20484 18090
rect 20444 17332 20496 17338
rect 20444 17274 20496 17280
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20364 16182 20392 16594
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20364 15706 20392 15914
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20352 15564 20404 15570
rect 20352 15506 20404 15512
rect 20364 13938 20392 15506
rect 20442 13968 20498 13977
rect 20352 13932 20404 13938
rect 20442 13903 20498 13912
rect 20352 13874 20404 13880
rect 20456 13870 20484 13903
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20364 12442 20392 13670
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20456 12850 20484 13262
rect 20548 12986 20576 19071
rect 20732 18329 20760 19110
rect 20824 18834 20852 19858
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20916 19310 20944 19790
rect 21008 19786 21036 20266
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 20996 19780 21048 19786
rect 20996 19722 21048 19728
rect 21100 19666 21128 19858
rect 21546 19816 21602 19825
rect 21546 19751 21548 19760
rect 21600 19751 21602 19760
rect 21548 19722 21600 19728
rect 21928 19718 21956 22200
rect 21008 19638 21128 19666
rect 21916 19712 21968 19718
rect 21916 19654 21968 19660
rect 20904 19304 20956 19310
rect 20904 19246 20956 19252
rect 21008 19174 21036 19638
rect 21546 19408 21602 19417
rect 21546 19343 21602 19352
rect 21560 19310 21588 19343
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21548 19304 21600 19310
rect 21548 19246 21600 19252
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20812 18828 20864 18834
rect 20812 18770 20864 18776
rect 21100 18630 21128 19246
rect 21272 19236 21324 19242
rect 21272 19178 21324 19184
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20718 18320 20774 18329
rect 20718 18255 20774 18264
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20640 17610 20668 18158
rect 21100 17814 21128 18566
rect 21180 18148 21232 18154
rect 21180 18090 21232 18096
rect 21192 18057 21220 18090
rect 21178 18048 21234 18057
rect 21178 17983 21234 17992
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20916 16810 20944 17682
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 21008 17134 21036 17478
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20824 16782 20944 16810
rect 20732 16250 20760 16730
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20640 14618 20668 15506
rect 20824 15094 20852 16782
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20916 15706 20944 16594
rect 21008 16590 21036 16934
rect 21100 16794 21128 17614
rect 21178 17096 21234 17105
rect 21178 17031 21180 17040
rect 21232 17031 21234 17040
rect 21180 17002 21232 17008
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 21008 16114 21036 16526
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21100 15994 21128 16730
rect 21008 15966 21128 15994
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20628 14612 20680 14618
rect 21008 14600 21036 15966
rect 21088 15904 21140 15910
rect 21088 15846 21140 15852
rect 20628 14554 20680 14560
rect 20824 14572 21036 14600
rect 20628 14340 20680 14346
rect 20628 14282 20680 14288
rect 20640 13734 20668 14282
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 20732 13802 20760 14214
rect 20720 13796 20772 13802
rect 20720 13738 20772 13744
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20640 13297 20668 13466
rect 20626 13288 20682 13297
rect 20626 13223 20682 13232
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20628 12912 20680 12918
rect 20680 12872 20760 12900
rect 20628 12854 20680 12860
rect 20444 12844 20496 12850
rect 20496 12804 20576 12832
rect 20444 12786 20496 12792
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20364 12102 20392 12242
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20456 11914 20484 12650
rect 20548 12170 20576 12804
rect 20732 12374 20760 12872
rect 20824 12646 20852 14572
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20916 12850 20944 13330
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20720 12368 20772 12374
rect 20720 12310 20772 12316
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20364 11886 20484 11914
rect 20364 11218 20392 11886
rect 20536 11280 20588 11286
rect 20536 11222 20588 11228
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20364 8974 20392 11154
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20456 9450 20484 9998
rect 20548 9926 20576 11222
rect 20640 10606 20668 12310
rect 21008 11898 21036 14418
rect 21100 13258 21128 15846
rect 21178 15192 21234 15201
rect 21178 15127 21234 15136
rect 21192 15094 21220 15127
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 21284 14618 21312 19178
rect 22296 19174 22324 22200
rect 22756 20534 22784 22200
rect 22744 20528 22796 20534
rect 22744 20470 22796 20476
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 21546 18864 21602 18873
rect 21364 18828 21416 18834
rect 21546 18799 21548 18808
rect 21364 18770 21416 18776
rect 21600 18799 21602 18808
rect 21548 18770 21600 18776
rect 21376 18426 21404 18770
rect 21546 18456 21602 18465
rect 21364 18420 21416 18426
rect 21546 18391 21602 18400
rect 21364 18362 21416 18368
rect 21560 18358 21588 18391
rect 21548 18352 21600 18358
rect 21548 18294 21600 18300
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21560 17513 21588 17546
rect 21546 17504 21602 17513
rect 21546 17439 21602 17448
rect 21364 17060 21416 17066
rect 21364 17002 21416 17008
rect 21376 15162 21404 17002
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21468 16561 21496 16934
rect 21548 16652 21600 16658
rect 21548 16594 21600 16600
rect 21454 16552 21510 16561
rect 21454 16487 21510 16496
rect 21560 16153 21588 16594
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 21546 16144 21602 16153
rect 21546 16079 21602 16088
rect 21546 15600 21602 15609
rect 21546 15535 21548 15544
rect 21600 15535 21602 15544
rect 21548 15506 21600 15512
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21364 15156 21416 15162
rect 21364 15098 21416 15104
rect 21364 14884 21416 14890
rect 21364 14826 21416 14832
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21272 14476 21324 14482
rect 21272 14418 21324 14424
rect 21180 14340 21232 14346
rect 21180 14282 21232 14288
rect 21192 14249 21220 14282
rect 21178 14240 21234 14249
rect 21178 14175 21234 14184
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 21192 12434 21220 13874
rect 21100 12406 21220 12434
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20904 11824 20956 11830
rect 20904 11766 20956 11772
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20732 10674 20760 11086
rect 20916 11082 20944 11766
rect 20996 11688 21048 11694
rect 20996 11630 21048 11636
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 21008 10810 21036 11630
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21100 10690 21128 12406
rect 21180 12300 21232 12306
rect 21180 12242 21232 12248
rect 21192 11393 21220 12242
rect 21178 11384 21234 11393
rect 21178 11319 21234 11328
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 21008 10662 21128 10690
rect 21180 10736 21232 10742
rect 21180 10678 21232 10684
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20904 10600 20956 10606
rect 20904 10542 20956 10548
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20548 9489 20576 9862
rect 20534 9480 20590 9489
rect 20444 9444 20496 9450
rect 20534 9415 20590 9424
rect 20444 9386 20496 9392
rect 20352 8968 20404 8974
rect 20352 8910 20404 8916
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 20364 8022 20392 8434
rect 20076 8016 20128 8022
rect 20076 7958 20128 7964
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 20456 7886 20484 9386
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 9178 20576 9318
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20640 9058 20668 10542
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20824 9722 20852 10066
rect 20916 9994 20944 10542
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20548 9030 20668 9058
rect 20548 8294 20576 9030
rect 20732 8974 20760 9522
rect 20810 9480 20866 9489
rect 20810 9415 20866 9424
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20732 8786 20760 8910
rect 20640 8758 20760 8786
rect 20640 8498 20668 8758
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20824 8378 20852 9415
rect 20904 8900 20956 8906
rect 20904 8842 20956 8848
rect 20640 8350 20852 8378
rect 20536 8288 20588 8294
rect 20536 8230 20588 8236
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20548 7698 20576 8230
rect 20456 7670 20576 7698
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20180 5574 20208 5714
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20180 4622 20208 5510
rect 20168 4616 20220 4622
rect 20168 4558 20220 4564
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 20456 3194 20484 7670
rect 20640 7562 20668 8350
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20548 7534 20668 7562
rect 20824 7546 20852 7890
rect 20812 7540 20864 7546
rect 20444 3188 20496 3194
rect 20444 3130 20496 3136
rect 20548 3074 20576 7534
rect 20812 7482 20864 7488
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20732 6866 20760 7142
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20732 5642 20760 6802
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20916 5302 20944 8842
rect 21008 8634 21036 10662
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 21100 9178 21128 9590
rect 21192 9518 21220 10678
rect 21284 10266 21312 14418
rect 21376 13530 21404 14826
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21468 13410 21496 15438
rect 21548 14884 21600 14890
rect 21548 14826 21600 14832
rect 21560 14657 21588 14826
rect 21546 14648 21602 14657
rect 21546 14583 21602 14592
rect 21548 14340 21600 14346
rect 21548 14282 21600 14288
rect 21560 13841 21588 14282
rect 21546 13832 21602 13841
rect 21546 13767 21602 13776
rect 21376 13382 21496 13410
rect 21548 13388 21600 13394
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21376 9654 21404 13382
rect 21548 13330 21600 13336
rect 21560 13297 21588 13330
rect 21546 13288 21602 13297
rect 21546 13223 21602 13232
rect 21560 13190 21588 13223
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21454 12880 21510 12889
rect 21454 12815 21510 12824
rect 21468 12782 21496 12815
rect 21456 12776 21508 12782
rect 21456 12718 21508 12724
rect 21638 12472 21694 12481
rect 21638 12407 21694 12416
rect 21454 12336 21510 12345
rect 21454 12271 21456 12280
rect 21508 12271 21510 12280
rect 21456 12242 21508 12248
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21468 11937 21496 12038
rect 21454 11928 21510 11937
rect 21454 11863 21510 11872
rect 21468 11694 21496 11863
rect 21456 11688 21508 11694
rect 21456 11630 21508 11636
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21468 10538 21496 11494
rect 21560 11218 21588 11562
rect 21652 11370 21680 12407
rect 21744 11898 21772 16390
rect 21824 15360 21876 15366
rect 21824 15302 21876 15308
rect 21732 11892 21784 11898
rect 21732 11834 21784 11840
rect 21652 11342 21772 11370
rect 21640 11280 21692 11286
rect 21640 11222 21692 11228
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21560 10985 21588 11154
rect 21546 10976 21602 10985
rect 21546 10911 21602 10920
rect 21456 10532 21508 10538
rect 21456 10474 21508 10480
rect 21468 10441 21496 10474
rect 21454 10432 21510 10441
rect 21454 10367 21510 10376
rect 21652 10169 21680 11222
rect 21638 10160 21694 10169
rect 21456 10124 21508 10130
rect 21638 10095 21694 10104
rect 21456 10066 21508 10072
rect 21468 10033 21496 10066
rect 21454 10024 21510 10033
rect 21454 9959 21510 9968
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21364 9648 21416 9654
rect 21364 9590 21416 9596
rect 21560 9518 21588 9930
rect 21180 9512 21232 9518
rect 21548 9512 21600 9518
rect 21180 9454 21232 9460
rect 21546 9480 21548 9489
rect 21600 9480 21602 9489
rect 21546 9415 21602 9424
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21454 9072 21510 9081
rect 21454 9007 21456 9016
rect 21508 9007 21510 9016
rect 21456 8978 21508 8984
rect 21086 8664 21142 8673
rect 20996 8628 21048 8634
rect 21086 8599 21142 8608
rect 20996 8570 21048 8576
rect 21100 8362 21128 8599
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 21456 8356 21508 8362
rect 21456 8298 21508 8304
rect 21468 8129 21496 8298
rect 21454 8120 21510 8129
rect 21454 8055 21510 8064
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21088 7744 21140 7750
rect 21192 7721 21220 7890
rect 21088 7686 21140 7692
rect 21178 7712 21234 7721
rect 20996 7336 21048 7342
rect 20996 7278 21048 7284
rect 21008 7002 21036 7278
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 21100 6390 21128 7686
rect 21178 7647 21234 7656
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21272 7200 21324 7206
rect 21468 7177 21496 7890
rect 21272 7142 21324 7148
rect 21454 7168 21510 7177
rect 21088 6384 21140 6390
rect 21088 6326 21140 6332
rect 21192 6322 21220 7142
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 21284 5914 21312 7142
rect 21454 7103 21510 7112
rect 21456 6860 21508 6866
rect 21456 6802 21508 6808
rect 21468 6769 21496 6802
rect 21454 6760 21510 6769
rect 21454 6695 21510 6704
rect 21454 6216 21510 6225
rect 21454 6151 21456 6160
rect 21508 6151 21510 6160
rect 21456 6122 21508 6128
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 21546 5808 21602 5817
rect 21546 5743 21548 5752
rect 21600 5743 21602 5752
rect 21548 5714 21600 5720
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 20904 5296 20956 5302
rect 20904 5238 20956 5244
rect 21270 4856 21326 4865
rect 21376 4826 21404 5646
rect 21454 5264 21510 5273
rect 21454 5199 21510 5208
rect 21468 5166 21496 5199
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21270 4791 21326 4800
rect 21364 4820 21416 4826
rect 21284 4690 21312 4791
rect 21364 4762 21416 4768
rect 21272 4684 21324 4690
rect 21272 4626 21324 4632
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 21560 4457 21588 4626
rect 21546 4448 21602 4457
rect 21546 4383 21602 4392
rect 21548 4072 21600 4078
rect 21548 4014 21600 4020
rect 21560 3913 21588 4014
rect 21546 3904 21602 3913
rect 21546 3839 21602 3848
rect 21652 3738 21680 10095
rect 21744 8634 21772 11342
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21836 8090 21864 15302
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 21548 3596 21600 3602
rect 21548 3538 21600 3544
rect 21456 3528 21508 3534
rect 21560 3505 21588 3538
rect 21456 3470 21508 3476
rect 21546 3496 21602 3505
rect 20996 3460 21048 3466
rect 20996 3402 21048 3408
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20456 3046 20576 3074
rect 20640 3058 20668 3334
rect 21008 3194 21036 3402
rect 20996 3188 21048 3194
rect 20996 3130 21048 3136
rect 20628 3052 20680 3058
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 17960 2576 18012 2582
rect 17960 2518 18012 2524
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 6920 2372 6972 2378
rect 6920 2314 6972 2320
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4160 2100 4212 2106
rect 4160 2042 4212 2048
rect 3514 2000 3570 2009
rect 3514 1935 3570 1944
rect 6932 800 6960 2314
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11716 1578 11744 2450
rect 16132 2310 16160 2450
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 11532 1550 11744 1578
rect 11532 800 11560 1550
rect 16132 800 16160 2246
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 20364 1601 20392 2450
rect 20456 2310 20484 3046
rect 20628 2994 20680 3000
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 20444 2304 20496 2310
rect 20444 2246 20496 2252
rect 20548 2009 20576 2926
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 20640 2514 20668 2858
rect 20628 2508 20680 2514
rect 20628 2450 20680 2456
rect 20720 2508 20772 2514
rect 20824 2496 20852 2926
rect 20772 2468 20852 2496
rect 21178 2544 21234 2553
rect 21178 2479 21180 2488
rect 20720 2450 20772 2456
rect 21232 2479 21234 2488
rect 21180 2450 21232 2456
rect 20534 2000 20590 2009
rect 20534 1935 20590 1944
rect 20350 1592 20406 1601
rect 20350 1527 20406 1536
rect 20640 1057 20668 2450
rect 20626 1048 20682 1057
rect 20626 983 20682 992
rect 20732 800 20760 2450
rect 2870 232 2926 241
rect 2870 167 2926 176
rect 6918 0 6974 800
rect 11518 0 11574 800
rect 16118 0 16174 800
rect 20718 0 20774 800
rect 21284 241 21312 2926
rect 21468 2514 21496 3470
rect 21546 3431 21602 3440
rect 21548 3392 21600 3398
rect 21548 3334 21600 3340
rect 21560 2990 21588 3334
rect 21548 2984 21600 2990
rect 21546 2952 21548 2961
rect 21600 2952 21602 2961
rect 21546 2887 21602 2896
rect 21928 2650 21956 11018
rect 21916 2644 21968 2650
rect 21916 2586 21968 2592
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 21468 649 21496 2450
rect 21454 640 21510 649
rect 21454 575 21510 584
rect 21270 232 21326 241
rect 21270 167 21326 176
<< via2 >>
rect 3330 22208 3386 22264
rect 1858 20712 1914 20768
rect 2134 20324 2190 20360
rect 2134 20304 2136 20324
rect 2136 20304 2188 20324
rect 2188 20304 2190 20324
rect 1398 19780 1454 19816
rect 1398 19760 1400 19780
rect 1400 19760 1452 19780
rect 1452 19760 1454 19780
rect 1398 19352 1454 19408
rect 2962 21664 3018 21720
rect 2778 21256 2834 21312
rect 2594 20460 2650 20496
rect 2594 20440 2596 20460
rect 2596 20440 2648 20460
rect 2648 20440 2650 20460
rect 2778 20460 2834 20496
rect 2778 20440 2780 20460
rect 2780 20440 2832 20460
rect 2832 20440 2834 20460
rect 2502 20324 2558 20360
rect 2502 20304 2504 20324
rect 2504 20304 2556 20324
rect 2556 20304 2558 20324
rect 2594 19780 2650 19816
rect 2594 19760 2596 19780
rect 2596 19760 2648 19780
rect 2648 19760 2650 19780
rect 1398 18828 1454 18864
rect 1398 18808 1400 18828
rect 1400 18808 1452 18828
rect 1452 18808 1454 18828
rect 1490 18420 1546 18456
rect 1490 18400 1492 18420
rect 1492 18400 1544 18420
rect 1544 18400 1546 18420
rect 1490 17484 1492 17504
rect 1492 17484 1544 17504
rect 1544 17484 1546 17504
rect 1490 17448 1546 17484
rect 1398 17060 1454 17096
rect 1398 17040 1400 17060
rect 1400 17040 1452 17060
rect 1452 17040 1454 17060
rect 1398 16496 1454 16552
rect 1398 16108 1454 16144
rect 1398 16088 1400 16108
rect 1400 16088 1452 16108
rect 1452 16088 1454 16108
rect 1398 15564 1454 15600
rect 1398 15544 1400 15564
rect 1400 15544 1452 15564
rect 1452 15544 1454 15564
rect 1490 15156 1546 15192
rect 1490 15136 1492 15156
rect 1492 15136 1544 15156
rect 1544 15136 1546 15156
rect 1490 14220 1492 14240
rect 1492 14220 1544 14240
rect 1544 14220 1546 14240
rect 1490 14184 1546 14220
rect 1306 13640 1362 13696
rect 1398 13232 1454 13288
rect 1306 12824 1362 12880
rect 1490 12144 1546 12200
rect 1490 10920 1546 10976
rect 1398 10376 1454 10432
rect 1950 19216 2006 19272
rect 1858 18028 1860 18048
rect 1860 18028 1912 18048
rect 1912 18028 1914 18048
rect 1858 17992 1914 18028
rect 2226 18692 2282 18728
rect 2226 18672 2228 18692
rect 2228 18672 2280 18692
rect 2280 18672 2282 18692
rect 2502 18808 2558 18864
rect 2962 19624 3018 19680
rect 2870 18964 2926 19000
rect 2870 18944 2872 18964
rect 2872 18944 2924 18964
rect 2924 18944 2926 18964
rect 1858 14612 1914 14648
rect 1858 14592 1860 14612
rect 1860 14592 1912 14612
rect 1912 14592 1914 14612
rect 1766 13812 1768 13832
rect 1768 13812 1820 13832
rect 1820 13812 1822 13832
rect 1766 13776 1822 13812
rect 1950 12844 2006 12880
rect 1950 12824 1952 12844
rect 1952 12824 2004 12844
rect 2004 12824 2006 12844
rect 1858 12280 1914 12336
rect 1766 11328 1822 11384
rect 1674 10532 1730 10568
rect 1674 10512 1676 10532
rect 1676 10512 1728 10532
rect 1728 10512 1730 10532
rect 1490 9968 1546 10024
rect 1490 9016 1546 9072
rect 1398 8064 1454 8120
rect 1398 7112 1454 7168
rect 3882 22616 3938 22672
rect 3238 20304 3294 20360
rect 3146 18264 3202 18320
rect 3422 19916 3478 19952
rect 3422 19896 3424 19916
rect 3424 19896 3476 19916
rect 3476 19896 3478 19916
rect 18970 22616 19026 22672
rect 2686 13640 2742 13696
rect 2962 12824 3018 12880
rect 2042 9424 2098 9480
rect 1858 8608 1914 8664
rect 1766 7656 1822 7712
rect 1490 6704 1546 6760
rect 1490 6180 1546 6216
rect 1490 6160 1492 6180
rect 1492 6160 1544 6180
rect 1544 6160 1546 6180
rect 1398 5772 1454 5808
rect 1398 5752 1400 5772
rect 1400 5752 1452 5772
rect 1452 5752 1454 5772
rect 1490 5208 1546 5264
rect 1674 4800 1730 4856
rect 1398 4392 1454 4448
rect 1398 3848 1454 3904
rect 1398 3440 1454 3496
rect 1398 2932 1400 2952
rect 1400 2932 1452 2952
rect 1452 2932 1454 2952
rect 1398 2896 1454 2932
rect 1398 2508 1454 2544
rect 1398 2488 1400 2508
rect 1400 2488 1452 2508
rect 1452 2488 1454 2508
rect 2870 8880 2926 8936
rect 2778 8064 2834 8120
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4158 19896 4214 19952
rect 4250 19624 4306 19680
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4066 17604 4122 17640
rect 4066 17584 4068 17604
rect 4068 17584 4120 17604
rect 4120 17584 4122 17604
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 1950 1536 2006 1592
rect 1674 992 1730 1048
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 3974 12180 3976 12200
rect 3976 12180 4028 12200
rect 4028 12180 4030 12200
rect 3974 12144 4030 12180
rect 4710 12180 4712 12200
rect 4712 12180 4764 12200
rect 4764 12180 4766 12200
rect 4710 12144 4766 12180
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4894 12008 4950 12064
rect 5722 12688 5778 12744
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4526 9580 4582 9616
rect 4526 9560 4528 9580
rect 4528 9560 4580 9580
rect 4580 9560 4582 9580
rect 4342 9288 4398 9344
rect 2778 584 2834 640
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4894 8472 4950 8528
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 5262 11464 5318 11520
rect 5722 9560 5778 9616
rect 5262 7384 5318 7440
rect 5446 8472 5502 8528
rect 6458 12180 6460 12200
rect 6460 12180 6512 12200
rect 6512 12180 6514 12200
rect 6458 12144 6514 12180
rect 5446 6976 5502 7032
rect 7102 17856 7158 17912
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7654 18944 7710 19000
rect 7286 18164 7288 18184
rect 7288 18164 7340 18184
rect 7340 18164 7342 18184
rect 7286 18128 7342 18164
rect 7470 17720 7526 17776
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7930 18284 7986 18320
rect 7930 18264 7932 18284
rect 7932 18264 7984 18284
rect 7984 18264 7986 18284
rect 8390 18128 8446 18184
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 8206 15000 8262 15056
rect 7654 14864 7710 14920
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7010 8880 7066 8936
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7562 9324 7564 9344
rect 7564 9324 7616 9344
rect 7616 9324 7618 9344
rect 7562 9288 7618 9324
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7654 8064 7710 8120
rect 9218 13776 9274 13832
rect 9586 17992 9642 18048
rect 9954 17312 10010 17368
rect 9954 16496 10010 16552
rect 9770 14900 9772 14920
rect 9772 14900 9824 14920
rect 9824 14900 9826 14920
rect 9770 14864 9826 14900
rect 9678 14340 9734 14376
rect 9678 14320 9680 14340
rect 9680 14320 9732 14340
rect 9732 14320 9734 14340
rect 9586 13912 9642 13968
rect 9126 10648 9182 10704
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 10138 18264 10194 18320
rect 10138 16496 10194 16552
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 10690 17312 10746 17368
rect 10598 16532 10600 16552
rect 10600 16532 10652 16552
rect 10652 16532 10654 16552
rect 10598 16496 10654 16532
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11610 17604 11666 17640
rect 11610 17584 11612 17604
rect 11612 17584 11664 17604
rect 11664 17584 11666 17604
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 10874 12824 10930 12880
rect 10506 11192 10562 11248
rect 9862 8880 9918 8936
rect 11058 11600 11114 11656
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 10782 8880 10838 8936
rect 11334 8916 11336 8936
rect 11336 8916 11388 8936
rect 11388 8916 11390 8936
rect 11334 8880 11390 8916
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11978 15020 12034 15056
rect 12254 18128 12310 18184
rect 11978 15000 11980 15020
rect 11980 15000 12032 15020
rect 12032 15000 12034 15020
rect 12530 18300 12532 18320
rect 12532 18300 12584 18320
rect 12584 18300 12586 18320
rect 12530 18264 12586 18300
rect 12438 18128 12494 18184
rect 12622 14320 12678 14376
rect 13450 18264 13506 18320
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 14830 19624 14886 19680
rect 15382 19624 15438 19680
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14646 18264 14702 18320
rect 12346 10548 12348 10568
rect 12348 10548 12400 10568
rect 12400 10548 12402 10568
rect 12346 10512 12402 10548
rect 12990 10512 13046 10568
rect 13726 12688 13782 12744
rect 14186 12552 14242 12608
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 15474 16496 15530 16552
rect 16670 20032 16726 20088
rect 16210 18808 16266 18864
rect 16762 19760 16818 19816
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 16762 18672 16818 18728
rect 16670 18400 16726 18456
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 14830 12688 14886 12744
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 15106 11736 15162 11792
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 15106 9832 15162 9888
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 19798 22208 19854 22264
rect 19706 21664 19762 21720
rect 19062 20032 19118 20088
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18510 18944 18566 19000
rect 18050 18536 18106 18592
rect 18418 18672 18474 18728
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18694 19216 18750 19272
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18878 19116 18880 19136
rect 18880 19116 18932 19136
rect 18932 19116 18934 19136
rect 18878 19080 18934 19116
rect 19246 19080 19302 19136
rect 19614 19116 19616 19136
rect 19616 19116 19668 19136
rect 19668 19116 19670 19136
rect 19614 19080 19670 19116
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 15382 11600 15438 11656
rect 17866 12824 17922 12880
rect 20442 21256 20498 21312
rect 20534 20712 20590 20768
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18326 12860 18328 12880
rect 18328 12860 18380 12880
rect 18380 12860 18382 12880
rect 18326 12824 18382 12860
rect 17958 11736 18014 11792
rect 17774 11600 17830 11656
rect 18694 12416 18750 12472
rect 17958 11212 18014 11248
rect 17958 11192 17960 11212
rect 17960 11192 18012 11212
rect 18012 11192 18014 11212
rect 16670 9968 16726 10024
rect 17222 9832 17278 9888
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18510 11464 18566 11520
rect 18878 12144 18934 12200
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 19154 12280 19210 12336
rect 19338 13912 19394 13968
rect 19430 12688 19486 12744
rect 19062 10648 19118 10704
rect 19338 10140 19340 10160
rect 19340 10140 19392 10160
rect 19392 10140 19394 10160
rect 19338 10104 19394 10140
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18602 8900 18658 8936
rect 18602 8880 18604 8900
rect 18604 8880 18656 8900
rect 18656 8880 18658 8900
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 19614 13252 19670 13288
rect 19614 13232 19616 13252
rect 19616 13232 19668 13252
rect 19668 13232 19670 13252
rect 19522 11736 19578 11792
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 19982 12316 19984 12336
rect 19984 12316 20036 12336
rect 20036 12316 20038 12336
rect 19982 12280 20038 12316
rect 20074 11500 20076 11520
rect 20076 11500 20128 11520
rect 20128 11500 20130 11520
rect 20074 11464 20130 11500
rect 19982 8472 20038 8528
rect 21178 20324 21234 20360
rect 21178 20304 21180 20324
rect 21180 20304 21232 20324
rect 21232 20304 21234 20324
rect 20718 19216 20774 19272
rect 20534 19080 20590 19136
rect 20442 13912 20498 13968
rect 21546 19780 21602 19816
rect 21546 19760 21548 19780
rect 21548 19760 21600 19780
rect 21600 19760 21602 19780
rect 21546 19352 21602 19408
rect 20718 18264 20774 18320
rect 21178 17992 21234 18048
rect 21178 17060 21234 17096
rect 21178 17040 21180 17060
rect 21180 17040 21232 17060
rect 21232 17040 21234 17060
rect 20626 13232 20682 13288
rect 21178 15136 21234 15192
rect 21546 18828 21602 18864
rect 21546 18808 21548 18828
rect 21548 18808 21600 18828
rect 21600 18808 21602 18828
rect 21546 18400 21602 18456
rect 21546 17448 21602 17504
rect 21454 16496 21510 16552
rect 21546 16088 21602 16144
rect 21546 15564 21602 15600
rect 21546 15544 21548 15564
rect 21548 15544 21600 15564
rect 21600 15544 21602 15564
rect 21178 14184 21234 14240
rect 21178 11328 21234 11384
rect 20534 9424 20590 9480
rect 20810 9424 20866 9480
rect 21546 14592 21602 14648
rect 21546 13776 21602 13832
rect 21546 13232 21602 13288
rect 21454 12824 21510 12880
rect 21638 12416 21694 12472
rect 21454 12300 21510 12336
rect 21454 12280 21456 12300
rect 21456 12280 21508 12300
rect 21508 12280 21510 12300
rect 21454 11872 21510 11928
rect 21546 10920 21602 10976
rect 21454 10376 21510 10432
rect 21638 10104 21694 10160
rect 21454 9968 21510 10024
rect 21546 9460 21548 9480
rect 21548 9460 21600 9480
rect 21600 9460 21602 9480
rect 21546 9424 21602 9460
rect 21454 9036 21510 9072
rect 21454 9016 21456 9036
rect 21456 9016 21508 9036
rect 21508 9016 21510 9036
rect 21086 8608 21142 8664
rect 21454 8064 21510 8120
rect 21178 7656 21234 7712
rect 21454 7112 21510 7168
rect 21454 6704 21510 6760
rect 21454 6180 21510 6216
rect 21454 6160 21456 6180
rect 21456 6160 21508 6180
rect 21508 6160 21510 6180
rect 21546 5772 21602 5808
rect 21546 5752 21548 5772
rect 21548 5752 21600 5772
rect 21600 5752 21602 5772
rect 21270 4800 21326 4856
rect 21454 5208 21510 5264
rect 21546 4392 21602 4448
rect 21546 3848 21602 3904
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 3514 1944 3570 2000
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 21178 2508 21234 2544
rect 21178 2488 21180 2508
rect 21180 2488 21232 2508
rect 21232 2488 21234 2508
rect 20534 1944 20590 2000
rect 20350 1536 20406 1592
rect 20626 992 20682 1048
rect 2870 176 2926 232
rect 21546 3440 21602 3496
rect 21546 2932 21548 2952
rect 21548 2932 21600 2952
rect 21600 2932 21602 2952
rect 21546 2896 21602 2932
rect 21454 584 21510 640
rect 21270 176 21326 232
<< metal3 >>
rect 0 22674 800 22704
rect 3877 22674 3943 22677
rect 0 22672 3943 22674
rect 0 22616 3882 22672
rect 3938 22616 3943 22672
rect 0 22614 3943 22616
rect 0 22584 800 22614
rect 3877 22611 3943 22614
rect 18965 22674 19031 22677
rect 22200 22674 23000 22704
rect 18965 22672 23000 22674
rect 18965 22616 18970 22672
rect 19026 22616 23000 22672
rect 18965 22614 23000 22616
rect 18965 22611 19031 22614
rect 22200 22584 23000 22614
rect 0 22266 800 22296
rect 3325 22266 3391 22269
rect 0 22264 3391 22266
rect 0 22208 3330 22264
rect 3386 22208 3391 22264
rect 0 22206 3391 22208
rect 0 22176 800 22206
rect 3325 22203 3391 22206
rect 19793 22266 19859 22269
rect 22200 22266 23000 22296
rect 19793 22264 23000 22266
rect 19793 22208 19798 22264
rect 19854 22208 23000 22264
rect 19793 22206 23000 22208
rect 19793 22203 19859 22206
rect 22200 22176 23000 22206
rect 0 21722 800 21752
rect 2957 21722 3023 21725
rect 0 21720 3023 21722
rect 0 21664 2962 21720
rect 3018 21664 3023 21720
rect 0 21662 3023 21664
rect 0 21632 800 21662
rect 2957 21659 3023 21662
rect 19701 21722 19767 21725
rect 22200 21722 23000 21752
rect 19701 21720 23000 21722
rect 19701 21664 19706 21720
rect 19762 21664 23000 21720
rect 19701 21662 23000 21664
rect 19701 21659 19767 21662
rect 22200 21632 23000 21662
rect 0 21314 800 21344
rect 2773 21314 2839 21317
rect 0 21312 2839 21314
rect 0 21256 2778 21312
rect 2834 21256 2839 21312
rect 0 21254 2839 21256
rect 0 21224 800 21254
rect 2773 21251 2839 21254
rect 20437 21314 20503 21317
rect 22200 21314 23000 21344
rect 20437 21312 23000 21314
rect 20437 21256 20442 21312
rect 20498 21256 23000 21312
rect 20437 21254 23000 21256
rect 20437 21251 20503 21254
rect 22200 21224 23000 21254
rect 0 20770 800 20800
rect 1853 20770 1919 20773
rect 0 20768 1919 20770
rect 0 20712 1858 20768
rect 1914 20712 1919 20768
rect 0 20710 1919 20712
rect 0 20680 800 20710
rect 1853 20707 1919 20710
rect 20529 20770 20595 20773
rect 22200 20770 23000 20800
rect 20529 20768 23000 20770
rect 20529 20712 20534 20768
rect 20590 20712 23000 20768
rect 20529 20710 23000 20712
rect 20529 20707 20595 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 22200 20680 23000 20710
rect 18270 20639 18590 20640
rect 2589 20498 2655 20501
rect 2773 20498 2839 20501
rect 2589 20496 2839 20498
rect 2589 20440 2594 20496
rect 2650 20440 2778 20496
rect 2834 20440 2839 20496
rect 2589 20438 2839 20440
rect 2589 20435 2655 20438
rect 2773 20435 2839 20438
rect 0 20362 800 20392
rect 2129 20362 2195 20365
rect 0 20360 2195 20362
rect 0 20304 2134 20360
rect 2190 20304 2195 20360
rect 0 20302 2195 20304
rect 0 20272 800 20302
rect 2129 20299 2195 20302
rect 2497 20362 2563 20365
rect 3233 20362 3299 20365
rect 2497 20360 3299 20362
rect 2497 20304 2502 20360
rect 2558 20304 3238 20360
rect 3294 20304 3299 20360
rect 2497 20302 3299 20304
rect 2497 20299 2563 20302
rect 3233 20299 3299 20302
rect 21173 20362 21239 20365
rect 22200 20362 23000 20392
rect 21173 20360 23000 20362
rect 21173 20304 21178 20360
rect 21234 20304 23000 20360
rect 21173 20302 23000 20304
rect 21173 20299 21239 20302
rect 22200 20272 23000 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 16665 20090 16731 20093
rect 19057 20090 19123 20093
rect 16665 20088 19123 20090
rect 16665 20032 16670 20088
rect 16726 20032 19062 20088
rect 19118 20032 19123 20088
rect 16665 20030 19123 20032
rect 16665 20027 16731 20030
rect 19057 20027 19123 20030
rect 3417 19954 3483 19957
rect 4153 19954 4219 19957
rect 3417 19952 4219 19954
rect 3417 19896 3422 19952
rect 3478 19896 4158 19952
rect 4214 19896 4219 19952
rect 3417 19894 4219 19896
rect 3417 19891 3483 19894
rect 4153 19891 4219 19894
rect 0 19818 800 19848
rect 1393 19818 1459 19821
rect 0 19816 1459 19818
rect 0 19760 1398 19816
rect 1454 19760 1459 19816
rect 0 19758 1459 19760
rect 0 19728 800 19758
rect 1393 19755 1459 19758
rect 2589 19818 2655 19821
rect 16757 19818 16823 19821
rect 2589 19816 16823 19818
rect 2589 19760 2594 19816
rect 2650 19760 16762 19816
rect 16818 19760 16823 19816
rect 2589 19758 16823 19760
rect 2589 19755 2655 19758
rect 16757 19755 16823 19758
rect 21541 19818 21607 19821
rect 22200 19818 23000 19848
rect 21541 19816 23000 19818
rect 21541 19760 21546 19816
rect 21602 19760 23000 19816
rect 21541 19758 23000 19760
rect 21541 19755 21607 19758
rect 22200 19728 23000 19758
rect 2957 19682 3023 19685
rect 4245 19682 4311 19685
rect 2957 19680 4311 19682
rect 2957 19624 2962 19680
rect 3018 19624 4250 19680
rect 4306 19624 4311 19680
rect 2957 19622 4311 19624
rect 2957 19619 3023 19622
rect 4245 19619 4311 19622
rect 14825 19682 14891 19685
rect 15377 19682 15443 19685
rect 14825 19680 15443 19682
rect 14825 19624 14830 19680
rect 14886 19624 15382 19680
rect 15438 19624 15443 19680
rect 14825 19622 15443 19624
rect 14825 19619 14891 19622
rect 15377 19619 15443 19622
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 0 19410 800 19440
rect 1393 19410 1459 19413
rect 0 19408 1459 19410
rect 0 19352 1398 19408
rect 1454 19352 1459 19408
rect 0 19350 1459 19352
rect 0 19320 800 19350
rect 1393 19347 1459 19350
rect 21541 19410 21607 19413
rect 22200 19410 23000 19440
rect 21541 19408 23000 19410
rect 21541 19352 21546 19408
rect 21602 19352 23000 19408
rect 21541 19350 23000 19352
rect 21541 19347 21607 19350
rect 22200 19320 23000 19350
rect 1945 19274 2011 19277
rect 18689 19274 18755 19277
rect 20713 19274 20779 19277
rect 1945 19272 20779 19274
rect 1945 19216 1950 19272
rect 2006 19216 18694 19272
rect 18750 19216 20718 19272
rect 20774 19216 20779 19272
rect 1945 19214 20779 19216
rect 1945 19211 2011 19214
rect 18689 19211 18755 19214
rect 20713 19211 20779 19214
rect 18873 19138 18939 19141
rect 19241 19138 19307 19141
rect 18873 19136 19307 19138
rect 18873 19080 18878 19136
rect 18934 19080 19246 19136
rect 19302 19080 19307 19136
rect 18873 19078 19307 19080
rect 18873 19075 18939 19078
rect 19241 19075 19307 19078
rect 19609 19138 19675 19141
rect 20529 19138 20595 19141
rect 19609 19136 20595 19138
rect 19609 19080 19614 19136
rect 19670 19080 20534 19136
rect 20590 19080 20595 19136
rect 19609 19078 20595 19080
rect 19609 19075 19675 19078
rect 20529 19075 20595 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 2865 19002 2931 19005
rect 7649 19002 7715 19005
rect 2865 19000 7715 19002
rect 2865 18944 2870 19000
rect 2926 18944 7654 19000
rect 7710 18944 7715 19000
rect 2865 18942 7715 18944
rect 2865 18939 2931 18942
rect 7649 18939 7715 18942
rect 18505 19002 18571 19005
rect 19612 19002 19672 19075
rect 18505 19000 19672 19002
rect 18505 18944 18510 19000
rect 18566 18944 19672 19000
rect 18505 18942 19672 18944
rect 18505 18939 18571 18942
rect 0 18866 800 18896
rect 1393 18866 1459 18869
rect 0 18864 1459 18866
rect 0 18808 1398 18864
rect 1454 18808 1459 18864
rect 0 18806 1459 18808
rect 0 18776 800 18806
rect 1393 18803 1459 18806
rect 2497 18866 2563 18869
rect 16205 18866 16271 18869
rect 2497 18864 16271 18866
rect 2497 18808 2502 18864
rect 2558 18808 16210 18864
rect 16266 18808 16271 18864
rect 2497 18806 16271 18808
rect 2497 18803 2563 18806
rect 16205 18803 16271 18806
rect 21541 18866 21607 18869
rect 22200 18866 23000 18896
rect 21541 18864 23000 18866
rect 21541 18808 21546 18864
rect 21602 18808 23000 18864
rect 21541 18806 23000 18808
rect 21541 18803 21607 18806
rect 22200 18776 23000 18806
rect 2221 18730 2287 18733
rect 16757 18730 16823 18733
rect 18413 18730 18479 18733
rect 2221 18728 12450 18730
rect 2221 18672 2226 18728
rect 2282 18672 12450 18728
rect 2221 18670 12450 18672
rect 2221 18667 2287 18670
rect 12390 18594 12450 18670
rect 16757 18728 18479 18730
rect 16757 18672 16762 18728
rect 16818 18672 18418 18728
rect 18474 18672 18479 18728
rect 16757 18670 18479 18672
rect 16757 18667 16823 18670
rect 18413 18667 18479 18670
rect 18045 18594 18111 18597
rect 12390 18592 18111 18594
rect 12390 18536 18050 18592
rect 18106 18536 18111 18592
rect 12390 18534 18111 18536
rect 18045 18531 18111 18534
rect 4409 18528 4729 18529
rect 0 18458 800 18488
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 1485 18458 1551 18461
rect 16665 18458 16731 18461
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 12390 18456 16731 18458
rect 12390 18400 16670 18456
rect 16726 18400 16731 18456
rect 12390 18398 16731 18400
rect 3141 18322 3207 18325
rect 7925 18322 7991 18325
rect 3141 18320 7991 18322
rect 3141 18264 3146 18320
rect 3202 18264 7930 18320
rect 7986 18264 7991 18320
rect 3141 18262 7991 18264
rect 3141 18259 3207 18262
rect 7925 18259 7991 18262
rect 10133 18322 10199 18325
rect 12390 18322 12450 18398
rect 16665 18395 16731 18398
rect 21541 18458 21607 18461
rect 22200 18458 23000 18488
rect 21541 18456 23000 18458
rect 21541 18400 21546 18456
rect 21602 18400 23000 18456
rect 21541 18398 23000 18400
rect 21541 18395 21607 18398
rect 22200 18368 23000 18398
rect 10133 18320 12450 18322
rect 10133 18264 10138 18320
rect 10194 18264 12450 18320
rect 10133 18262 12450 18264
rect 12525 18322 12591 18325
rect 13445 18322 13511 18325
rect 12525 18320 13511 18322
rect 12525 18264 12530 18320
rect 12586 18264 13450 18320
rect 13506 18264 13511 18320
rect 12525 18262 13511 18264
rect 10133 18259 10199 18262
rect 12525 18259 12591 18262
rect 13445 18259 13511 18262
rect 14641 18322 14707 18325
rect 20713 18322 20779 18325
rect 14641 18320 20779 18322
rect 14641 18264 14646 18320
rect 14702 18264 20718 18320
rect 20774 18264 20779 18320
rect 14641 18262 20779 18264
rect 14641 18259 14707 18262
rect 20713 18259 20779 18262
rect 7281 18186 7347 18189
rect 8385 18186 8451 18189
rect 7281 18184 8451 18186
rect 7281 18128 7286 18184
rect 7342 18128 8390 18184
rect 8446 18128 8451 18184
rect 7281 18126 8451 18128
rect 7281 18123 7347 18126
rect 8385 18123 8451 18126
rect 12249 18186 12315 18189
rect 12433 18186 12499 18189
rect 12249 18184 12499 18186
rect 12249 18128 12254 18184
rect 12310 18128 12438 18184
rect 12494 18128 12499 18184
rect 12249 18126 12499 18128
rect 12249 18123 12315 18126
rect 12433 18123 12499 18126
rect 0 18050 800 18080
rect 1853 18050 1919 18053
rect 0 18048 1919 18050
rect 0 17992 1858 18048
rect 1914 17992 1919 18048
rect 0 17990 1919 17992
rect 0 17960 800 17990
rect 1853 17987 1919 17990
rect 9438 17988 9444 18052
rect 9508 18050 9514 18052
rect 9581 18050 9647 18053
rect 9508 18048 9647 18050
rect 9508 17992 9586 18048
rect 9642 17992 9647 18048
rect 9508 17990 9647 17992
rect 9508 17988 9514 17990
rect 9581 17987 9647 17990
rect 21173 18050 21239 18053
rect 22200 18050 23000 18080
rect 21173 18048 23000 18050
rect 21173 17992 21178 18048
rect 21234 17992 23000 18048
rect 21173 17990 23000 17992
rect 21173 17987 21239 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 7097 17914 7163 17917
rect 7097 17912 7298 17914
rect 7097 17856 7102 17912
rect 7158 17856 7298 17912
rect 7097 17854 7298 17856
rect 7097 17851 7163 17854
rect 7238 17778 7298 17854
rect 7465 17778 7531 17781
rect 7238 17776 7531 17778
rect 7238 17720 7470 17776
rect 7526 17720 7531 17776
rect 7238 17718 7531 17720
rect 7465 17715 7531 17718
rect 4061 17642 4127 17645
rect 11605 17642 11671 17645
rect 4061 17640 11671 17642
rect 4061 17584 4066 17640
rect 4122 17584 11610 17640
rect 11666 17584 11671 17640
rect 4061 17582 11671 17584
rect 4061 17579 4127 17582
rect 11605 17579 11671 17582
rect 0 17506 800 17536
rect 1485 17506 1551 17509
rect 0 17504 1551 17506
rect 0 17448 1490 17504
rect 1546 17448 1551 17504
rect 0 17446 1551 17448
rect 0 17416 800 17446
rect 1485 17443 1551 17446
rect 21541 17506 21607 17509
rect 22200 17506 23000 17536
rect 21541 17504 23000 17506
rect 21541 17448 21546 17504
rect 21602 17448 23000 17504
rect 21541 17446 23000 17448
rect 21541 17443 21607 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 22200 17416 23000 17446
rect 18270 17375 18590 17376
rect 9949 17370 10015 17373
rect 10685 17370 10751 17373
rect 9949 17368 10751 17370
rect 9949 17312 9954 17368
rect 10010 17312 10690 17368
rect 10746 17312 10751 17368
rect 9949 17310 10751 17312
rect 9949 17307 10015 17310
rect 10685 17307 10751 17310
rect 0 17098 800 17128
rect 1393 17098 1459 17101
rect 0 17096 1459 17098
rect 0 17040 1398 17096
rect 1454 17040 1459 17096
rect 0 17038 1459 17040
rect 0 17008 800 17038
rect 1393 17035 1459 17038
rect 21173 17098 21239 17101
rect 22200 17098 23000 17128
rect 21173 17096 23000 17098
rect 21173 17040 21178 17096
rect 21234 17040 23000 17096
rect 21173 17038 23000 17040
rect 21173 17035 21239 17038
rect 22200 17008 23000 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 0 16554 800 16584
rect 1393 16554 1459 16557
rect 0 16552 1459 16554
rect 0 16496 1398 16552
rect 1454 16496 1459 16552
rect 0 16494 1459 16496
rect 0 16464 800 16494
rect 1393 16491 1459 16494
rect 9949 16554 10015 16557
rect 10133 16554 10199 16557
rect 9949 16552 10199 16554
rect 9949 16496 9954 16552
rect 10010 16496 10138 16552
rect 10194 16496 10199 16552
rect 9949 16494 10199 16496
rect 9949 16491 10015 16494
rect 10133 16491 10199 16494
rect 10593 16554 10659 16557
rect 15469 16554 15535 16557
rect 10593 16552 15535 16554
rect 10593 16496 10598 16552
rect 10654 16496 15474 16552
rect 15530 16496 15535 16552
rect 10593 16494 15535 16496
rect 10593 16491 10659 16494
rect 15469 16491 15535 16494
rect 21449 16554 21515 16557
rect 22200 16554 23000 16584
rect 21449 16552 23000 16554
rect 21449 16496 21454 16552
rect 21510 16496 23000 16552
rect 21449 16494 23000 16496
rect 21449 16491 21515 16494
rect 22200 16464 23000 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 800 16176
rect 1393 16146 1459 16149
rect 0 16144 1459 16146
rect 0 16088 1398 16144
rect 1454 16088 1459 16144
rect 0 16086 1459 16088
rect 0 16056 800 16086
rect 1393 16083 1459 16086
rect 21541 16146 21607 16149
rect 22200 16146 23000 16176
rect 21541 16144 23000 16146
rect 21541 16088 21546 16144
rect 21602 16088 23000 16144
rect 21541 16086 23000 16088
rect 21541 16083 21607 16086
rect 22200 16056 23000 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15602 800 15632
rect 1393 15602 1459 15605
rect 0 15600 1459 15602
rect 0 15544 1398 15600
rect 1454 15544 1459 15600
rect 0 15542 1459 15544
rect 0 15512 800 15542
rect 1393 15539 1459 15542
rect 21541 15602 21607 15605
rect 22200 15602 23000 15632
rect 21541 15600 23000 15602
rect 21541 15544 21546 15600
rect 21602 15544 23000 15600
rect 21541 15542 23000 15544
rect 21541 15539 21607 15542
rect 22200 15512 23000 15542
rect 4409 15264 4729 15265
rect 0 15194 800 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 21173 15194 21239 15197
rect 22200 15194 23000 15224
rect 21173 15192 23000 15194
rect 21173 15136 21178 15192
rect 21234 15136 23000 15192
rect 21173 15134 23000 15136
rect 21173 15131 21239 15134
rect 22200 15104 23000 15134
rect 8201 15058 8267 15061
rect 11973 15058 12039 15061
rect 8201 15056 12039 15058
rect 8201 15000 8206 15056
rect 8262 15000 11978 15056
rect 12034 15000 12039 15056
rect 8201 14998 12039 15000
rect 8201 14995 8267 14998
rect 11973 14995 12039 14998
rect 7649 14922 7715 14925
rect 9765 14922 9831 14925
rect 7649 14920 9831 14922
rect 7649 14864 7654 14920
rect 7710 14864 9770 14920
rect 9826 14864 9831 14920
rect 7649 14862 9831 14864
rect 7649 14859 7715 14862
rect 9765 14859 9831 14862
rect 7874 14720 8194 14721
rect 0 14650 800 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 1853 14650 1919 14653
rect 0 14648 1919 14650
rect 0 14592 1858 14648
rect 1914 14592 1919 14648
rect 0 14590 1919 14592
rect 0 14560 800 14590
rect 1853 14587 1919 14590
rect 21541 14650 21607 14653
rect 22200 14650 23000 14680
rect 21541 14648 23000 14650
rect 21541 14592 21546 14648
rect 21602 14592 23000 14648
rect 21541 14590 23000 14592
rect 21541 14587 21607 14590
rect 22200 14560 23000 14590
rect 9673 14378 9739 14381
rect 12617 14378 12683 14381
rect 9673 14376 12683 14378
rect 9673 14320 9678 14376
rect 9734 14320 12622 14376
rect 12678 14320 12683 14376
rect 9673 14318 12683 14320
rect 9673 14315 9739 14318
rect 12617 14315 12683 14318
rect 0 14242 800 14272
rect 1485 14242 1551 14245
rect 0 14240 1551 14242
rect 0 14184 1490 14240
rect 1546 14184 1551 14240
rect 0 14182 1551 14184
rect 0 14152 800 14182
rect 1485 14179 1551 14182
rect 21173 14242 21239 14245
rect 22200 14242 23000 14272
rect 21173 14240 23000 14242
rect 21173 14184 21178 14240
rect 21234 14184 23000 14240
rect 21173 14182 23000 14184
rect 21173 14179 21239 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 22200 14152 23000 14182
rect 18270 14111 18590 14112
rect 9581 13970 9647 13973
rect 9262 13968 9647 13970
rect 9262 13912 9586 13968
rect 9642 13912 9647 13968
rect 9262 13910 9647 13912
rect 0 13834 800 13864
rect 9262 13837 9322 13910
rect 9581 13907 9647 13910
rect 19333 13970 19399 13973
rect 20437 13970 20503 13973
rect 19333 13968 20503 13970
rect 19333 13912 19338 13968
rect 19394 13912 20442 13968
rect 20498 13912 20503 13968
rect 19333 13910 20503 13912
rect 19333 13907 19399 13910
rect 20437 13907 20503 13910
rect 1761 13834 1827 13837
rect 0 13832 1827 13834
rect 0 13776 1766 13832
rect 1822 13776 1827 13832
rect 0 13774 1827 13776
rect 0 13744 800 13774
rect 1761 13771 1827 13774
rect 9213 13832 9322 13837
rect 9213 13776 9218 13832
rect 9274 13776 9322 13832
rect 9213 13774 9322 13776
rect 21541 13834 21607 13837
rect 22200 13834 23000 13864
rect 21541 13832 23000 13834
rect 21541 13776 21546 13832
rect 21602 13776 23000 13832
rect 21541 13774 23000 13776
rect 9213 13771 9279 13774
rect 21541 13771 21607 13774
rect 22200 13744 23000 13774
rect 1301 13698 1367 13701
rect 2681 13698 2747 13701
rect 1301 13696 2747 13698
rect 1301 13640 1306 13696
rect 1362 13640 2686 13696
rect 2742 13640 2747 13696
rect 1301 13638 2747 13640
rect 1301 13635 1367 13638
rect 2681 13635 2747 13638
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 0 13290 800 13320
rect 1393 13290 1459 13293
rect 0 13288 1459 13290
rect 0 13232 1398 13288
rect 1454 13232 1459 13288
rect 0 13230 1459 13232
rect 0 13200 800 13230
rect 1393 13227 1459 13230
rect 19609 13290 19675 13293
rect 20621 13290 20687 13293
rect 19609 13288 20687 13290
rect 19609 13232 19614 13288
rect 19670 13232 20626 13288
rect 20682 13232 20687 13288
rect 19609 13230 20687 13232
rect 19609 13227 19675 13230
rect 20621 13227 20687 13230
rect 21541 13290 21607 13293
rect 22200 13290 23000 13320
rect 21541 13288 23000 13290
rect 21541 13232 21546 13288
rect 21602 13232 23000 13288
rect 21541 13230 23000 13232
rect 21541 13227 21607 13230
rect 22200 13200 23000 13230
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12882 800 12912
rect 1301 12882 1367 12885
rect 0 12880 1367 12882
rect 0 12824 1306 12880
rect 1362 12824 1367 12880
rect 0 12822 1367 12824
rect 0 12792 800 12822
rect 1301 12819 1367 12822
rect 1945 12882 2011 12885
rect 2957 12882 3023 12885
rect 1945 12880 3023 12882
rect 1945 12824 1950 12880
rect 2006 12824 2962 12880
rect 3018 12824 3023 12880
rect 1945 12822 3023 12824
rect 1945 12819 2011 12822
rect 2957 12819 3023 12822
rect 10869 12882 10935 12885
rect 17861 12882 17927 12885
rect 18321 12882 18387 12885
rect 10869 12880 18387 12882
rect 10869 12824 10874 12880
rect 10930 12824 17866 12880
rect 17922 12824 18326 12880
rect 18382 12824 18387 12880
rect 10869 12822 18387 12824
rect 10869 12819 10935 12822
rect 17861 12819 17927 12822
rect 18321 12819 18387 12822
rect 21449 12882 21515 12885
rect 22200 12882 23000 12912
rect 21449 12880 23000 12882
rect 21449 12824 21454 12880
rect 21510 12824 23000 12880
rect 21449 12822 23000 12824
rect 21449 12819 21515 12822
rect 22200 12792 23000 12822
rect 5717 12746 5783 12749
rect 13721 12746 13787 12749
rect 14825 12746 14891 12749
rect 19425 12746 19491 12749
rect 5717 12744 13787 12746
rect 5717 12688 5722 12744
rect 5778 12688 13726 12744
rect 13782 12688 13787 12744
rect 5717 12686 13787 12688
rect 5717 12683 5783 12686
rect 13721 12683 13787 12686
rect 14598 12744 19491 12746
rect 14598 12688 14830 12744
rect 14886 12688 19430 12744
rect 19486 12688 19491 12744
rect 14598 12686 19491 12688
rect 14181 12610 14247 12613
rect 14598 12610 14658 12686
rect 14825 12683 14891 12686
rect 19425 12683 19491 12686
rect 14181 12608 14658 12610
rect 14181 12552 14186 12608
rect 14242 12552 14658 12608
rect 14181 12550 14658 12552
rect 14181 12547 14247 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 18689 12474 18755 12477
rect 21633 12474 21699 12477
rect 18689 12472 21699 12474
rect 18689 12416 18694 12472
rect 18750 12416 21638 12472
rect 21694 12416 21699 12472
rect 18689 12414 21699 12416
rect 18689 12411 18755 12414
rect 21633 12411 21699 12414
rect 0 12338 800 12368
rect 1853 12338 1919 12341
rect 19149 12338 19215 12341
rect 0 12336 1919 12338
rect 0 12280 1858 12336
rect 1914 12280 1919 12336
rect 0 12278 1919 12280
rect 0 12248 800 12278
rect 1853 12275 1919 12278
rect 19014 12336 19215 12338
rect 19014 12280 19154 12336
rect 19210 12280 19215 12336
rect 19014 12278 19215 12280
rect 1485 12200 1551 12205
rect 1485 12144 1490 12200
rect 1546 12144 1551 12200
rect 1485 12139 1551 12144
rect 3969 12202 4035 12205
rect 4705 12202 4771 12205
rect 6453 12202 6519 12205
rect 3969 12200 6519 12202
rect 3969 12144 3974 12200
rect 4030 12144 4710 12200
rect 4766 12144 6458 12200
rect 6514 12144 6519 12200
rect 3969 12142 6519 12144
rect 3969 12139 4035 12142
rect 4705 12139 4771 12142
rect 6453 12139 6519 12142
rect 18873 12202 18939 12205
rect 19014 12202 19074 12278
rect 19149 12275 19215 12278
rect 19977 12338 20043 12341
rect 21449 12338 21515 12341
rect 22200 12338 23000 12368
rect 19977 12336 23000 12338
rect 19977 12280 19982 12336
rect 20038 12280 21454 12336
rect 21510 12280 23000 12336
rect 19977 12278 23000 12280
rect 19977 12275 20043 12278
rect 21449 12275 21515 12278
rect 22200 12248 23000 12278
rect 18873 12200 19074 12202
rect 18873 12144 18878 12200
rect 18934 12144 19074 12200
rect 18873 12142 19074 12144
rect 18873 12139 18939 12142
rect 0 11930 800 11960
rect 1488 11930 1548 12139
rect 4889 12066 4955 12069
rect 4889 12064 5274 12066
rect 4889 12008 4894 12064
rect 4950 12008 5274 12064
rect 4889 12006 5274 12008
rect 4889 12003 4955 12006
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 0 11870 1548 11930
rect 0 11840 800 11870
rect 5214 11525 5274 12006
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 21449 11930 21515 11933
rect 22200 11930 23000 11960
rect 21449 11928 23000 11930
rect 21449 11872 21454 11928
rect 21510 11872 23000 11928
rect 21449 11870 23000 11872
rect 21449 11867 21515 11870
rect 22200 11840 23000 11870
rect 15101 11794 15167 11797
rect 17953 11794 18019 11797
rect 19517 11794 19583 11797
rect 15101 11792 19583 11794
rect 15101 11736 15106 11792
rect 15162 11736 17958 11792
rect 18014 11736 19522 11792
rect 19578 11736 19583 11792
rect 15101 11734 19583 11736
rect 15101 11731 15167 11734
rect 17953 11731 18019 11734
rect 19517 11731 19583 11734
rect 11053 11658 11119 11661
rect 15377 11658 15443 11661
rect 17769 11658 17835 11661
rect 11053 11656 17835 11658
rect 11053 11600 11058 11656
rect 11114 11600 15382 11656
rect 15438 11600 17774 11656
rect 17830 11600 17835 11656
rect 11053 11598 17835 11600
rect 11053 11595 11119 11598
rect 15377 11595 15443 11598
rect 17769 11595 17835 11598
rect 5214 11520 5323 11525
rect 5214 11464 5262 11520
rect 5318 11464 5323 11520
rect 5214 11462 5323 11464
rect 5257 11459 5323 11462
rect 18505 11522 18571 11525
rect 20069 11524 20135 11525
rect 20069 11522 20116 11524
rect 18505 11520 20116 11522
rect 18505 11464 18510 11520
rect 18566 11464 20074 11520
rect 18505 11462 20116 11464
rect 18505 11459 18571 11462
rect 20069 11460 20116 11462
rect 20180 11460 20186 11524
rect 20069 11459 20135 11460
rect 7874 11456 8194 11457
rect 0 11386 800 11416
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 1761 11386 1827 11389
rect 0 11384 1827 11386
rect 0 11328 1766 11384
rect 1822 11328 1827 11384
rect 0 11326 1827 11328
rect 0 11296 800 11326
rect 1761 11323 1827 11326
rect 21173 11386 21239 11389
rect 22200 11386 23000 11416
rect 21173 11384 23000 11386
rect 21173 11328 21178 11384
rect 21234 11328 23000 11384
rect 21173 11326 23000 11328
rect 21173 11323 21239 11326
rect 22200 11296 23000 11326
rect 10501 11250 10567 11253
rect 17953 11250 18019 11253
rect 10501 11248 18019 11250
rect 10501 11192 10506 11248
rect 10562 11192 17958 11248
rect 18014 11192 18019 11248
rect 10501 11190 18019 11192
rect 10501 11187 10567 11190
rect 17953 11187 18019 11190
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 21541 10978 21607 10981
rect 22200 10978 23000 11008
rect 21541 10976 23000 10978
rect 21541 10920 21546 10976
rect 21602 10920 23000 10976
rect 21541 10918 23000 10920
rect 21541 10915 21607 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 22200 10888 23000 10918
rect 18270 10847 18590 10848
rect 9121 10706 9187 10709
rect 19057 10706 19123 10709
rect 9121 10704 19123 10706
rect 9121 10648 9126 10704
rect 9182 10648 19062 10704
rect 19118 10648 19123 10704
rect 9121 10646 19123 10648
rect 9121 10643 9187 10646
rect 19057 10643 19123 10646
rect 1669 10570 1735 10573
rect 9438 10570 9444 10572
rect 1669 10568 9444 10570
rect 1669 10512 1674 10568
rect 1730 10512 9444 10568
rect 1669 10510 9444 10512
rect 1669 10507 1735 10510
rect 9438 10508 9444 10510
rect 9508 10508 9514 10572
rect 12341 10570 12407 10573
rect 12985 10570 13051 10573
rect 12341 10568 13051 10570
rect 12341 10512 12346 10568
rect 12402 10512 12990 10568
rect 13046 10512 13051 10568
rect 12341 10510 13051 10512
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 0 10026 800 10056
rect 1485 10026 1551 10029
rect 0 10024 1551 10026
rect 0 9968 1490 10024
rect 1546 9968 1551 10024
rect 0 9966 1551 9968
rect 9446 10026 9506 10508
rect 12341 10507 12407 10510
rect 12985 10507 13051 10510
rect 21449 10434 21515 10437
rect 22200 10434 23000 10464
rect 21449 10432 23000 10434
rect 21449 10376 21454 10432
rect 21510 10376 23000 10432
rect 21449 10374 23000 10376
rect 21449 10371 21515 10374
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 22200 10344 23000 10374
rect 14805 10303 15125 10304
rect 19333 10162 19399 10165
rect 21633 10162 21699 10165
rect 19333 10160 21699 10162
rect 19333 10104 19338 10160
rect 19394 10104 21638 10160
rect 21694 10104 21699 10160
rect 19333 10102 21699 10104
rect 19333 10099 19399 10102
rect 21633 10099 21699 10102
rect 16665 10026 16731 10029
rect 9446 10024 16731 10026
rect 9446 9968 16670 10024
rect 16726 9968 16731 10024
rect 9446 9966 16731 9968
rect 0 9936 800 9966
rect 1485 9963 1551 9966
rect 16665 9963 16731 9966
rect 21449 10026 21515 10029
rect 22200 10026 23000 10056
rect 21449 10024 23000 10026
rect 21449 9968 21454 10024
rect 21510 9968 23000 10024
rect 21449 9966 23000 9968
rect 21449 9963 21515 9966
rect 22200 9936 23000 9966
rect 15101 9890 15167 9893
rect 17217 9890 17283 9893
rect 15101 9888 17283 9890
rect 15101 9832 15106 9888
rect 15162 9832 17222 9888
rect 17278 9832 17283 9888
rect 15101 9830 17283 9832
rect 15101 9827 15167 9830
rect 17217 9827 17283 9830
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 4521 9618 4587 9621
rect 5717 9618 5783 9621
rect 4521 9616 5783 9618
rect 4521 9560 4526 9616
rect 4582 9560 5722 9616
rect 5778 9560 5783 9616
rect 4521 9558 5783 9560
rect 4521 9555 4587 9558
rect 5717 9555 5783 9558
rect 0 9482 800 9512
rect 2037 9482 2103 9485
rect 0 9480 2103 9482
rect 0 9424 2042 9480
rect 2098 9424 2103 9480
rect 0 9422 2103 9424
rect 0 9392 800 9422
rect 2037 9419 2103 9422
rect 20529 9482 20595 9485
rect 20805 9482 20871 9485
rect 20529 9480 20871 9482
rect 20529 9424 20534 9480
rect 20590 9424 20810 9480
rect 20866 9424 20871 9480
rect 20529 9422 20871 9424
rect 20529 9419 20595 9422
rect 20805 9419 20871 9422
rect 21541 9482 21607 9485
rect 22200 9482 23000 9512
rect 21541 9480 23000 9482
rect 21541 9424 21546 9480
rect 21602 9424 23000 9480
rect 21541 9422 23000 9424
rect 21541 9419 21607 9422
rect 22200 9392 23000 9422
rect 4337 9346 4403 9349
rect 7557 9346 7623 9349
rect 4337 9344 7623 9346
rect 4337 9288 4342 9344
rect 4398 9288 7562 9344
rect 7618 9288 7623 9344
rect 4337 9286 7623 9288
rect 4337 9283 4403 9286
rect 7557 9283 7623 9286
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 0 9074 800 9104
rect 1485 9074 1551 9077
rect 0 9072 1551 9074
rect 0 9016 1490 9072
rect 1546 9016 1551 9072
rect 0 9014 1551 9016
rect 0 8984 800 9014
rect 1485 9011 1551 9014
rect 21449 9074 21515 9077
rect 22200 9074 23000 9104
rect 21449 9072 23000 9074
rect 21449 9016 21454 9072
rect 21510 9016 23000 9072
rect 21449 9014 23000 9016
rect 21449 9011 21515 9014
rect 22200 8984 23000 9014
rect 2865 8938 2931 8941
rect 7005 8938 7071 8941
rect 2865 8936 7071 8938
rect 2865 8880 2870 8936
rect 2926 8880 7010 8936
rect 7066 8880 7071 8936
rect 2865 8878 7071 8880
rect 2865 8875 2931 8878
rect 7005 8875 7071 8878
rect 9857 8938 9923 8941
rect 10777 8938 10843 8941
rect 11329 8938 11395 8941
rect 18597 8938 18663 8941
rect 9857 8936 18663 8938
rect 9857 8880 9862 8936
rect 9918 8880 10782 8936
rect 10838 8880 11334 8936
rect 11390 8880 18602 8936
rect 18658 8880 18663 8936
rect 9857 8878 18663 8880
rect 9857 8875 9923 8878
rect 10777 8875 10843 8878
rect 11329 8875 11395 8878
rect 18597 8875 18663 8878
rect 4409 8736 4729 8737
rect 0 8666 800 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 1853 8666 1919 8669
rect 0 8664 1919 8666
rect 0 8608 1858 8664
rect 1914 8608 1919 8664
rect 0 8606 1919 8608
rect 0 8576 800 8606
rect 1853 8603 1919 8606
rect 21081 8666 21147 8669
rect 22200 8666 23000 8696
rect 21081 8664 23000 8666
rect 21081 8608 21086 8664
rect 21142 8608 23000 8664
rect 21081 8606 23000 8608
rect 21081 8603 21147 8606
rect 22200 8576 23000 8606
rect 4889 8530 4955 8533
rect 5441 8530 5507 8533
rect 4889 8528 5507 8530
rect 4889 8472 4894 8528
rect 4950 8472 5446 8528
rect 5502 8472 5507 8528
rect 4889 8470 5507 8472
rect 4889 8467 4955 8470
rect 5441 8467 5507 8470
rect 19977 8530 20043 8533
rect 20110 8530 20116 8532
rect 19977 8528 20116 8530
rect 19977 8472 19982 8528
rect 20038 8472 20116 8528
rect 19977 8470 20116 8472
rect 19977 8467 20043 8470
rect 20110 8468 20116 8470
rect 20180 8468 20186 8532
rect 7874 8192 8194 8193
rect 0 8122 800 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 1393 8122 1459 8125
rect 0 8120 1459 8122
rect 0 8064 1398 8120
rect 1454 8064 1459 8120
rect 0 8062 1459 8064
rect 0 8032 800 8062
rect 1393 8059 1459 8062
rect 2773 8122 2839 8125
rect 7649 8122 7715 8125
rect 2773 8120 7715 8122
rect 2773 8064 2778 8120
rect 2834 8064 7654 8120
rect 7710 8064 7715 8120
rect 2773 8062 7715 8064
rect 2773 8059 2839 8062
rect 7649 8059 7715 8062
rect 21449 8122 21515 8125
rect 22200 8122 23000 8152
rect 21449 8120 23000 8122
rect 21449 8064 21454 8120
rect 21510 8064 23000 8120
rect 21449 8062 23000 8064
rect 21449 8059 21515 8062
rect 22200 8032 23000 8062
rect 0 7714 800 7744
rect 1761 7714 1827 7717
rect 0 7712 1827 7714
rect 0 7656 1766 7712
rect 1822 7656 1827 7712
rect 0 7654 1827 7656
rect 0 7624 800 7654
rect 1761 7651 1827 7654
rect 21173 7714 21239 7717
rect 22200 7714 23000 7744
rect 21173 7712 23000 7714
rect 21173 7656 21178 7712
rect 21234 7656 23000 7712
rect 21173 7654 23000 7656
rect 21173 7651 21239 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 22200 7624 23000 7654
rect 18270 7583 18590 7584
rect 5257 7442 5323 7445
rect 5257 7440 5458 7442
rect 5257 7384 5262 7440
rect 5318 7384 5458 7440
rect 5257 7382 5458 7384
rect 5257 7379 5323 7382
rect 0 7170 800 7200
rect 1393 7170 1459 7173
rect 0 7168 1459 7170
rect 0 7112 1398 7168
rect 1454 7112 1459 7168
rect 0 7110 1459 7112
rect 0 7080 800 7110
rect 1393 7107 1459 7110
rect 5398 7037 5458 7382
rect 21449 7170 21515 7173
rect 22200 7170 23000 7200
rect 21449 7168 23000 7170
rect 21449 7112 21454 7168
rect 21510 7112 23000 7168
rect 21449 7110 23000 7112
rect 21449 7107 21515 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 22200 7080 23000 7110
rect 14805 7039 15125 7040
rect 5398 7032 5507 7037
rect 5398 6976 5446 7032
rect 5502 6976 5507 7032
rect 5398 6974 5507 6976
rect 5441 6971 5507 6974
rect 0 6762 800 6792
rect 1485 6762 1551 6765
rect 0 6760 1551 6762
rect 0 6704 1490 6760
rect 1546 6704 1551 6760
rect 0 6702 1551 6704
rect 0 6672 800 6702
rect 1485 6699 1551 6702
rect 21449 6762 21515 6765
rect 22200 6762 23000 6792
rect 21449 6760 23000 6762
rect 21449 6704 21454 6760
rect 21510 6704 23000 6760
rect 21449 6702 23000 6704
rect 21449 6699 21515 6702
rect 22200 6672 23000 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6218 800 6248
rect 1485 6218 1551 6221
rect 0 6216 1551 6218
rect 0 6160 1490 6216
rect 1546 6160 1551 6216
rect 0 6158 1551 6160
rect 0 6128 800 6158
rect 1485 6155 1551 6158
rect 21449 6218 21515 6221
rect 22200 6218 23000 6248
rect 21449 6216 23000 6218
rect 21449 6160 21454 6216
rect 21510 6160 23000 6216
rect 21449 6158 23000 6160
rect 21449 6155 21515 6158
rect 22200 6128 23000 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 21541 5810 21607 5813
rect 22200 5810 23000 5840
rect 21541 5808 23000 5810
rect 21541 5752 21546 5808
rect 21602 5752 23000 5808
rect 21541 5750 23000 5752
rect 21541 5747 21607 5750
rect 22200 5720 23000 5750
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 0 5266 800 5296
rect 1485 5266 1551 5269
rect 0 5264 1551 5266
rect 0 5208 1490 5264
rect 1546 5208 1551 5264
rect 0 5206 1551 5208
rect 0 5176 800 5206
rect 1485 5203 1551 5206
rect 21449 5266 21515 5269
rect 22200 5266 23000 5296
rect 21449 5264 23000 5266
rect 21449 5208 21454 5264
rect 21510 5208 23000 5264
rect 21449 5206 23000 5208
rect 21449 5203 21515 5206
rect 22200 5176 23000 5206
rect 7874 4928 8194 4929
rect 0 4858 800 4888
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 1669 4858 1735 4861
rect 0 4856 1735 4858
rect 0 4800 1674 4856
rect 1730 4800 1735 4856
rect 0 4798 1735 4800
rect 0 4768 800 4798
rect 1669 4795 1735 4798
rect 21265 4858 21331 4861
rect 22200 4858 23000 4888
rect 21265 4856 23000 4858
rect 21265 4800 21270 4856
rect 21326 4800 23000 4856
rect 21265 4798 23000 4800
rect 21265 4795 21331 4798
rect 22200 4768 23000 4798
rect 0 4450 800 4480
rect 1393 4450 1459 4453
rect 0 4448 1459 4450
rect 0 4392 1398 4448
rect 1454 4392 1459 4448
rect 0 4390 1459 4392
rect 0 4360 800 4390
rect 1393 4387 1459 4390
rect 21541 4450 21607 4453
rect 22200 4450 23000 4480
rect 21541 4448 23000 4450
rect 21541 4392 21546 4448
rect 21602 4392 23000 4448
rect 21541 4390 23000 4392
rect 21541 4387 21607 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 22200 4360 23000 4390
rect 18270 4319 18590 4320
rect 0 3906 800 3936
rect 1393 3906 1459 3909
rect 0 3904 1459 3906
rect 0 3848 1398 3904
rect 1454 3848 1459 3904
rect 0 3846 1459 3848
rect 0 3816 800 3846
rect 1393 3843 1459 3846
rect 21541 3906 21607 3909
rect 22200 3906 23000 3936
rect 21541 3904 23000 3906
rect 21541 3848 21546 3904
rect 21602 3848 23000 3904
rect 21541 3846 23000 3848
rect 21541 3843 21607 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22200 3816 23000 3846
rect 14805 3775 15125 3776
rect 0 3498 800 3528
rect 1393 3498 1459 3501
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3408 800 3438
rect 1393 3435 1459 3438
rect 21541 3498 21607 3501
rect 22200 3498 23000 3528
rect 21541 3496 23000 3498
rect 21541 3440 21546 3496
rect 21602 3440 23000 3496
rect 21541 3438 23000 3440
rect 21541 3435 21607 3438
rect 22200 3408 23000 3438
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 0 2954 800 2984
rect 1393 2954 1459 2957
rect 0 2952 1459 2954
rect 0 2896 1398 2952
rect 1454 2896 1459 2952
rect 0 2894 1459 2896
rect 0 2864 800 2894
rect 1393 2891 1459 2894
rect 21541 2954 21607 2957
rect 22200 2954 23000 2984
rect 21541 2952 23000 2954
rect 21541 2896 21546 2952
rect 21602 2896 23000 2952
rect 21541 2894 23000 2896
rect 21541 2891 21607 2894
rect 22200 2864 23000 2894
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 0 2546 800 2576
rect 1393 2546 1459 2549
rect 0 2544 1459 2546
rect 0 2488 1398 2544
rect 1454 2488 1459 2544
rect 0 2486 1459 2488
rect 0 2456 800 2486
rect 1393 2483 1459 2486
rect 21173 2546 21239 2549
rect 22200 2546 23000 2576
rect 21173 2544 23000 2546
rect 21173 2488 21178 2544
rect 21234 2488 23000 2544
rect 21173 2486 23000 2488
rect 21173 2483 21239 2486
rect 22200 2456 23000 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 0 2002 800 2032
rect 3509 2002 3575 2005
rect 0 2000 3575 2002
rect 0 1944 3514 2000
rect 3570 1944 3575 2000
rect 0 1942 3575 1944
rect 0 1912 800 1942
rect 3509 1939 3575 1942
rect 20529 2002 20595 2005
rect 22200 2002 23000 2032
rect 20529 2000 23000 2002
rect 20529 1944 20534 2000
rect 20590 1944 23000 2000
rect 20529 1942 23000 1944
rect 20529 1939 20595 1942
rect 22200 1912 23000 1942
rect 0 1594 800 1624
rect 1945 1594 2011 1597
rect 0 1592 2011 1594
rect 0 1536 1950 1592
rect 2006 1536 2011 1592
rect 0 1534 2011 1536
rect 0 1504 800 1534
rect 1945 1531 2011 1534
rect 20345 1594 20411 1597
rect 22200 1594 23000 1624
rect 20345 1592 23000 1594
rect 20345 1536 20350 1592
rect 20406 1536 23000 1592
rect 20345 1534 23000 1536
rect 20345 1531 20411 1534
rect 22200 1504 23000 1534
rect 0 1050 800 1080
rect 1669 1050 1735 1053
rect 0 1048 1735 1050
rect 0 992 1674 1048
rect 1730 992 1735 1048
rect 0 990 1735 992
rect 0 960 800 990
rect 1669 987 1735 990
rect 20621 1050 20687 1053
rect 22200 1050 23000 1080
rect 20621 1048 23000 1050
rect 20621 992 20626 1048
rect 20682 992 23000 1048
rect 20621 990 23000 992
rect 20621 987 20687 990
rect 22200 960 23000 990
rect 0 642 800 672
rect 2773 642 2839 645
rect 0 640 2839 642
rect 0 584 2778 640
rect 2834 584 2839 640
rect 0 582 2839 584
rect 0 552 800 582
rect 2773 579 2839 582
rect 21449 642 21515 645
rect 22200 642 23000 672
rect 21449 640 23000 642
rect 21449 584 21454 640
rect 21510 584 23000 640
rect 21449 582 23000 584
rect 21449 579 21515 582
rect 22200 552 23000 582
rect 0 234 800 264
rect 2865 234 2931 237
rect 0 232 2931 234
rect 0 176 2870 232
rect 2926 176 2931 232
rect 0 174 2931 176
rect 0 144 800 174
rect 2865 171 2931 174
rect 21265 234 21331 237
rect 22200 234 23000 264
rect 21265 232 23000 234
rect 21265 176 21270 232
rect 21326 176 23000 232
rect 21265 174 23000 176
rect 21265 171 21331 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 9444 17988 9508 18052
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 20116 11520 20180 11524
rect 20116 11464 20130 11520
rect 20130 11464 20180 11520
rect 20116 11460 20180 11464
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 9444 10508 9508 10572
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 20116 8468 20180 8532
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 9443 18052 9509 18053
rect 9443 17988 9444 18052
rect 9508 17988 9509 18052
rect 9443 17987 9509 17988
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 9446 10573 9506 17987
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 9443 10572 9509 10573
rect 9443 10508 9444 10572
rect 9508 10508 9509 10572
rect 9443 10507 9509 10508
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 20115 11524 20181 11525
rect 20115 11460 20116 11524
rect 20180 11460 20181 11524
rect 20115 11459 20181 11460
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 20118 8533 20178 11459
rect 20115 8532 20181 8533
rect 20115 8468 20116 8532
rect 20180 8468 20181 8532
rect 20115 8467 20181 8468
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__buf_1  input72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1624635492
transform 1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1624635492
transform 1 0 1932 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1624635492
transform 1 0 1656 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1624635492
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2208 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1624635492
transform -1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1624635492
transform -1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2300 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2760 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  Test_en_N_FTB01
timestamp 1624635492
transform -1 0 5060 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1624635492
transform -1 0 3588 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1624635492
transform -1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1624635492
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3864 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_43 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5060 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  prog_clk_3_N_FTB01
timestamp 1624635492
transform -1 0 5888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_56
timestamp 1624635492
transform 1 0 6256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56
timestamp 1624635492
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1624635492
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 7268 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_67
timestamp 1624635492
transform 1 0 7268 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79
timestamp 1624635492
transform 1 0 8372 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1624635492
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1624635492
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_100
timestamp 1624635492
transform 1 0 10304 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1624635492
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1624635492
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1624635492
transform -1 0 12052 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_112
timestamp 1624635492
transform 1 0 11408 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_119
timestamp 1624635492
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_106
timestamp 1624635492
transform 1 0 10856 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_131
timestamp 1624635492
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1624635492
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_127
timestamp 1624635492
transform 1 0 12788 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_139
timestamp 1624635492
transform 1 0 13892 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  clk_3_N_FTB01
timestamp 1624635492
transform -1 0 15732 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1624635492
transform 1 0 16100 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1624635492
transform -1 0 16560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_146
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_158
timestamp 1624635492
transform 1 0 15640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_162
timestamp 1624635492
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_151
timestamp 1624635492
transform 1 0 14996 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1624635492
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_168
timestamp 1624635492
transform 1 0 16560 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_175
timestamp 1624635492
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1624635492
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1624635492
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 1624635492
transform -1 0 20424 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1624635492
transform -1 0 20148 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1624635492
transform -1 0 20424 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1624635492
transform -1 0 19780 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_199
timestamp 1624635492
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_204
timestamp 1624635492
transform 1 0 19872 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1624635492
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1624635492
transform -1 0 20608 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 20792 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1624635492
transform -1 0 20700 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1624635492
transform -1 0 20976 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1624635492
transform -1 0 21068 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 1624635492
transform -1 0 21344 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input75
timestamp 1624635492
transform -1 0 21252 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1624635492
transform -1 0 21620 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1624635492
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1624635492
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1624635492
transform -1 0 1840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1624635492
transform -1 0 2024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1624635492
transform -1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1624635492
transform -1 0 2392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_14
timestamp 1624635492
transform 1 0 2392 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_26
timestamp 1624635492
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1624635492
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1624635492
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1624635492
transform 1 0 7176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1624635492
transform 1 0 8280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1624635492
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1624635492
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1624635492
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1624635492
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_156
timestamp 1624635492
transform 1 0 15456 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_168
timestamp 1624635492
transform 1 0 16560 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_180
timestamp 1624635492
transform 1 0 17664 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_192
timestamp 1624635492
transform 1 0 18768 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_201
timestamp 1624635492
transform 1 0 19596 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input77
timestamp 1624635492
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1624635492
transform -1 0 21344 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1624635492
transform -1 0 21160 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1624635492
transform -1 0 20976 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1624635492
transform -1 0 20792 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp 1624635492
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1624635492
transform -1 0 1840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_8
timestamp 1624635492
transform 1 0 1840 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_20
timestamp 1624635492
transform 1 0 2944 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1624635492
transform 1 0 4048 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1624635492
transform 1 0 5152 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_56
timestamp 1624635492
transform 1 0 6256 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1624635492
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1624635492
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1624635492
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1624635492
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1624635492
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1624635492
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_151
timestamp 1624635492
transform 1 0 14996 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_163
timestamp 1624635492
transform 1 0 16100 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_172
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1624635492
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1624635492
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_208
timestamp 1624635492
transform 1 0 20240 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input78
timestamp 1624635492
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1624635492
transform -1 0 21344 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_216
timestamp 1624635492
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624635492
transform 1 0 1656 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 2116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 2300 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_13
timestamp 1624635492
transform 1 0 2300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_25
timestamp 1624635492
transform 1 0 3404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1624635492
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1624635492
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1624635492
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1624635492
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_99
timestamp 1624635492
transform 1 0 10212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1624635492
transform 1 0 11316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1624635492
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1624635492
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_156
timestamp 1624635492
transform 1 0 15456 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_168
timestamp 1624635492
transform 1 0 16560 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_180
timestamp 1624635492
transform 1 0 17664 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_192
timestamp 1624635492
transform 1 0 18768 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_201
timestamp 1624635492
transform 1 0 19596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1624635492
transform 1 0 21344 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1624635492
transform -1 0 21344 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 21068 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 20884 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_9
timestamp 1624635492
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_21
timestamp 1624635492
transform 1 0 3036 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_33
timestamp 1624635492
transform 1 0 4140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_45
timestamp 1624635492
transform 1 0 5244 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1624635492
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1624635492
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1624635492
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1624635492
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_115
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_127
timestamp 1624635492
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_139
timestamp 1624635492
transform 1 0 13892 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_151
timestamp 1624635492
transform 1 0 14996 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1624635492
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_172
timestamp 1624635492
transform 1 0 16928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1624635492
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1624635492
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_208
timestamp 1624635492
transform 1 0 20240 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1624635492
transform -1 0 21620 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 21252 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_216
timestamp 1624635492
transform 1 0 20976 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 1840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_8
timestamp 1624635492
transform 1 0 1840 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_20
timestamp 1624635492
transform 1 0 2944 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_9
timestamp 1624635492
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_28
timestamp 1624635492
transform 1 0 3680 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_21
timestamp 1624635492
transform 1 0 3036 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_33
timestamp 1624635492
transform 1 0 4140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1624635492
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1624635492
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_45
timestamp 1624635492
transform 1 0 5244 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1624635492
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1624635492
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1624635492
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1624635492
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1624635492
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1624635492
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1624635492
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1624635492
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1624635492
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_135
timestamp 1624635492
transform 1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1624635492
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1624635492
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_156
timestamp 1624635492
transform 1 0 15456 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1624635492
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_163
timestamp 1624635492
transform 1 0 16100 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_168
timestamp 1624635492
transform 1 0 16560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_180
timestamp 1624635492
transform 1 0 17664 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1624635492
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_192
timestamp 1624635492
transform 1 0 18768 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_201
timestamp 1624635492
transform 1 0 19596 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1624635492
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_208
timestamp 1624635492
transform 1 0 20240 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 20792 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 21160 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1624635492
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1624635492
transform -1 0 21620 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 21344 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 21252 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_214
timestamp 1624635492
transform 1 0 20792 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 3312 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1624635492
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1624635492
transform 1 0 4876 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1624635492
transform 1 0 3312 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_28
timestamp 1624635492
transform 1 0 3680 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_30
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp 1624635492
transform 1 0 4600 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_50
timestamp 1624635492
transform 1 0 5704 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_62
timestamp 1624635492
transform 1 0 6808 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_74
timestamp 1624635492
transform 1 0 7912 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1624635492
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1624635492
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1624635492
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1624635492
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_156
timestamp 1624635492
transform 1 0 15456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_168
timestamp 1624635492
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_180
timestamp 1624635492
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 19596 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_192
timestamp 1624635492
transform 1 0 18768 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1624635492
transform -1 0 21620 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 21252 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1624635492
transform 1 0 2852 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_13
timestamp 1624635492
transform 1 0 2300 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1624635492
transform -1 0 3956 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1624635492
transform 1 0 4876 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_31
timestamp 1624635492
transform 1 0 3956 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1624635492
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1624635492
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_53
timestamp 1624635492
transform 1 0 5980 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_58
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8832 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1624635492
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_84
timestamp 1624635492
transform 1 0 8832 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_96
timestamp 1624635492
transform 1 0 9936 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_108
timestamp 1624635492
transform 1 0 11040 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1624635492
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1624635492
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_151
timestamp 1624635492
transform 1 0 14996 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_163
timestamp 1624635492
transform 1 0 16100 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 18400 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 19320 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_188
timestamp 1624635492
transform 1 0 18400 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_196
timestamp 1624635492
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1624635492
transform 1 0 20792 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3496 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1624635492
transform 1 0 1748 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 4692 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_26
timestamp 1624635492
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 6164 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7636 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_82
timestamp 1624635492
transform 1 0 8648 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1624635492
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1624635492
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1624635492
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1624635492
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_156
timestamp 1624635492
transform 1 0 15456 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1624635492
transform -1 0 18400 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_168
timestamp 1624635492
transform 1 0 16560 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_176
timestamp 1624635492
transform 1 0 17296 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1624635492
transform 1 0 19688 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_188
timestamp 1624635492
transform 1 0 18400 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_201
timestamp 1624635492
transform 1 0 19596 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20792 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1624635492
transform -1 0 21620 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1624635492
transform -1 0 21252 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 20976 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1624635492
transform -1 0 3312 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1624635492
transform -1 0 2484 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 1564 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_5
timestamp 1624635492
transform 1 0 1564 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1624635492
transform -1 0 5520 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 3312 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_35
timestamp 1624635492
transform 1 0 4324 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6532 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1624635492
transform -1 0 6348 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_58
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 9844 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_75
timestamp 1624635492
transform 1 0 8004 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_95
timestamp 1624635492
transform 1 0 9844 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_107
timestamp 1624635492
transform 1 0 10948 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1624635492
transform 1 0 11500 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1624635492
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1624635492
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_151
timestamp 1624635492
transform 1 0 14996 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_163
timestamp 1624635492
transform 1 0 16100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17112 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1624635492
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 19412 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 20056 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 20056 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_199
timestamp 1624635492
transform 1 0 19412 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1624635492
transform -1 0 21620 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1624635492
transform -1 0 21252 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 1656 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 1656 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1624635492
transform 1 0 3128 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_28
timestamp 1624635492
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_39
timestamp 1624635492
transform 1 0 4692 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1624635492
transform 1 0 6716 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 5796 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1624635492
transform 1 0 4968 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_60
timestamp 1624635492
transform 1 0 6624 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 7728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_72
timestamp 1624635492
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10396 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9292 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 9292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_98
timestamp 1624635492
transform 1 0 10120 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 13340 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_112
timestamp 1624635492
transform 1 0 11408 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1624635492
transform 1 0 11776 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13340 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_142
timestamp 1624635492
transform 1 0 14168 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1624635492
transform -1 0 16100 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 15088 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 16468 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1624635492
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1624635492
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 17572 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 17480 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 16652 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_178
timestamp 1624635492
transform 1 0 17480 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1624635492
transform 1 0 20148 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 20148 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_195
timestamp 1624635492
transform 1 0 19044 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_199
timestamp 1624635492
transform 1 0 19412 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_201
timestamp 1624635492
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1624635492
transform 1 0 20976 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1624635492
transform -1 0 21620 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1624635492
transform 1 0 1748 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1624635492
transform -1 0 2300 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1624635492
transform 1 0 1748 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 2668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 2484 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 2852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2392 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1624635492
transform 1 0 2116 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_17
timestamp 1624635492
transform 1 0 2668 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2852 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1624635492
transform -1 0 4508 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1624635492
transform 1 0 4508 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1624635492
transform -1 0 5428 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_30
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 6900 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 1624635492
transform 1 0 5428 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1624635492
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_58
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1624635492
transform 1 0 5336 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1624635492
transform -1 0 7176 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8648 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1624635492
transform -1 0 8004 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1624635492
transform 1 0 8004 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_82
timestamp 1624635492
transform 1 0 8648 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11408 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9752 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11408 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_84
timestamp 1624635492
transform 1 0 8832 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 1624635492
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11868 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13340 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1624635492
transform -1 0 12512 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1624635492
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_112
timestamp 1624635492
transform 1 0 11408 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 13432 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1624635492
transform -1 0 14260 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_133
timestamp 1624635492
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_133
timestamp 1624635492
transform 1 0 13340 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1624635492
transform -1 0 16560 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 16192 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 16192 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1624635492
transform 1 0 15456 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_13_150
timestamp 1624635492
transform 1 0 14904 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 19780 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_168
timestamp 1624635492
transform 1 0 16560 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_181
timestamp 1624635492
transform 1 0 17756 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_181
timestamp 1624635492
transform 1 0 17756 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1624635492
transform 1 0 20148 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1624635492
transform 1 0 19596 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_203
timestamp 1624635492
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_193
timestamp 1624635492
transform 1 0 18860 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_199
timestamp 1624635492
transform 1 0 19412 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 20792 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 21252 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 20976 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1624635492
transform -1 0 21068 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1624635492
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1624635492
transform -1 0 21620 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1624635492
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1624635492
transform 1 0 2852 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1624635492
transform -1 0 2852 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1624635492
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1624635492
transform 1 0 4324 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1624635492
transform -1 0 4324 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1624635492
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1624635492
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 6900 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_53
timestamp 1624635492
transform 1 0 5980 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7912 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7084 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_63
timestamp 1624635492
transform 1 0 6900 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9476 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11132 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_90
timestamp 1624635492
transform 1 0 9384 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 13156 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_111
timestamp 1624635492
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1624635492
transform 1 0 13156 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1624635492
transform 1 0 13708 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 13432 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1624635492
transform 1 0 14904 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1624635492
transform 1 0 15732 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_146
timestamp 1624635492
transform 1 0 14536 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1624635492
transform -1 0 17756 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 16836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1624635492
transform 1 0 17756 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1624635492
transform -1 0 20148 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1624635492
transform 1 0 20148 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1624635492
transform 1 0 18492 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 20976 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1624635492
transform -1 0 21620 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1624635492
transform -1 0 2852 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1624635492
transform 1 0 2852 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1624635492
transform -1 0 2024 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1624635492
transform 1 0 4784 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1624635492
transform -1 0 4784 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_28
timestamp 1624635492
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1624635492
transform 1 0 5612 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 7176 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_16_58
timestamp 1624635492
transform 1 0 6440 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1624635492
transform 1 0 7268 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 8924 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 8096 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_66
timestamp 1624635492
transform 1 0 7176 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_78
timestamp 1624635492
transform 1 0 8280 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9200 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1624635492
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_87
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1624635492
transform 1 0 10028 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 10764 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1624635492
transform 1 0 12236 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13064 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1624635492
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 15640 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 14904 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp 1624635492
transform 1 0 14996 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_16_150
timestamp 1624635492
transform 1 0 14904 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17112 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1624635492
transform -1 0 18400 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1624635492
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_183
timestamp 1624635492
transform 1 0 17940 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1624635492
transform -1 0 18676 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1624635492
transform 1 0 19596 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1624635492
transform 1 0 18676 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1624635492
transform 1 0 20424 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1624635492
transform -1 0 21620 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 3036 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 3956 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1624635492
transform 1 0 3036 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_30
timestamp 1624635492
transform 1 0 3864 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1624635492
transform 1 0 5428 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6532 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_56
timestamp 1624635492
transform 1 0 6256 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_58
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7452 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 8280 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_68
timestamp 1624635492
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_81
timestamp 1624635492
transform 1 0 8556 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9384 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11316 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_89
timestamp 1624635492
transform 1 0 9292 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_99
timestamp 1624635492
transform 1 0 10212 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1624635492
transform -1 0 12696 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_111
timestamp 1624635492
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 12696 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14168 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1624635492
transform 1 0 15640 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_167
timestamp 1624635492
transform 1 0 16468 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1624635492
transform 1 0 19412 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 18584 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1624635492
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_208
timestamp 1624635492
transform 1 0 20240 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1624635492
transform 1 0 20792 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 20332 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1624635492
transform -1 0 21620 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 20792 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 3036 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 4876 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1624635492
transform 1 0 3956 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_21
timestamp 1624635492
transform 1 0 3036 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_40
timestamp 1624635492
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_57
timestamp 1624635492
transform 1 0 6348 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6900 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_79
timestamp 1624635492
transform 1 0 8372 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10672 0 -1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1624635492
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_104
timestamp 1624635492
transform 1 0 10672 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11684 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_112
timestamp 1624635492
transform 1 0 11408 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_131
timestamp 1624635492
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1624635492
transform -1 0 16100 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_153
timestamp 1624635492
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_165
timestamp 1624635492
transform 1 0 16284 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1624635492
transform 1 0 17664 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1624635492
transform -1 0 17664 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1624635492
transform 1 0 18492 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1624635492
transform 1 0 20148 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624635492
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 20148 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 19964 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 19780 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1624635492
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1624635492
transform 1 0 20976 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1624635492
transform -1 0 21620 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2300 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1624635492
transform -1 0 3312 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1624635492
transform -1 0 2484 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1624635492
transform 1 0 1748 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1624635492
transform -1 0 1656 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 2300 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1624635492
transform 1 0 4600 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_30
timestamp 1624635492
transform 1 0 3864 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_38
timestamp 1624635492
transform 1 0 4600 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1624635492
transform 1 0 5428 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1624635492
transform -1 0 7636 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5704 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1624635492
transform 1 0 5520 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_56
timestamp 1624635492
transform 1 0 6256 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_58
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_52
timestamp 1624635492
transform 1 0 5888 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_60
timestamp 1624635492
transform 1 0 6624 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1624635492
transform 1 0 7636 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 8188 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1624635492
transform -1 0 7728 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1624635492
transform 1 0 7728 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 8740 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_74
timestamp 1624635492
transform 1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9568 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9660 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11316 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_87
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1624635492
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 11316 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  FILLER_19_111
timestamp 1624635492
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_108
timestamp 1624635492
transform 1 0 11040 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1624635492
transform 1 0 13616 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1624635492
transform -1 0 14260 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 14628 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1624635492
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_145
timestamp 1624635492
transform 1 0 14444 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_131
timestamp 1624635492
transform 1 0 13156 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1624635492
transform 1 0 15824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 16192 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1624635492
transform -1 0 15824 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_163
timestamp 1624635492
transform 1 0 16100 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_147
timestamp 1624635492
transform 1 0 14628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_164
timestamp 1624635492
transform 1 0 16192 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 18400 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 17572 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_176
timestamp 1624635492
transform 1 0 17296 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1624635492
transform 1 0 19044 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_197
timestamp 1624635492
transform 1 0 19228 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1624635492
transform -1 0 19320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1624635492
transform 1 0 18400 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1624635492
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 19504 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624635492
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1624635492
transform 1 0 20148 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1624635492
transform 1 0 20148 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19872 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20148 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1624635492
transform 1 0 20976 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1624635492
transform -1 0 21252 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1624635492
transform -1 0 21620 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1624635492
transform 1 0 21344 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1624635492
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1624635492
transform 1 0 2116 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2392 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform -1 0 2116 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 2852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1624635492
transform 1 0 4324 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1624635492
transform -1 0 4324 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_21
timestamp 1624635492
transform 1 0 3036 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_25
timestamp 1624635492
transform 1 0 3404 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1624635492
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_53
timestamp 1624635492
transform 1 0 5980 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8924 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1624635492
transform -1 0 9936 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9936 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_85
timestamp 1624635492
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11592 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12788 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1624635492
transform -1 0 13616 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1624635492
transform -1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_138
timestamp 1624635492
transform 1 0 13800 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1624635492
transform 1 0 15732 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1624635492
transform 1 0 14904 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_146
timestamp 1624635492
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1624635492
transform 1 0 16560 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 18400 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 19964 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1624635492
transform -1 0 20792 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_188
timestamp 1624635492
transform 1 0 18400 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1624635492
transform 1 0 20792 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1624635492
transform 1 0 2116 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2392 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1624635492
transform -1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2116 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_17
timestamp 1624635492
transform 1 0 2668 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 5336 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5520 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_46
timestamp 1624635492
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7268 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_22_64
timestamp 1624635492
transform 1 0 6992 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_83
timestamp 1624635492
transform 1 0 8740 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9936 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_98
timestamp 1624635492
transform 1 0 10120 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12604 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_110
timestamp 1624635492
transform 1 0 11224 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_122
timestamp 1624635492
transform 1 0 12328 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1624635492
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1624635492
transform 1 0 15824 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 17756 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_169
timestamp 1624635492
transform 1 0 16652 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_183
timestamp 1624635492
transform 1 0 17940 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1624635492
transform -1 0 20516 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19504 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624635492
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_195
timestamp 1624635492
transform 1 0 19044 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_201
timestamp 1624635492
transform 1 0 19596 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1624635492
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output115
timestamp 1624635492
transform 1 0 21252 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output126
timestamp 1624635492
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_211
timestamp 1624635492
transform 1 0 20516 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1624635492
transform 1 0 1748 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1624635492
transform -1 0 3772 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1624635492
transform -1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1624635492
transform -1 0 2208 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_12
timestamp 1624635492
transform 1 0 2208 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 4232 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1624635492
transform -1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_31
timestamp 1624635492
transform 1 0 3956 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1624635492
transform 1 0 5704 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1624635492
transform 1 0 5888 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_56
timestamp 1624635492
transform 1 0 6256 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7452 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 8280 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_67
timestamp 1624635492
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp 1624635492
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_87
timestamp 1624635492
transform 1 0 9108 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_99
timestamp 1624635492
transform 1 0 10212 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_104
timestamp 1624635492
transform 1 0 10672 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1624635492
transform 1 0 11684 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12972 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1624635492
transform -1 0 11592 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13800 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_138
timestamp 1624635492
transform 1 0 13800 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1624635492
transform -1 0 15548 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 15824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_146
timestamp 1624635492
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_162
timestamp 1624635492
transform 1 0 16008 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 17112 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1624635492
transform 1 0 17940 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624635492
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_170
timestamp 1624635492
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_172
timestamp 1624635492
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1624635492
transform -1 0 20332 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20056 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1624635492
transform 1 0 19596 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1624635492
transform 1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 19412 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_192
timestamp 1624635492
transform 1 0 18768 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_196
timestamp 1624635492
transform 1 0 19136 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1624635492
transform -1 0 20884 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1624635492
transform -1 0 20608 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output127
timestamp 1624635492
transform 1 0 21252 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output128
timestamp 1624635492
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1624635492
transform 1 0 1748 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1624635492
transform 1 0 2024 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 2300 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1624635492
transform -1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1624635492
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1624635492
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1624635492
transform 1 0 2944 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1624635492
transform -1 0 4324 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1624635492
transform 1 0 4324 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_28
timestamp 1624635492
transform 1 0 3680 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_30
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1624635492
transform 1 0 5152 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 5980 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1624635492
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1624635492
transform 1 0 8740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1624635492
transform 1 0 7912 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_68
timestamp 1624635492
transform 1 0 7360 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_71
timestamp 1624635492
transform 1 0 7636 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9200 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1624635492
transform -1 0 11500 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_87
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 11500 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_122
timestamp 1624635492
transform 1 0 12328 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1624635492
transform -1 0 14260 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16100 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1624635492
transform 1 0 14720 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 15548 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_159
timestamp 1624635492
transform 1 0 15732 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 19044 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1624635492
transform 1 0 19044 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1624635492
transform -1 0 20424 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624635492
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 19320 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1624635492
transform -1 0 21068 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1624635492
transform -1 0 20792 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output129
timestamp 1624635492
transform 1 0 21252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1624635492
transform -1 0 21252 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_210
timestamp 1624635492
transform 1 0 20424 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1624635492
transform 1 0 1748 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1624635492
transform 1 0 2024 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 3864 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1624635492
transform -1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_13
timestamp 1624635492
transform 1 0 2300 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1624635492
transform -1 0 5060 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_30
timestamp 1624635492
transform 1 0 3864 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1624635492
transform -1 0 5888 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1624635492
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1624635492
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_52
timestamp 1624635492
transform 1 0 5888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_58
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1624635492
transform 1 0 7636 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_80
timestamp 1624635492
transform 1 0 8464 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 10028 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1624635492
transform -1 0 10028 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11684 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1624635492
transform 1 0 11500 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 13156 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1624635492
transform -1 0 14904 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14904 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17756 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1624635492
transform -1 0 17756 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624635492
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 16836 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 19228 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1624635492
transform 1 0 20700 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1624635492
transform 1 0 21528 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_7
timestamp 1624635492
transform 1 0 1748 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1624635492
transform -1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1624635492
transform -1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1624635492
transform 1 0 1748 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_17
timestamp 1624635492
transform 1 0 2668 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_16
timestamp 1624635492
transform 1 0 2576 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_12
timestamp 1624635492
transform 1 0 2208 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1624635492
transform -1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1624635492
transform -1 0 2484 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1624635492
transform -1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 3680 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1624635492
transform 1 0 2024 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 3956 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3864 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_28
timestamp 1624635492
transform 1 0 3680 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_30
timestamp 1624635492
transform 1 0 3864 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 6164 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 5336 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1624635492
transform 1 0 5428 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_56
timestamp 1624635492
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_58
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_62
timestamp 1624635492
transform 1 0 6808 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 6900 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 8372 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1624635492
transform 1 0 7636 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_26_80
timestamp 1624635492
transform 1 0 8464 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10028 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9844 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform -1 0 9476 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_87
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_91
timestamp 1624635492
transform 1 0 9476 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_104
timestamp 1624635492
transform 1 0 10672 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1624635492
transform -1 0 11684 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13340 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624635492
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12328 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_115
timestamp 1624635492
transform 1 0 11684 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_121
timestamp 1624635492
transform 1 0 12236 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_110
timestamp 1624635492
transform 1 0 11224 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_115
timestamp 1624635492
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 14352 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 13064 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1624635492
transform -1 0 13892 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1624635492
transform -1 0 14168 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_left_track_1.prog_clk
timestamp 1624635492
transform 1 0 13892 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1624635492
transform 1 0 14168 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1624635492
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1624635492
transform 1 0 14536 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1624635492
transform 1 0 15824 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 16376 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_155
timestamp 1624635492
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_159
timestamp 1624635492
transform 1 0 15732 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_165
timestamp 1624635492
transform 1 0 16284 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_176
timestamp 1624635492
transform 1 0 17296 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_172
timestamp 1624635492
transform 1 0 16928 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1624635492
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_169
timestamp 1624635492
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624635492
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1624635492
transform 1 0 16836 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_26_183
timestamp 1624635492
transform 1 0 17940 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_180
timestamp 1624635492
transform 1 0 17664 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output141_A
timestamp 1624635492
transform -1 0 18216 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output92_A
timestamp 1624635492
transform -1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 17756 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 17848 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 17664 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 17388 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output144_A
timestamp 1624635492
transform -1 0 18676 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1624635492
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 18768 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1624635492
transform -1 0 19136 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1624635492
transform 1 0 18676 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1624635492
transform -1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624635492
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 20884 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 21068 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output130
timestamp 1624635492
transform 1 0 21252 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output131
timestamp 1624635492
transform 1 0 21252 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output132
timestamp 1624635492
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1624635492
transform -1 0 21252 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 2392 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output113
timestamp 1624635492
transform -1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_7
timestamp 1624635492
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_14
timestamp 1624635492
transform 1 0 2392 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624635492
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_26
timestamp 1624635492
transform 1 0 3496 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1624635492
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5152 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1624635492
transform -1 0 7544 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_42
timestamp 1624635492
transform 1 0 4968 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_60
timestamp 1624635492
transform 1 0 6624 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7544 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_81
timestamp 1624635492
transform 1 0 8556 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9752 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624635492
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1624635492
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_87
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1624635492
transform 1 0 9660 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1624635492
transform 1 0 12052 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1624635492
transform -1 0 12052 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_122
timestamp 1624635492
transform 1 0 12328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14720 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624635492
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_134
timestamp 1624635492
transform 1 0 13432 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_142
timestamp 1624635492
transform 1 0 14168 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_144
timestamp 1624635492
transform 1 0 14352 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15548 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16376 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1624635492
transform -1 0 17756 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17756 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_168
timestamp 1624635492
transform 1 0 16560 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1624635492
transform 1 0 19688 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 19228 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624635492
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1624635492
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1624635492
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1624635492
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_194
timestamp 1624635492
transform 1 0 18952 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_201
timestamp 1624635492
transform 1 0 19596 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1624635492
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1624635492
transform -1 0 21068 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output133
timestamp 1624635492
transform 1 0 21252 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1624635492
transform -1 0 21252 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1624635492
transform 1 0 2116 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1624635492
transform 1 0 2392 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform -1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output114
timestamp 1624635492
transform -1 0 2116 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1624635492
transform -1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1624635492
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1624635492
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_23
timestamp 1624635492
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_35
timestamp 1624635492
transform 1 0 4324 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 5428 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624635492
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_43
timestamp 1624635492
transform 1 0 5060 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_47
timestamp 1624635492
transform 1 0 5428 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_55
timestamp 1624635492
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_58
timestamp 1624635492
transform 1 0 6440 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1624635492
transform 1 0 7268 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 8372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_66
timestamp 1624635492
transform 1 0 7176 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_79
timestamp 1624635492
transform 1 0 8372 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11132 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_91
timestamp 1624635492
transform 1 0 9476 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_99
timestamp 1624635492
transform 1 0 10212 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1624635492
transform -1 0 12788 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12512 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624635492
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 11316 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_111
timestamp 1624635492
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1624635492
transform -1 0 13064 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 13064 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 13248 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_127
timestamp 1624635492
transform 1 0 12788 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_134
timestamp 1624635492
transform 1 0 13432 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_140
timestamp 1624635492
transform 1 0 13984 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_143
timestamp 1624635492
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14536 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1624635492
transform 1 0 16008 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16928 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624635492
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1624635492
transform 1 0 18400 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1624635492
transform -1 0 20056 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1624635492
transform 1 0 20056 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1624635492
transform -1 0 19780 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1624635492
transform -1 0 18952 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_191
timestamp 1624635492
transform 1 0 18676 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1624635492
transform -1 0 20884 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1624635492
transform -1 0 20608 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output116
timestamp 1624635492
transform 1 0 21252 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output134
timestamp 1624635492
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1624635492
transform -1 0 2024 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp 1624635492
transform 1 0 2024 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _113_
timestamp 1624635492
transform 1 0 2300 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _115_
timestamp 1624635492
transform 1 0 2576 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform -1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1624635492
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1624635492
transform -1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1624635492
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1624635492
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1624635492
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1624635492
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _097_
timestamp 1624635492
transform 1 0 5980 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 6440 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_42
timestamp 1624635492
transform 1 0 4968 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_50
timestamp 1624635492
transform 1 0 5704 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_56
timestamp 1624635492
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_61
timestamp 1624635492
transform 1 0 6716 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1624635492
transform -1 0 8832 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_73
timestamp 1624635492
transform 1 0 7820 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10672 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9108 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 10212 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1624635492
transform -1 0 10396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_103
timestamp 1624635492
transform 1 0 10580 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1624635492
transform 1 0 12144 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1624635492
transform -1 0 14168 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14352 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1624635492
transform 1 0 12972 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624635492
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_138
timestamp 1624635492
transform 1 0 13800 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_142
timestamp 1624635492
transform 1 0 14168 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15824 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1624635492
transform -1 0 17572 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17940 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17848 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_182
timestamp 1624635492
transform 1 0 17848 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 19596 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624635492
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_199
timestamp 1624635492
transform 1 0 19412 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output117
timestamp 1624635492
transform 1 0 21252 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 21252 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp 1624635492
transform 1 0 1748 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1624635492
transform 1 0 2024 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1624635492
transform 1 0 2300 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1624635492
transform -1 0 2852 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _114_
timestamp 1624635492
transform 1 0 2852 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform -1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1624635492
transform 1 0 3312 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3864 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1624635492
transform 1 0 3588 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 3312 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1624635492
transform 1 0 6072 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624635492
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform -1 0 5152 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_44
timestamp 1624635492
transform 1 0 5152 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_52
timestamp 1624635492
transform 1 0 5888 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_58
timestamp 1624635492
transform 1 0 6440 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 9200 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_70
timestamp 1624635492
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1624635492
transform 1 0 10672 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9200 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 13156 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624635492
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 11224 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform -1 0 11408 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_107
timestamp 1624635492
transform 1 0 10948 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 13156 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1624635492
transform -1 0 15732 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1624635492
transform 1 0 15732 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1624635492
transform 1 0 16100 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1624635492
transform 1 0 16376 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1624635492
transform -1 0 15456 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_31_162
timestamp 1624635492
transform 1 0 16008 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1624635492
transform 1 0 16928 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1624635492
transform -1 0 18308 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1624635492
transform 1 0 18308 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1624635492
transform -1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624635492
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1624635492
transform 1 0 18768 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1624635492
transform 1 0 19044 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1624635492
transform 1 0 19872 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1624635492
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output118
timestamp 1624635492
transform 1 0 21252 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output145
timestamp 1624635492
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1624635492
transform 1 0 20700 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1624635492
transform -1 0 2392 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _111_
timestamp 1624635492
transform 1 0 2392 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624635492
transform 1 0 2668 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1624635492
transform 1 0 2944 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform -1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1624635492
transform -1 0 2116 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624635492
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 1624635492
transform 1 0 3220 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1624635492
transform -1 0 3772 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1624635492
transform 1 0 3864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1624635492
transform 1 0 4140 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1624635492
transform -1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1624635492
transform -1 0 4784 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1624635492
transform -1 0 4968 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1624635492
transform -1 0 6532 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1624635492
transform -1 0 5152 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1624635492
transform -1 0 5336 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output155_A
timestamp 1624635492
transform 1 0 5336 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_48
timestamp 1624635492
transform 1 0 5520 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_56
timestamp 1624635492
transform 1 0 6256 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_59
timestamp 1624635492
transform 1 0 6532 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1624635492
transform -1 0 9016 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1624635492
transform -1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1624635492
transform -1 0 8188 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1624635492
transform -1 0 8004 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1624635492
transform -1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_69
timestamp 1624635492
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9936 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9108 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624635492
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12328 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12604 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1624635492
transform -1 0 12880 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_112
timestamp 1624635492
transform 1 0 11408 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1624635492
transform -1 0 13156 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14076 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1624635492
transform -1 0 15180 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624635492
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 14260 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_131
timestamp 1624635492
transform 1 0 13156 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1624635492
transform -1 0 15456 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 15732 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 16376 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 16652 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624635492
transform -1 0 15916 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 15916 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1624635492
transform -1 0 17020 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output152
timestamp 1624635492
transform -1 0 17572 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output153
timestamp 1624635492
transform -1 0 17940 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output154
timestamp 1624635492
transform -1 0 18400 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1624635492
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_169
timestamp 1624635492
transform 1 0 16652 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_183
timestamp 1624635492
transform 1 0 17940 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1624635492
transform -1 0 20240 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1624635492
transform -1 0 19964 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1624635492
transform -1 0 19504 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1624635492
transform -1 0 19228 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1624635492
transform 1 0 18676 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1624635492
transform -1 0 18676 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624635492
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output144
timestamp 1624635492
transform 1 0 20240 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1624635492
transform 1 0 19596 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1624635492
transform -1 0 21252 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output119
timestamp 1624635492
transform 1 0 21252 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output141
timestamp 1624635492
transform -1 0 20976 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1624635492
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1624635492
transform 1 0 1748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform -1 0 2484 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1624635492
transform -1 0 2852 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1624635492
transform -1 0 3220 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624635492
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform -1 0 4784 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1624635492
transform -1 0 3588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1624635492
transform -1 0 4232 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output155
timestamp 1624635492
transform -1 0 5152 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1624635492
transform -1 0 3772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1624635492
transform -1 0 4416 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_44
timestamp 1624635492
transform 1 0 5152 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output156
timestamp 1624635492
transform -1 0 5612 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_49
timestamp 1624635492
transform 1 0 5612 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1624635492
transform 1 0 5704 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_53
timestamp 1624635492
transform 1 0 5980 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1624635492
transform 1 0 6072 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1624635492
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1624635492
transform 1 0 6532 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624635492
transform 1 0 6440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 6992 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1624635492
transform -1 0 7268 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1624635492
transform 1 0 7360 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1624635492
transform 1 0 7820 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1624635492
transform 1 0 8188 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1624635492
transform 1 0 8648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1624635492
transform -1 0 7820 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1624635492
transform -1 0 8648 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_67
timestamp 1624635492
transform 1 0 7268 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_76
timestamp 1624635492
transform 1 0 8096 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624635492
transform 1 0 9108 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1624635492
transform -1 0 10212 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1624635492
transform -1 0 10672 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1624635492
transform 1 0 9200 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1624635492
transform -1 0 9752 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1624635492
transform -1 0 9936 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1624635492
transform -1 0 9108 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_104
timestamp 1624635492
transform 1 0 10672 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624635492
transform 1 0 11776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1624635492
transform -1 0 11040 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1624635492
transform -1 0 11500 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1624635492
transform 1 0 11868 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1624635492
transform 1 0 12144 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1624635492
transform -1 0 12788 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1624635492
transform -1 0 11776 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_123
timestamp 1624635492
transform 1 0 12420 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624635492
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1624635492
transform -1 0 13156 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output149
timestamp 1624635492
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output150
timestamp 1624635492
transform 1 0 13708 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output151
timestamp 1624635492
transform 1 0 13340 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 13340 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_127
timestamp 1624635492
transform 1 0 12788 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output135
timestamp 1624635492
transform -1 0 14904 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output142
timestamp 1624635492
transform 1 0 16376 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output143
timestamp 1624635492
transform 1 0 16008 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output146
timestamp 1624635492
transform -1 0 15272 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output147
timestamp 1624635492
transform -1 0 15640 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output148
timestamp 1624635492
transform -1 0 16008 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624635492
transform 1 0 17112 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output136
timestamp 1624635492
transform 1 0 18308 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output137
timestamp 1624635492
transform 1 0 17940 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output138
timestamp 1624635492
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output139
timestamp 1624635492
transform 1 0 17204 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output140
timestamp 1624635492
transform 1 0 16744 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1624635492
transform -1 0 20148 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624635492
transform 1 0 19780 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output122
timestamp 1624635492
transform 1 0 20148 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output123
timestamp 1624635492
transform 1 0 19412 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output124
timestamp 1624635492
transform 1 0 19044 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output125
timestamp 1624635492
transform 1 0 18676 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform 1 0 21252 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output120
timestamp 1624635492
transform 1 0 20884 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output121
timestamp 1624635492
transform 1 0 20516 0 1 20128
box -38 -48 406 592
<< labels >>
rlabel metal2 s 202 22200 258 23000 6 SC_IN_TOP
port 0 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 SC_OUT_TOP
port 1 nsew signal tristate
rlabel metal2 s 4434 22200 4490 23000 6 Test_en_N_out
port 2 nsew signal tristate
rlabel metal2 s 20718 0 20774 800 6 Test_en_S_in
port 3 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 ccff_head
port 4 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 ccff_tail
port 5 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[0]
port 6 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[10]
port 7 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[11]
port 8 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[12]
port 9 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[13]
port 10 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[14]
port 11 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[15]
port 12 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[16]
port 13 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 14 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[18]
port 15 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_in[19]
port 16 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[1]
port 17 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[2]
port 18 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[3]
port 19 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[4]
port 20 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[5]
port 21 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[6]
port 22 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[7]
port 23 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[8]
port 24 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[9]
port 25 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[0]
port 26 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[10]
port 27 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 28 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[12]
port 29 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 30 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[14]
port 31 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[15]
port 32 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[16]
port 33 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[17]
port 34 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[18]
port 35 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 chanx_left_out[19]
port 36 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[1]
port 37 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[2]
port 38 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[3]
port 39 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[4]
port 40 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[5]
port 41 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[6]
port 42 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[7]
port 43 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[8]
port 44 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[9]
port 45 nsew signal tristate
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[0]
port 46 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[10]
port 47 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[11]
port 48 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[12]
port 49 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[13]
port 50 nsew signal input
rlabel metal3 s 22200 10888 23000 11008 6 chanx_right_in[14]
port 51 nsew signal input
rlabel metal3 s 22200 11296 23000 11416 6 chanx_right_in[15]
port 52 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[16]
port 53 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[17]
port 54 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_in[18]
port 55 nsew signal input
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_in[19]
port 56 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[1]
port 57 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[2]
port 58 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[3]
port 59 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[4]
port 60 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[5]
port 61 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[6]
port 62 nsew signal input
rlabel metal3 s 22200 7624 23000 7744 6 chanx_right_in[7]
port 63 nsew signal input
rlabel metal3 s 22200 8032 23000 8152 6 chanx_right_in[8]
port 64 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[9]
port 65 nsew signal input
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[0]
port 66 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[10]
port 67 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[11]
port 68 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[12]
port 69 nsew signal tristate
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[13]
port 70 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[14]
port 71 nsew signal tristate
rlabel metal3 s 22200 20680 23000 20800 6 chanx_right_out[15]
port 72 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[16]
port 73 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[17]
port 74 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[18]
port 75 nsew signal tristate
rlabel metal3 s 22200 22584 23000 22704 6 chanx_right_out[19]
port 76 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[1]
port 77 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[2]
port 78 nsew signal tristate
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[3]
port 79 nsew signal tristate
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[4]
port 80 nsew signal tristate
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[5]
port 81 nsew signal tristate
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[6]
port 82 nsew signal tristate
rlabel metal3 s 22200 17008 23000 17128 6 chanx_right_out[7]
port 83 nsew signal tristate
rlabel metal3 s 22200 17416 23000 17536 6 chanx_right_out[8]
port 84 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[9]
port 85 nsew signal tristate
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[0]
port 86 nsew signal input
rlabel metal2 s 9954 22200 10010 23000 6 chany_top_in[10]
port 87 nsew signal input
rlabel metal2 s 10414 22200 10470 23000 6 chany_top_in[11]
port 88 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[12]
port 89 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[13]
port 90 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[14]
port 91 nsew signal input
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_in[15]
port 92 nsew signal input
rlabel metal2 s 12530 22200 12586 23000 6 chany_top_in[16]
port 93 nsew signal input
rlabel metal2 s 12898 22200 12954 23000 6 chany_top_in[17]
port 94 nsew signal input
rlabel metal2 s 13358 22200 13414 23000 6 chany_top_in[18]
port 95 nsew signal input
rlabel metal2 s 13818 22200 13874 23000 6 chany_top_in[19]
port 96 nsew signal input
rlabel metal2 s 6090 22200 6146 23000 6 chany_top_in[1]
port 97 nsew signal input
rlabel metal2 s 6550 22200 6606 23000 6 chany_top_in[2]
port 98 nsew signal input
rlabel metal2 s 7010 22200 7066 23000 6 chany_top_in[3]
port 99 nsew signal input
rlabel metal2 s 7378 22200 7434 23000 6 chany_top_in[4]
port 100 nsew signal input
rlabel metal2 s 7838 22200 7894 23000 6 chany_top_in[5]
port 101 nsew signal input
rlabel metal2 s 8206 22200 8262 23000 6 chany_top_in[6]
port 102 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[7]
port 103 nsew signal input
rlabel metal2 s 9126 22200 9182 23000 6 chany_top_in[8]
port 104 nsew signal input
rlabel metal2 s 9494 22200 9550 23000 6 chany_top_in[9]
port 105 nsew signal input
rlabel metal2 s 14186 22200 14242 23000 6 chany_top_out[0]
port 106 nsew signal tristate
rlabel metal2 s 18510 22200 18566 23000 6 chany_top_out[10]
port 107 nsew signal tristate
rlabel metal2 s 18878 22200 18934 23000 6 chany_top_out[11]
port 108 nsew signal tristate
rlabel metal2 s 19338 22200 19394 23000 6 chany_top_out[12]
port 109 nsew signal tristate
rlabel metal2 s 19706 22200 19762 23000 6 chany_top_out[13]
port 110 nsew signal tristate
rlabel metal2 s 20166 22200 20222 23000 6 chany_top_out[14]
port 111 nsew signal tristate
rlabel metal2 s 20626 22200 20682 23000 6 chany_top_out[15]
port 112 nsew signal tristate
rlabel metal2 s 20994 22200 21050 23000 6 chany_top_out[16]
port 113 nsew signal tristate
rlabel metal2 s 21454 22200 21510 23000 6 chany_top_out[17]
port 114 nsew signal tristate
rlabel metal2 s 21914 22200 21970 23000 6 chany_top_out[18]
port 115 nsew signal tristate
rlabel metal2 s 22282 22200 22338 23000 6 chany_top_out[19]
port 116 nsew signal tristate
rlabel metal2 s 14646 22200 14702 23000 6 chany_top_out[1]
port 117 nsew signal tristate
rlabel metal2 s 15106 22200 15162 23000 6 chany_top_out[2]
port 118 nsew signal tristate
rlabel metal2 s 15474 22200 15530 23000 6 chany_top_out[3]
port 119 nsew signal tristate
rlabel metal2 s 15934 22200 15990 23000 6 chany_top_out[4]
port 120 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[5]
port 121 nsew signal tristate
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[6]
port 122 nsew signal tristate
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[7]
port 123 nsew signal tristate
rlabel metal2 s 17590 22200 17646 23000 6 chany_top_out[8]
port 124 nsew signal tristate
rlabel metal2 s 18050 22200 18106 23000 6 chany_top_out[9]
port 125 nsew signal tristate
rlabel metal2 s 4802 22200 4858 23000 6 clk_3_N_out
port 126 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 clk_3_S_in
port 127 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_11_
port 128 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_13_
port 129 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_15_
port 130 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 left_bottom_grid_pin_17_
port 131 nsew signal input
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_1_
port 132 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_3_
port 133 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_5_
port 134 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_7_
port 135 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_9_
port 136 nsew signal input
rlabel metal2 s 3974 22200 4030 23000 6 prog_clk_0_N_in
port 137 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 prog_clk_3_N_out
port 138 nsew signal tristate
rlabel metal2 s 11518 0 11574 800 6 prog_clk_3_S_in
port 139 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_11_
port 140 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_13_
port 141 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_15_
port 142 nsew signal input
rlabel metal3 s 22200 3816 23000 3936 6 right_bottom_grid_pin_17_
port 143 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_1_
port 144 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_3_
port 145 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_5_
port 146 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_7_
port 147 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_9_
port 148 nsew signal input
rlabel metal2 s 570 22200 626 23000 6 top_left_grid_pin_42_
port 149 nsew signal input
rlabel metal2 s 1030 22200 1086 23000 6 top_left_grid_pin_43_
port 150 nsew signal input
rlabel metal2 s 1398 22200 1454 23000 6 top_left_grid_pin_44_
port 151 nsew signal input
rlabel metal2 s 1858 22200 1914 23000 6 top_left_grid_pin_45_
port 152 nsew signal input
rlabel metal2 s 2318 22200 2374 23000 6 top_left_grid_pin_46_
port 153 nsew signal input
rlabel metal2 s 2686 22200 2742 23000 6 top_left_grid_pin_47_
port 154 nsew signal input
rlabel metal2 s 3146 22200 3202 23000 6 top_left_grid_pin_48_
port 155 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 top_left_grid_pin_49_
port 156 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 157 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 158 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 159 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 160 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 161 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
