* NGSPICE file created from bottom_left_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

.subckt bottom_left_tile VGND VPWR ccff_head ccff_tail chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[20] chanx_right_in[21] chanx_right_in[22] chanx_right_in[23] chanx_right_in[24]
+ chanx_right_in[25] chanx_right_in[26] chanx_right_in[27] chanx_right_in[28] chanx_right_in[29]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[20] chanx_right_out[21] chanx_right_out[22]
+ chanx_right_out[23] chanx_right_out[24] chanx_right_out[25] chanx_right_out[26]
+ chanx_right_out[27] chanx_right_out[28] chanx_right_out[29] chanx_right_out[2] chanx_right_out[3]
+ chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8]
+ chanx_right_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[20] chany_top_in[21]
+ chany_top_in[22] chany_top_in[23] chany_top_in[24] chany_top_in[25] chany_top_in[26]
+ chany_top_in[27] chany_top_in[28] chany_top_in[29] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[20] chany_top_out[21]
+ chany_top_out[22] chany_top_out[23] chany_top_out[24] chany_top_out[25] chany_top_out[26]
+ chany_top_out[27] chany_top_out[28] chany_top_out[29] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] prog_clk prog_reset_top_in reset_top_in right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_ right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_ test_enable_top_in
+ top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
+ top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_ top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_0.mux_l1_in_1_ net141 net22 sb_0__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_49_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_131_ sb_0__0_.mux_top_track_0.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_32.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_34.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_10.mux_l2_in_0_ net160 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_10.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_114_ sb_0__0_.mux_top_track_34.out VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_2.mux_l1_in_0_ net64 net53 sb_0__0_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_44_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_5 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_top_track_12.mux_l2_in_0_ net143 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_12.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput75 net75 VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_12
Xoutput97 net97 VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_12
Xoutput86 net86 VGND VGND VPWR VPWR chanx_right_out[22] sky130_fd_sc_hd__buf_12
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk
+ sb_0__0_.mem_right_track_44.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_44.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_0.mux_l1_in_0_ net70 net67 sb_0__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_130_ sb_0__0_.mux_top_track_2.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_113_ net3 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_44.mux_l2_in_0__153 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_44.mux_l2_in_0__153/HI
+ net153 sky130_fd_sc_hd__conb_1
XFILLER_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_right_track_10.mux_l1_in_0_ net65 net49 sb_0__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_6 net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_12.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_12.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_89_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput76 net76 VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_12
Xoutput98 net98 VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput87 net87 VGND VGND VPWR VPWR chanx_right_out[23] sky130_fd_sc_hd__buf_12
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_34.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_44.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk
+ sb_0__0_.mem_right_track_0.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_12.mux_l1_in_0_ net16 net67 sb_0__0_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_27_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__0_.mux_top_track_28.mux_l2_in_0__148 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_28.mux_l2_in_0__148/HI
+ net148 sky130_fd_sc_hd__conb_1
XFILLER_14_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_32.out sky130_fd_sc_hd__clkbuf_1
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_112_ net31 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_494 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_7 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_10.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_12.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput99 net99 VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_12
Xoutput77 net77 VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_12
Xoutput88 net88 VGND VGND VPWR VPWR chanx_right_out[24] sky130_fd_sc_hd__buf_12
XFILLER_88_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk
+ sb_0__0_.mem_right_track_0.ccff_head net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_34.mux_l2_in_0_ net133 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_34.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_2__leaf_prog_clk
+ sb_0__0_.mem_right_track_18.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_18.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_6.mux_l1_in_1__139 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_6.mux_l1_in_1__139/HI
+ net139 sky130_fd_sc_hd__conb_1
XFILLER_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_6.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_6.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_111_ net30 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_8 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_48.out sky130_fd_sc_hd__clkbuf_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput78 net78 VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_12
Xoutput89 net89 VGND VGND VPWR VPWR chanx_right_out[25] sky130_fd_sc_hd__buf_12
XFILLER_88_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_14.out sky130_fd_sc_hd__clkbuf_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_16.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_18.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_34.mux_l1_in_0_ net66 net36 sb_0__0_.mem_right_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_4.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_6.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_64_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_30.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_30.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_right_track_46.mux_l2_in_0_ net136 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_46.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__0_.mux_top_track_12.mux_l2_in_0__143 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_12.mux_l2_in_0__143/HI
+ net143 sky130_fd_sc_hd__conb_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_110_ net29 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_9 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_right_track_16.mux_l2_in_0__163 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_16.mux_l2_in_0__163/HI
+ net163 sky130_fd_sc_hd__conb_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput79 net79 VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mux_top_track_48.mux_l2_in_0_ net155 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_48.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_50.mux_l2_in_0_ net156 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_0.ccff_head VGND VGND VPWR VPWR sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_28.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_30.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_right_track_46.mux_l1_in_0_ net64 net59 sb_0__0_.mem_right_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_0.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_top_track_48.mux_l1_in_0_ net26 net69 sb_0__0_.mem_top_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_top_track_50.mux_l1_in_0_ net25 net70 sb_0__0_.mem_top_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_78_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_34.mux_l2_in_0__133 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_34.mux_l2_in_0__133/HI
+ net133 sky130_fd_sc_hd__conb_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_099_ sb_0__0_.mux_right_track_4.out VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk sb_0__0_.mem_top_track_44.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk net1
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_8.mux_l2_in_0_ net140 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_10.ccff_head VGND VGND VPWR VPWR sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_55_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_6.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_19_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_098_ sb_0__0_.mux_right_track_6.out VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_6.mux_l2_in_0_ sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__0_.mem_top_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_4.mux_l2_in_0__134 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_4.mux_l2_in_0__134/HI
+ net134 sky130_fd_sc_hd__conb_1
XFILLER_86_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk sb_0__0_.mem_top_track_12.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_74_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_0.mux_l1_in_1__141 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_0.mux_l1_in_1__141/HI
+ net141 sky130_fd_sc_hd__conb_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_34.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_79_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_top_track_6.mux_l1_in_1_ net157 net19 sb_0__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_16.mux_l2_in_0_ net163 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_16.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_4.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_8.mux_l1_in_0_ net64 net50 sb_0__0_.mem_right_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_27_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_097_ sb_0__0_.mux_right_track_8.out VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_4__leaf_prog_clk sb_0__0_.mem_top_track_10.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_18.mux_l2_in_0_ net146 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_18.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_30.mux_l2_in_0__149 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_30.mux_l2_in_0__149/HI
+ net149 sky130_fd_sc_hd__conb_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_top_track_6.mux_l1_in_0_ net70 net67 sb_0__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_18.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_18.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_top_track_2.mux_l2_in_0__147 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_2.mux_l2_in_0__147/HI
+ net147 sky130_fd_sc_hd__conb_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_16.out sky130_fd_sc_hd__clkbuf_1
XFILLER_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_096_ sb_0__0_.mux_right_track_10.out VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_16.mux_l1_in_0_ net65 net46 sb_0__0_.mem_right_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_28.mux_l2_in_0_ net166 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_28.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_079_ sb_0__0_.mux_right_track_44.out VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_30.mux_l2_in_0_ net167 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_30.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_48.mux_l2_in_0__137 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_48.mux_l2_in_0__137/HI
+ net137 sky130_fd_sc_hd__conb_1
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_50.out sky130_fd_sc_hd__clkbuf_1
XFILLER_88_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_18.mux_l1_in_0_ net12 net70 sb_0__0_.mem_top_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_16.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_18.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_32.mux_l2_in_0_ net150 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_32.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk sb_0__0_.mem_top_track_30.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_30.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_10.mux_l2_in_0__142 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_10.mux_l2_in_0__142/HI
+ net142 sky130_fd_sc_hd__conb_1
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_59_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_095_ sb_0__0_.mux_right_track_12.out VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_28.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_28.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_078_ sb_0__0_.mux_right_track_46.out VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_14.mux_l2_in_0__162 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_14.mux_l2_in_0__162/HI
+ net162 sky130_fd_sc_hd__conb_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_28.mux_l1_in_0_ net63 net39 sb_0__0_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_30.mux_l1_in_0_ net64 net38 sb_0__0_.mem_right_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_28.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_30.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_77_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_0__0_.mux_top_track_32.mux_l1_in_0_ net5 net69 sb_0__0_.mem_top_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_44.mux_l2_in_0_ net153 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_44.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_91_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_094_ sb_0__0_.mux_right_track_14.out VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
XFILLER_49_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_2__leaf_prog_clk
+ sb_0__0_.mem_right_track_18.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_28.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_32.out sky130_fd_sc_hd__clkbuf_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_077_ sb_0__0_.mux_right_track_48.out VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_129_ sb_0__0_.mux_top_track_4.out VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_32.mux_l2_in_0__132 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_32.mux_l2_in_0__132/HI
+ net132 sky130_fd_sc_hd__conb_1
XFILLER_67_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_093_ sb_0__0_.mux_right_track_16.out VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput1 ccff_head VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_2.mux_l2_in_0__165 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_2.mux_l2_in_0__165/HI
+ net165 sky130_fd_sc_hd__conb_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_076_ sb_0__0_.mux_right_track_50.out VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_44.mux_l1_in_0_ net28 net67 sb_0__0_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_128_ sb_0__0_.mux_top_track_6.out VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput70 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND VPWR
+ VPWR net70 sky130_fd_sc_hd__buf_2
XFILLER_67_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_48.out sky130_fd_sc_hd__clkbuf_1
XFILLER_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_46.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_46.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_57_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_092_ sb_0__0_.mux_right_track_18.out VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
XFILLER_40_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 chanx_right_in[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_68_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_075_ net56 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_127_ sb_0__0_.mux_top_track_8.out VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_right_track_4.mux_l2_in_0_ net134 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_4.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_87_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput60 chany_top_in[8] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_14.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_14.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_top_track_2.mux_l2_in_0_ net147 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_2.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_44.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_46.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_3__leaf_prog_clk
+ sb_0__0_.mem_right_track_2.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_0__0_.mux_right_track_28.mux_l2_in_0__166 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_28.mux_l2_in_0__166/HI
+ net166 sky130_fd_sc_hd__conb_1
XFILLER_59_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_091_ net44 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
XFILLER_40_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput3 chanx_right_in[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_074_ net55 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_126_ sb_0__0_.mux_top_track_10.out VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput50 chany_top_in[26] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
Xinput61 chany_top_in[9] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_12.mux_l2_in_0_ net161 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_12.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_109_ sb_0__0_.mux_top_track_44.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_12.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_14.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_4.mux_l1_in_0_ net65 net52 sb_0__0_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_14.mux_l2_in_0_ net144 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_14.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_95_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_3__leaf_prog_clk
+ sb_0__0_.mem_right_track_0.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_54_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_090_ net42 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput4 chanx_right_in[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_2.mux_l1_in_0_ net21 net68 sb_0__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_073_ net54 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_8.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_10.ccff_head
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_125_ sb_0__0_.mux_top_track_12.out VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_46.mux_l2_in_0__136 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_46.mux_l2_in_0__136/HI
+ net136 sky130_fd_sc_hd__conb_1
Xinput40 chany_top_in[17] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput62 prog_reset_top_in VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_12
Xinput51 chany_top_in[27] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_108_ sb_0__0_.mux_top_track_46.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_2
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_12.mux_l1_in_0_ net63 net48 sb_0__0_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_22_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 chanx_right_in[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_83_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_28.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_14.mux_l1_in_0_ net15 net68 sb_0__0_.mem_top_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_072_ net43 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xsb_0__0_.mux_right_track_50.mux_l2_in_0__138 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_50.mux_l2_in_0__138/HI
+ net138 sky130_fd_sc_hd__conb_1
XFILLER_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_12.mux_l2_in_0__161 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_12.mux_l2_in_0__161/HI
+ net161 sky130_fd_sc_hd__conb_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_10 clknet_3_6__leaf_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_6.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_8.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_32.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_32.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_124_ sb_0__0_.mux_top_track_14.out VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_93_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput30 chanx_right_in[8] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 chany_top_in[28] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
Xinput41 chany_top_in[18] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
Xinput63 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND
+ VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_34.out sky130_fd_sc_hd__clkbuf_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_107_ sb_0__0_.mux_top_track_48.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput6 chanx_right_in[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_18.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_30.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_32.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_123_ sb_0__0_.mux_top_track_16.out VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput31 chanx_right_in[9] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 chanx_right_in[26] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput53 chany_top_in[29] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput42 chany_top_in[19] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND
+ VPWR VPWR net64 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_106_ sb_0__0_.mux_top_track_50.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_2.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput7 chanx_right_in[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_16.out sky130_fd_sc_hd__clkbuf_1
XFILLER_46_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput130 net130 VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_12
XFILLER_75_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_122_ sb_0__0_.mux_top_track_18.out VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput21 chanx_right_in[27] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 chanx_right_in[17] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput43 chany_top_in[1] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xinput54 chany_top_in[2] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 chany_top_in[0] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput65 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND
+ VPWR VPWR net65 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_105_ net24 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_48.mux_l2_in_0_ net137 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_48.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_50.mux_l2_in_0_ net138 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
+ net71 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_84_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_6__leaf_prog_clk sb_0__0_.mem_top_track_46.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_46.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_89_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_50.out sky130_fd_sc_hd__clkbuf_1
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_50.mem_out\[0\] net62 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfrtp_4
XFILLER_58_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_0.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 chanx_right_in[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput131 net131 VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_12
Xoutput120 net120 VGND VGND VPWR VPWR chany_top_out[26] sky130_fd_sc_hd__buf_12
XFILLER_28_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_121_ net11 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 chanx_right_in[28] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xsb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk sb_0__0_.mem_top_track_8.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xinput11 chanx_right_in[18] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 chany_top_in[20] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput55 chany_top_in[3] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput33 chany_top_in[10] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput66 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND
+ VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_104_ net13 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk sb_0__0_.mem_top_track_14.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk sb_0__0_.mem_top_track_44.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_46.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_89_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_48.mux_l1_in_0_ net65 net58 sb_0__0_.mem_right_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_50.mux_l1_in_0_ net66 net57 sb_0__0_.mem_right_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_67_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_48.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_50.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 chanx_right_in[16] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_0.mux_l2_in_0_ sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__0_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput110 net110 VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_12
Xoutput121 net121 VGND VGND VPWR VPWR chany_top_out[27] sky130_fd_sc_hd__buf_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_120_ net10 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_right_track_0.mux_l1_in_1_ net159 net66 sb_0__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_6.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xinput12 chanx_right_in[19] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput45 chany_top_in[21] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput34 chany_top_in[11] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput23 chanx_right_in[29] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput56 chany_top_in[4] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput67 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND VPWR
+ VPWR net67 sky130_fd_sc_hd__buf_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_103_ net2 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_4__leaf_prog_clk sb_0__0_.mem_top_track_12.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_30.mux_l2_in_0__167 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_30.mux_l2_in_0__167/HI
+ net167 sky130_fd_sc_hd__conb_1
XFILLER_31_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput100 net100 VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_12
Xoutput122 net122 VGND VGND VPWR VPWR chany_top_out[28] sky130_fd_sc_hd__buf_12
Xoutput111 net111 VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_0.mux_l1_in_0_ net63 net32 sb_0__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_34.mux_l2_in_0__151 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_34.mux_l2_in_0__151/HI
+ net151 sky130_fd_sc_hd__conb_1
XFILLER_46_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput13 chanx_right_in[1] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
Xinput46 chany_top_in[22] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput35 chany_top_in[12] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 chanx_right_in[2] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput57 chany_top_in[5] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput68 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND VPWR
+ VPWR net68 sky130_fd_sc_hd__buf_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_44.mux_l2_in_0__135 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_44.mux_l2_in_0__135/HI
+ net135 sky130_fd_sc_hd__conb_1
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_102_ net23 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_10.mux_l2_in_0_ net142 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_10.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_8.mux_l2_in_0_ net158 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_10.ccff_head VGND VGND VPWR VPWR sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_0__0_.mux_right_track_0.mux_l1_in_1__159 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_0.mux_l1_in_1__159/HI
+ net159 sky130_fd_sc_hd__conb_1
XFILLER_89_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_top_track_18.mux_l2_in_0__146 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_18.mux_l2_in_0__146/HI
+ net146 sky130_fd_sc_hd__conb_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_0__0_.mux_right_track_10.mux_l2_in_0__160 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_10.mux_l2_in_0__160/HI
+ net160 sky130_fd_sc_hd__conb_1
XFILLER_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput101 net101 VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chany_top_out[29] sky130_fd_sc_hd__buf_12
Xoutput112 net112 VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_32.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_32.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_87_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput36 chany_top_in[13] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 chanx_right_in[3] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 chanx_right_in[20] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput47 chany_top_in[23] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
Xinput58 chany_top_in[6] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
Xinput69 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND VPWR
+ VPWR net69 sky130_fd_sc_hd__buf_2
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_18.mux_l2_in_0_ net164 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_18.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_101_ sb_0__0_.mux_right_track_0.out VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_10.mux_l1_in_0_ net17 net69 sb_0__0_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_29_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_30.out sky130_fd_sc_hd__clkbuf_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_8.mux_l1_in_0_ net18 net68 sb_0__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput124 net124 VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_12
Xoutput102 net102 VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_12
XFILLER_87_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_30.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_32.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput37 chany_top_in[14] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput26 chanx_right_in[4] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 chanx_right_in[21] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xinput59 chany_top_in[7] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
Xinput48 chany_top_in[24] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_18.out sky130_fd_sc_hd__clkbuf_1
XFILLER_83_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_100_ sb_0__0_.mux_right_track_2.out VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_8.mux_l2_in_0__158 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_8.mux_l2_in_0__158/HI
+ net158 sky130_fd_sc_hd__conb_1
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_7__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_7__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_right_track_18.mux_l1_in_0_ net66 net45 sb_0__0_.mem_right_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_32.mux_l2_in_0_ net132 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_32.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_8.mux_l2_in_0__140 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_8.mux_l2_in_0__140/HI
+ net140 sky130_fd_sc_hd__conb_1
XFILLER_50_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_top_track_34.mux_l2_in_0_ net151 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_34.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput114 net114 VGND VGND VPWR VPWR chany_top_out[20] sky130_fd_sc_hd__buf_12
Xoutput103 net103 VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_12
Xoutput125 net125 VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_12
XFILLER_87_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput27 chanx_right_in[5] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput16 chanx_right_in[22] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput49 chany_top_in[25] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput38 chany_top_in[15] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_6__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_6__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_46.out sky130_fd_sc_hd__clkbuf_1
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_12_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_10.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_10.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_50.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_0.ccff_head sky130_fd_sc_hd__dfrtp_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_48.mux_l2_in_0__155 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_48.mux_l2_in_0__155/HI
+ net155 sky130_fd_sc_hd__conb_1
XFILLER_67_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_32.mux_l1_in_0_ net65 net37 sb_0__0_.mem_right_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_5__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_44.mux_l2_in_0_ net135 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_44.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput115 net115 VGND VGND VPWR VPWR chany_top_out[21] sky130_fd_sc_hd__buf_12
Xoutput104 net104 VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_12
Xoutput126 net126 VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk
+ sb_0__0_.mem_right_track_48.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_48.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput28 chanx_right_in[6] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput17 chanx_right_in[23] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput39 chany_top_in[16] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_34.mux_l1_in_0_ net4 net70 sb_0__0_.mem_top_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_19_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_089_ net41 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_0__0_.mux_top_track_46.mux_l2_in_0_ net154 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_46.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_92_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_10.ccff_head net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_10.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_34.out sky130_fd_sc_hd__clkbuf_1
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_48.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_50.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_4__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_16.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_16.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput116 net116 VGND VGND VPWR VPWR chany_top_out[22] sky130_fd_sc_hd__buf_12
Xoutput105 net105 VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_12
XFILLER_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput127 net127 VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_12
Xsb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_46.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_48.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_4.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_4.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput18 chanx_right_in[24] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 chanx_right_in[7] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_44.mux_l1_in_0_ net63 net60 sb_0__0_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_088_ net40 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_3__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_3__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_46.mux_l1_in_0_ net27 net68 sb_0__0_.mem_top_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk
+ sb_0__0_.mem_right_track_14.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_16.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_6.mux_l1_in_1__157 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_6.mux_l1_in_1__157/HI
+ net157 sky130_fd_sc_hd__conb_1
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput106 net106 VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_12
Xoutput117 net117 VGND VGND VPWR VPWR chany_top_out[23] sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_5__leaf_prog_clk
+ sb_0__0_.mem_right_track_2.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_4.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_32.mux_l2_in_0__150 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_32.mux_l2_in_0__150/HI
+ net150 sky130_fd_sc_hd__conb_1
XFILLER_52_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput19 chanx_right_in[25] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_087_ sb_0__0_.mux_right_track_28.out VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_2__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_top_track_16.mux_l2_in_0__145 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_16.mux_l2_in_0__145/HI
+ net145 sky130_fd_sc_hd__conb_1
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_6.mux_l2_in_0_ sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_0__0_.mem_right_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput107 net107 VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_12
Xoutput129 net129 VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_12
Xoutput118 net118 VGND VGND VPWR VPWR chany_top_out[24] sky130_fd_sc_hd__buf_12
XFILLER_95_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_6.mux_l1_in_1_ net139 net66 sb_0__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_31_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_1__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_1__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_4.mux_l2_in_0_ net152 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_4.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_086_ sb_0__0_.mux_right_track_30.out VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_2
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_2__leaf_prog_clk
+ sb_0__0_.mem_right_track_34.mem_out\[0\] net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_34.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_14.mux_l2_in_0_ net162 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_14.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_3_0__leaf_prog_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_82_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput119 net119 VGND VGND VPWR VPWR chany_top_out[25] sky130_fd_sc_hd__buf_12
Xoutput108 net108 VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_12
XFILLER_95_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput90 net90 VGND VGND VPWR VPWR chanx_right_out[26] sky130_fd_sc_hd__buf_12
XFILLER_68_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_right_track_6.mux_l1_in_0_ net63 net51 sb_0__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_23_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_top_track_16.mux_l2_in_0_ net145 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_16.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_085_ sb_0__0_.mux_right_track_32.out VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_8.out sky130_fd_sc_hd__clkbuf_1
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_4.mux_l1_in_0_ net20 net69 sb_0__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_6__leaf_prog_clk
+ sb_0__0_.mem_right_track_32.ccff_tail net62 VGND VGND VPWR VPWR sb_0__0_.mem_right_track_34.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_14.out sky130_fd_sc_hd__clkbuf_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput109 net109 VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_12
Xoutput80 net80 VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_12
Xoutput91 net91 VGND VGND VPWR VPWR chanx_right_out[27] sky130_fd_sc_hd__buf_12
XFILLER_95_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_14.mux_l1_in_0_ net64 net47 sb_0__0_.mem_right_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_4__leaf_prog_clk sb_0__0_.mem_top_track_4.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_084_ sb_0__0_.mux_right_track_34.out VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_7__leaf_prog_clk sb_0__0_.mem_top_track_10.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_24_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_16.mux_l1_in_0_ net14 net69 sb_0__0_.mem_top_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_21_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_28.mux_l2_in_0_ net148 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_28.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_119_ net9 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xsb_0__0_.mux_top_track_30.mux_l2_in_0_ net149 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_top_track_30.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_46.mux_l2_in_0__154 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_46.mux_l2_in_0__154/HI
+ net154 sky130_fd_sc_hd__conb_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_468 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_8.out sky130_fd_sc_hd__clkbuf_1
XFILLER_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_48.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_48.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput81 net81 VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_12
Xoutput92 net92 VGND VGND VPWR VPWR chanx_right_out[28] sky130_fd_sc_hd__buf_12
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_2.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_68_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_4.mux_l2_in_0__152 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_4.mux_l2_in_0__152/HI
+ net152 sky130_fd_sc_hd__conb_1
X_083_ net35 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_7__leaf_prog_clk sb_0__0_.mem_top_track_10.ccff_head
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mux_top_track_50.mux_l2_in_0__156 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_50.mux_l2_in_0__156/HI
+ net156 sky130_fd_sc_hd__conb_1
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_118_ net8 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_3__leaf_prog_clk sb_0__0_.mem_top_track_16.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_16.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_top_track_28.mux_l1_in_0_ net7 net67 sb_0__0_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_top_track_30.mux_l1_in_0_ net6 net68 sb_0__0_.mem_top_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_0__leaf_prog_clk sb_0__0_.mem_top_track_46.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_48.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput71 net71 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xoutput82 net82 VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_12
Xoutput93 net93 VGND VGND VPWR VPWR chanx_right_out[29] sky130_fd_sc_hd__buf_12
XFILLER_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_30.out sky130_fd_sc_hd__clkbuf_1
XFILLER_77_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_082_ net34 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_18.out sky130_fd_sc_hd__clkbuf_1
XFILLER_11_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_117_ sb_0__0_.mux_top_track_28.out VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_3_1__leaf_prog_clk sb_0__0_.mem_top_track_14.ccff_tail
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_16.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_48_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_2 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput94 net94 VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_12
Xoutput72 net72 VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_12
Xoutput83 net83 VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_12
XFILLER_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_081_ net33 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_top_track_14.mux_l2_in_0__144 VGND VGND VPWR VPWR sb_0__0_.mux_top_track_14.mux_l2_in_0__144/HI
+ net144 sky130_fd_sc_hd__conb_1
Xsb_0__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_ sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_46.out sky130_fd_sc_hd__clkbuf_1
XFILLER_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_116_ sb_0__0_.mux_top_track_30.out VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_0__0_.mux_right_track_18.mux_l2_in_0__164 VGND VGND VPWR VPWR sb_0__0_.mux_right_track_18.mux_l2_in_0__164/HI
+ net164 sky130_fd_sc_hd__conb_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput73 net73 VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_12
Xoutput84 net84 VGND VGND VPWR VPWR chanx_right_out[20] sky130_fd_sc_hd__buf_12
Xoutput95 net95 VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_12
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_080_ net61 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mux_right_track_2.mux_l2_in_0_ net165 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
+ sb_0__0_.mem_right_track_2.ccff_tail VGND VGND VPWR VPWR sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_3_2__leaf_prog_clk sb_0__0_.mem_top_track_34.mem_out\[0\]
+ net62 VGND VGND VPWR VPWR sb_0__0_.mem_top_track_34.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ sb_0__0_.mux_top_track_32.out VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_4 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_0__0_.mux_top_track_0.mux_l2_in_0_ sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_0__0_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput74 net74 VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_12
Xoutput85 net85 VGND VGND VPWR VPWR chanx_right_out[21] sky130_fd_sc_hd__buf_12
Xoutput96 net96 VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_12
XFILLER_48_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
.ends

