magic
tech sky130A
magscale 1 2
timestamp 1656945746
<< viali >>
rect 21189 20553 21223 20587
rect 15853 20485 15887 20519
rect 17233 20485 17267 20519
rect 16129 20417 16163 20451
rect 17765 20417 17799 20451
rect 20462 20417 20496 20451
rect 21005 20417 21039 20451
rect 17509 20349 17543 20383
rect 20729 20349 20763 20383
rect 18889 20213 18923 20247
rect 19349 20213 19383 20247
rect 6561 20009 6595 20043
rect 19257 20009 19291 20043
rect 5181 19941 5215 19975
rect 11437 19873 11471 19907
rect 4261 19805 4295 19839
rect 5365 19805 5399 19839
rect 6193 19805 6227 19839
rect 6745 19805 6779 19839
rect 9321 19805 9355 19839
rect 9597 19805 9631 19839
rect 9873 19805 9907 19839
rect 11713 19805 11747 19839
rect 15485 19805 15519 19839
rect 16037 19805 16071 19839
rect 18061 19805 18095 19839
rect 18889 19805 18923 19839
rect 20637 19805 20671 19839
rect 20913 19805 20947 19839
rect 5917 19737 5951 19771
rect 10149 19737 10183 19771
rect 15240 19737 15274 19771
rect 16304 19737 16338 19771
rect 20370 19737 20404 19771
rect 4077 19669 4111 19703
rect 14105 19669 14139 19703
rect 17417 19669 17451 19703
rect 21097 19669 21131 19703
rect 10425 19465 10459 19499
rect 11529 19465 11563 19499
rect 15761 19465 15795 19499
rect 16221 19465 16255 19499
rect 18337 19465 18371 19499
rect 19993 19465 20027 19499
rect 9965 19397 9999 19431
rect 11989 19397 12023 19431
rect 13860 19397 13894 19431
rect 10057 19329 10091 19363
rect 10701 19329 10735 19363
rect 10977 19329 11011 19363
rect 11897 19329 11931 19363
rect 14648 19329 14682 19363
rect 16037 19329 16071 19363
rect 16948 19329 16982 19363
rect 19450 19329 19484 19363
rect 19717 19329 19751 19363
rect 21106 19329 21140 19363
rect 21373 19329 21407 19363
rect 9873 19261 9907 19295
rect 12173 19261 12207 19295
rect 14105 19261 14139 19295
rect 14381 19261 14415 19295
rect 16681 19261 16715 19295
rect 12725 19125 12759 19159
rect 18061 19125 18095 19159
rect 10057 18785 10091 18819
rect 11253 18785 11287 18819
rect 12357 18717 12391 18751
rect 12613 18717 12647 18751
rect 14105 18717 14139 18751
rect 15761 18717 15795 18751
rect 18797 18717 18831 18751
rect 19257 18717 19291 18751
rect 14350 18649 14384 18683
rect 16006 18649 16040 18683
rect 18530 18649 18564 18683
rect 19502 18649 19536 18683
rect 13737 18581 13771 18615
rect 15485 18581 15519 18615
rect 17141 18581 17175 18615
rect 17417 18581 17451 18615
rect 20637 18581 20671 18615
rect 13952 18309 13986 18343
rect 14197 18241 14231 18275
rect 17417 18241 17451 18275
rect 17673 18241 17707 18275
rect 20462 18241 20496 18275
rect 20729 18241 20763 18275
rect 12817 18037 12851 18071
rect 18797 18037 18831 18071
rect 19349 18037 19383 18071
rect 16405 17833 16439 17867
rect 17785 17697 17819 17731
rect 17518 17629 17552 17663
rect 19901 17629 19935 17663
rect 18153 17561 18187 17595
rect 20146 17561 20180 17595
rect 21281 17493 21315 17527
rect 11529 17289 11563 17323
rect 14013 17289 14047 17323
rect 17693 17289 17727 17323
rect 19533 17289 19567 17323
rect 14556 17221 14590 17255
rect 18806 17221 18840 17255
rect 11897 17153 11931 17187
rect 12633 17153 12667 17187
rect 12900 17153 12934 17187
rect 14289 17153 14323 17187
rect 19073 17153 19107 17187
rect 21025 17153 21059 17187
rect 21281 17153 21315 17187
rect 11989 17085 12023 17119
rect 12173 17085 12207 17119
rect 15669 16949 15703 16983
rect 19901 16949 19935 16983
rect 19349 16745 19383 16779
rect 11897 16609 11931 16643
rect 12357 16609 12391 16643
rect 17233 16609 17267 16643
rect 15117 16541 15151 16575
rect 17500 16541 17534 16575
rect 19901 16541 19935 16575
rect 20157 16541 20191 16575
rect 12624 16473 12658 16507
rect 15384 16473 15418 16507
rect 13737 16405 13771 16439
rect 16497 16405 16531 16439
rect 18613 16405 18647 16439
rect 21281 16405 21315 16439
rect 9873 16201 9907 16235
rect 10333 16201 10367 16235
rect 15761 16201 15795 16235
rect 17816 16133 17850 16167
rect 10241 16065 10275 16099
rect 10885 16065 10919 16099
rect 12725 16065 12759 16099
rect 12992 16065 13026 16099
rect 14381 16065 14415 16099
rect 14648 16065 14682 16099
rect 20076 16065 20110 16099
rect 10517 15997 10551 16031
rect 18061 15997 18095 16031
rect 19809 15997 19843 16031
rect 14105 15861 14139 15895
rect 16681 15861 16715 15895
rect 21189 15861 21223 15895
rect 16497 15521 16531 15555
rect 19533 15453 19567 15487
rect 19789 15453 19823 15487
rect 16230 15385 16264 15419
rect 15117 15317 15151 15351
rect 20913 15317 20947 15351
rect 10149 15113 10183 15147
rect 10517 14977 10551 15011
rect 10609 14977 10643 15011
rect 14114 14977 14148 15011
rect 14381 14977 14415 15011
rect 20565 14977 20599 15011
rect 10793 14909 10827 14943
rect 20821 14909 20855 14943
rect 13001 14773 13035 14807
rect 19441 14773 19475 14807
rect 10241 14569 10275 14603
rect 16313 14501 16347 14535
rect 9689 14433 9723 14467
rect 10517 14433 10551 14467
rect 15485 14433 15519 14467
rect 12357 14365 12391 14399
rect 17693 14365 17727 14399
rect 20637 14365 20671 14399
rect 9873 14297 9907 14331
rect 12624 14297 12658 14331
rect 15218 14297 15252 14331
rect 17448 14297 17482 14331
rect 20370 14297 20404 14331
rect 9229 14229 9263 14263
rect 9781 14229 9815 14263
rect 11069 14229 11103 14263
rect 13737 14229 13771 14263
rect 14105 14229 14139 14263
rect 19257 14229 19291 14263
rect 12449 14025 12483 14059
rect 14105 14025 14139 14059
rect 18061 14025 18095 14059
rect 19993 14025 20027 14059
rect 16948 13957 16982 13991
rect 13573 13889 13607 13923
rect 13829 13889 13863 13923
rect 15218 13889 15252 13923
rect 15485 13889 15519 13923
rect 16681 13889 16715 13923
rect 18337 13889 18371 13923
rect 18604 13889 18638 13923
rect 21117 13889 21151 13923
rect 21373 13821 21407 13855
rect 19717 13685 19751 13719
rect 14289 13481 14323 13515
rect 21097 13481 21131 13515
rect 16773 13413 16807 13447
rect 15669 13345 15703 13379
rect 18153 13345 18187 13379
rect 19257 13345 19291 13379
rect 17886 13277 17920 13311
rect 20913 13277 20947 13311
rect 15402 13209 15436 13243
rect 19524 13209 19558 13243
rect 20637 13141 20671 13175
rect 11897 12937 11931 12971
rect 12725 12937 12759 12971
rect 14749 12937 14783 12971
rect 17233 12937 17267 12971
rect 19993 12937 20027 12971
rect 21106 12869 21140 12903
rect 11989 12801 12023 12835
rect 13001 12801 13035 12835
rect 13268 12801 13302 12835
rect 15862 12801 15896 12835
rect 16129 12801 16163 12835
rect 18346 12801 18380 12835
rect 18613 12801 18647 12835
rect 21373 12801 21407 12835
rect 11805 12733 11839 12767
rect 11069 12665 11103 12699
rect 12357 12597 12391 12631
rect 14381 12597 14415 12631
rect 18705 12393 18739 12427
rect 19993 12393 20027 12427
rect 20545 12393 20579 12427
rect 21097 12393 21131 12427
rect 14841 12325 14875 12359
rect 16497 12325 16531 12359
rect 14197 12257 14231 12291
rect 15853 12257 15887 12291
rect 17325 12257 17359 12291
rect 17049 12189 17083 12223
rect 17785 12189 17819 12223
rect 18521 12189 18555 12223
rect 19809 12189 19843 12223
rect 20361 12189 20395 12223
rect 20913 12189 20947 12223
rect 18061 12121 18095 12155
rect 14381 12053 14415 12087
rect 14473 12053 14507 12087
rect 15485 12053 15519 12087
rect 16037 12053 16071 12087
rect 16129 12053 16163 12087
rect 12817 11849 12851 11883
rect 13277 11849 13311 11883
rect 14197 11849 14231 11883
rect 15577 11849 15611 11883
rect 16681 11849 16715 11883
rect 17141 11849 17175 11883
rect 18521 11849 18555 11883
rect 21005 11849 21039 11883
rect 12909 11713 12943 11747
rect 13553 11713 13587 11747
rect 14473 11713 14507 11747
rect 17509 11713 17543 11747
rect 18337 11713 18371 11747
rect 18889 11713 18923 11747
rect 19625 11713 19659 11747
rect 20821 11713 20855 11747
rect 12725 11645 12759 11679
rect 14749 11645 14783 11679
rect 15301 11645 15335 11679
rect 15485 11645 15519 11679
rect 17601 11645 17635 11679
rect 17693 11645 17727 11679
rect 19165 11645 19199 11679
rect 19901 11645 19935 11679
rect 15945 11577 15979 11611
rect 16313 11509 16347 11543
rect 12173 11305 12207 11339
rect 12449 11305 12483 11339
rect 14841 11305 14875 11339
rect 15393 11305 15427 11339
rect 19441 11305 19475 11339
rect 21005 11305 21039 11339
rect 18889 11237 18923 11271
rect 11621 11169 11655 11203
rect 13093 11169 13127 11203
rect 14289 11169 14323 11203
rect 15945 11169 15979 11203
rect 17509 11169 17543 11203
rect 17969 11169 18003 11203
rect 14381 11101 14415 11135
rect 19257 11101 19291 11135
rect 20821 11101 20855 11135
rect 11069 11033 11103 11067
rect 11805 11033 11839 11067
rect 12909 11033 12943 11067
rect 13737 11033 13771 11067
rect 14473 11033 14507 11067
rect 15853 11033 15887 11067
rect 16589 11033 16623 11067
rect 17325 11033 17359 11067
rect 17417 11033 17451 11067
rect 19809 11033 19843 11067
rect 20269 11033 20303 11067
rect 11713 10965 11747 10999
rect 12817 10965 12851 10999
rect 15761 10965 15795 10999
rect 16957 10965 16991 10999
rect 18521 10965 18555 10999
rect 13737 10761 13771 10795
rect 16681 10761 16715 10795
rect 17141 10761 17175 10795
rect 17693 10761 17727 10795
rect 20177 10761 20211 10795
rect 21005 10761 21039 10795
rect 12357 10693 12391 10727
rect 13369 10693 13403 10727
rect 17049 10693 17083 10727
rect 18061 10693 18095 10727
rect 19165 10693 19199 10727
rect 14105 10625 14139 10659
rect 14749 10625 14783 10659
rect 15853 10625 15887 10659
rect 16129 10625 16163 10659
rect 19073 10625 19107 10659
rect 20085 10625 20119 10659
rect 20821 10625 20855 10659
rect 12725 10557 12759 10591
rect 14197 10557 14231 10591
rect 14289 10557 14323 10591
rect 15025 10557 15059 10591
rect 17233 10557 17267 10591
rect 18153 10557 18187 10591
rect 18337 10557 18371 10591
rect 19257 10557 19291 10591
rect 20269 10557 20303 10591
rect 15485 10421 15519 10455
rect 18705 10421 18739 10455
rect 19717 10421 19751 10455
rect 13645 10217 13679 10251
rect 14841 10217 14875 10251
rect 15945 10217 15979 10251
rect 20453 10217 20487 10251
rect 21005 10217 21039 10251
rect 12449 10149 12483 10183
rect 13093 10081 13127 10115
rect 14289 10081 14323 10115
rect 16497 10081 16531 10115
rect 17509 10081 17543 10115
rect 17693 10081 17727 10115
rect 19533 10081 19567 10115
rect 19257 10013 19291 10047
rect 20821 10013 20855 10047
rect 12817 9945 12851 9979
rect 15577 9945 15611 9979
rect 17417 9945 17451 9979
rect 18061 9945 18095 9979
rect 12081 9877 12115 9911
rect 12909 9877 12943 9911
rect 14381 9877 14415 9911
rect 14473 9877 14507 9911
rect 15117 9877 15151 9911
rect 16313 9877 16347 9911
rect 16405 9877 16439 9911
rect 17049 9877 17083 9911
rect 18521 9877 18555 9911
rect 19993 9877 20027 9911
rect 14381 9673 14415 9707
rect 12357 9605 12391 9639
rect 16681 9605 16715 9639
rect 18245 9605 18279 9639
rect 20821 9605 20855 9639
rect 21373 9605 21407 9639
rect 12449 9537 12483 9571
rect 14473 9537 14507 9571
rect 17969 9537 18003 9571
rect 19073 9537 19107 9571
rect 19717 9537 19751 9571
rect 20545 9537 20579 9571
rect 12265 9469 12299 9503
rect 14289 9469 14323 9503
rect 15117 9469 15151 9503
rect 15577 9469 15611 9503
rect 19809 9469 19843 9503
rect 19901 9469 19935 9503
rect 12817 9401 12851 9435
rect 14841 9401 14875 9435
rect 19349 9401 19383 9435
rect 11713 9333 11747 9367
rect 13369 9333 13403 9367
rect 13645 9333 13679 9367
rect 17509 9333 17543 9367
rect 16405 8993 16439 9027
rect 18061 8993 18095 9027
rect 20269 8993 20303 9027
rect 16313 8925 16347 8959
rect 19257 8925 19291 8959
rect 19993 8925 20027 8959
rect 21097 8925 21131 8959
rect 16221 8857 16255 8891
rect 16865 8857 16899 8891
rect 18245 8857 18279 8891
rect 19533 8857 19567 8891
rect 14565 8789 14599 8823
rect 15853 8789 15887 8823
rect 17601 8789 17635 8823
rect 18153 8789 18187 8823
rect 18613 8789 18647 8823
rect 20913 8789 20947 8823
rect 14565 8585 14599 8619
rect 14933 8585 14967 8619
rect 17049 8585 17083 8619
rect 17141 8585 17175 8619
rect 17693 8585 17727 8619
rect 19349 8585 19383 8619
rect 20453 8585 20487 8619
rect 21005 8585 21039 8619
rect 14473 8449 14507 8483
rect 15853 8449 15887 8483
rect 15945 8449 15979 8483
rect 18061 8449 18095 8483
rect 19165 8449 19199 8483
rect 20085 8449 20119 8483
rect 20821 8449 20855 8483
rect 13829 8381 13863 8415
rect 14381 8381 14415 8415
rect 15761 8381 15795 8415
rect 17233 8381 17267 8415
rect 18153 8381 18187 8415
rect 18245 8381 18279 8415
rect 19809 8381 19843 8415
rect 19993 8381 20027 8415
rect 15209 8313 15243 8347
rect 16313 8313 16347 8347
rect 16681 8245 16715 8279
rect 18705 8245 18739 8279
rect 14841 8041 14875 8075
rect 18429 8041 18463 8075
rect 20361 8041 20395 8075
rect 14197 7905 14231 7939
rect 15853 7905 15887 7939
rect 17877 7905 17911 7939
rect 19533 7905 19567 7939
rect 21005 7905 21039 7939
rect 5825 7837 5859 7871
rect 6101 7837 6135 7871
rect 16773 7837 16807 7871
rect 17049 7837 17083 7871
rect 19257 7837 19291 7871
rect 14473 7769 14507 7803
rect 16497 7769 16531 7803
rect 17969 7769 18003 7803
rect 19993 7769 20027 7803
rect 5641 7701 5675 7735
rect 13645 7701 13679 7735
rect 14381 7701 14415 7735
rect 15209 7701 15243 7735
rect 15577 7701 15611 7735
rect 18061 7701 18095 7735
rect 18705 7701 18739 7735
rect 20729 7701 20763 7735
rect 20821 7701 20855 7735
rect 13645 7497 13679 7531
rect 14105 7497 14139 7531
rect 14749 7497 14783 7531
rect 17325 7497 17359 7531
rect 17785 7497 17819 7531
rect 19073 7497 19107 7531
rect 20085 7497 20119 7531
rect 20637 7497 20671 7531
rect 21097 7497 21131 7531
rect 18705 7429 18739 7463
rect 13369 7361 13403 7395
rect 14013 7361 14047 7395
rect 15669 7361 15703 7395
rect 17693 7361 17727 7395
rect 19717 7361 19751 7395
rect 21005 7361 21039 7395
rect 14289 7293 14323 7327
rect 15393 7293 15427 7327
rect 15577 7293 15611 7327
rect 16681 7293 16715 7327
rect 17877 7293 17911 7327
rect 18429 7293 18463 7327
rect 18613 7293 18647 7327
rect 19533 7293 19567 7327
rect 19625 7293 19659 7327
rect 21281 7293 21315 7327
rect 16037 7225 16071 7259
rect 20637 6953 20671 6987
rect 17509 6885 17543 6919
rect 20269 6885 20303 6919
rect 15025 6817 15059 6851
rect 15485 6817 15519 6851
rect 16313 6817 16347 6851
rect 16957 6817 16991 6851
rect 18337 6817 18371 6851
rect 19441 6817 19475 6851
rect 21281 6817 21315 6851
rect 16129 6749 16163 6783
rect 18245 6749 18279 6783
rect 21005 6749 21039 6783
rect 16221 6681 16255 6715
rect 18153 6681 18187 6715
rect 18797 6681 18831 6715
rect 14657 6613 14691 6647
rect 15761 6613 15795 6647
rect 17049 6613 17083 6647
rect 17141 6613 17175 6647
rect 17785 6613 17819 6647
rect 19533 6613 19567 6647
rect 19625 6613 19659 6647
rect 19993 6613 20027 6647
rect 21097 6613 21131 6647
rect 15853 6409 15887 6443
rect 16313 6409 16347 6443
rect 17417 6409 17451 6443
rect 18429 6409 18463 6443
rect 19257 6409 19291 6443
rect 19993 6409 20027 6443
rect 20545 6409 20579 6443
rect 21005 6409 21039 6443
rect 14749 6273 14783 6307
rect 15945 6273 15979 6307
rect 17049 6273 17083 6307
rect 18061 6273 18095 6307
rect 19901 6273 19935 6307
rect 20913 6273 20947 6307
rect 14473 6205 14507 6239
rect 15761 6205 15795 6239
rect 16865 6205 16899 6239
rect 16957 6205 16991 6239
rect 17785 6205 17819 6239
rect 17969 6205 18003 6239
rect 20085 6205 20119 6239
rect 21189 6205 21223 6239
rect 19533 6137 19567 6171
rect 15301 6069 15335 6103
rect 18797 6069 18831 6103
rect 16221 5865 16255 5899
rect 18889 5865 18923 5899
rect 19533 5865 19567 5899
rect 20545 5865 20579 5899
rect 17785 5797 17819 5831
rect 15669 5729 15703 5763
rect 17233 5729 17267 5763
rect 18337 5729 18371 5763
rect 20177 5729 20211 5763
rect 21189 5729 21223 5763
rect 14565 5661 14599 5695
rect 14289 5593 14323 5627
rect 15853 5593 15887 5627
rect 16497 5593 16531 5627
rect 17417 5593 17451 5627
rect 20913 5593 20947 5627
rect 15209 5525 15243 5559
rect 15761 5525 15795 5559
rect 17325 5525 17359 5559
rect 18429 5525 18463 5559
rect 18521 5525 18555 5559
rect 19901 5525 19935 5559
rect 19993 5525 20027 5559
rect 21005 5525 21039 5559
rect 15577 5321 15611 5355
rect 16313 5321 16347 5355
rect 18245 5321 18279 5355
rect 18705 5321 18739 5355
rect 19533 5321 19567 5355
rect 21005 5321 21039 5355
rect 15209 5253 15243 5287
rect 17877 5253 17911 5287
rect 20269 5253 20303 5287
rect 17141 5185 17175 5219
rect 20821 5185 20855 5219
rect 16865 5117 16899 5151
rect 17693 5117 17727 5151
rect 17785 5117 17819 5151
rect 15945 5049 15979 5083
rect 19165 4981 19199 5015
rect 19901 4981 19935 5015
rect 15761 4777 15795 4811
rect 18153 4777 18187 4811
rect 18797 4777 18831 4811
rect 19349 4777 19383 4811
rect 21005 4777 21039 4811
rect 20453 4709 20487 4743
rect 15117 4641 15151 4675
rect 15301 4641 15335 4675
rect 17601 4641 17635 4675
rect 16129 4573 16163 4607
rect 20637 4573 20671 4607
rect 15393 4505 15427 4539
rect 16405 4505 16439 4539
rect 17785 4505 17819 4539
rect 18521 4505 18555 4539
rect 14657 4437 14691 4471
rect 16957 4437 16991 4471
rect 17693 4437 17727 4471
rect 19625 4437 19659 4471
rect 20085 4437 20119 4471
rect 21373 4437 21407 4471
rect 15945 4233 15979 4267
rect 18153 4165 18187 4199
rect 19441 4097 19475 4131
rect 19993 4097 20027 4131
rect 20545 4097 20579 4131
rect 21097 4097 21131 4131
rect 17417 4029 17451 4063
rect 17969 4029 18003 4063
rect 18061 4029 18095 4063
rect 18521 3961 18555 3995
rect 19257 3961 19291 3995
rect 20361 3961 20395 3995
rect 16773 3893 16807 3927
rect 17141 3893 17175 3927
rect 18889 3893 18923 3927
rect 19809 3893 19843 3927
rect 20913 3893 20947 3927
rect 19349 3689 19383 3723
rect 21189 3689 21223 3723
rect 17969 3621 18003 3655
rect 19901 3621 19935 3655
rect 18705 3553 18739 3587
rect 16681 3485 16715 3519
rect 16957 3485 16991 3519
rect 17325 3485 17359 3519
rect 19533 3485 19567 3519
rect 20085 3485 20119 3519
rect 20913 3485 20947 3519
rect 17509 3349 17543 3383
rect 18337 3349 18371 3383
rect 20729 3349 20763 3383
rect 17325 3145 17359 3179
rect 18061 3145 18095 3179
rect 20269 3145 20303 3179
rect 12909 3009 12943 3043
rect 13461 3009 13495 3043
rect 16037 3009 16071 3043
rect 17693 3009 17727 3043
rect 18429 3009 18463 3043
rect 19349 3009 19383 3043
rect 19901 3009 19935 3043
rect 20453 3009 20487 3043
rect 21097 3009 21131 3043
rect 16957 2941 16991 2975
rect 13277 2873 13311 2907
rect 15853 2873 15887 2907
rect 19717 2873 19751 2907
rect 20913 2873 20947 2907
rect 12725 2805 12759 2839
rect 18797 2805 18831 2839
rect 19165 2805 19199 2839
rect 19625 2601 19659 2635
rect 20913 2601 20947 2635
rect 20361 2533 20395 2567
rect 17417 2465 17451 2499
rect 18521 2397 18555 2431
rect 19809 2397 19843 2431
rect 20545 2397 20579 2431
rect 21097 2397 21131 2431
rect 17785 2329 17819 2363
rect 17049 2261 17083 2295
rect 18153 2261 18187 2295
rect 18889 2261 18923 2295
<< metal1 >>
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 21174 20584 21180 20596
rect 16546 20556 21036 20584
rect 21135 20556 21180 20584
rect 15841 20519 15899 20525
rect 15841 20485 15853 20519
rect 15887 20516 15899 20519
rect 16546 20516 16574 20556
rect 15887 20488 16574 20516
rect 17221 20519 17279 20525
rect 15887 20485 15899 20488
rect 15841 20479 15899 20485
rect 17221 20485 17233 20519
rect 17267 20516 17279 20519
rect 18874 20516 18880 20528
rect 17267 20488 18880 20516
rect 17267 20485 17279 20488
rect 17221 20479 17279 20485
rect 18874 20476 18880 20488
rect 18932 20476 18938 20528
rect 16117 20451 16175 20457
rect 16117 20417 16129 20451
rect 16163 20448 16175 20451
rect 17034 20448 17040 20460
rect 16163 20420 17040 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 17753 20451 17811 20457
rect 17753 20448 17765 20451
rect 17144 20420 17765 20448
rect 16206 20340 16212 20392
rect 16264 20380 16270 20392
rect 17144 20380 17172 20420
rect 17753 20417 17765 20420
rect 17799 20417 17811 20451
rect 17753 20411 17811 20417
rect 19702 20408 19708 20460
rect 19760 20448 19766 20460
rect 21008 20457 21036 20556
rect 21174 20544 21180 20556
rect 21232 20544 21238 20596
rect 20450 20451 20508 20457
rect 20450 20448 20462 20451
rect 19760 20420 20462 20448
rect 19760 20408 19766 20420
rect 20450 20417 20462 20420
rect 20496 20417 20508 20451
rect 20450 20411 20508 20417
rect 20993 20451 21051 20457
rect 20993 20417 21005 20451
rect 21039 20417 21051 20451
rect 20993 20411 21051 20417
rect 17494 20380 17500 20392
rect 16264 20352 17172 20380
rect 17455 20352 17500 20380
rect 16264 20340 16270 20352
rect 17494 20340 17500 20352
rect 17552 20340 17558 20392
rect 20714 20380 20720 20392
rect 20675 20352 20720 20380
rect 20714 20340 20720 20352
rect 20772 20340 20778 20392
rect 18877 20247 18935 20253
rect 18877 20213 18889 20247
rect 18923 20244 18935 20247
rect 18966 20244 18972 20256
rect 18923 20216 18972 20244
rect 18923 20213 18935 20216
rect 18877 20207 18935 20213
rect 18966 20204 18972 20216
rect 19024 20204 19030 20256
rect 19337 20247 19395 20253
rect 19337 20213 19349 20247
rect 19383 20244 19395 20247
rect 19518 20244 19524 20256
rect 19383 20216 19524 20244
rect 19383 20213 19395 20216
rect 19337 20207 19395 20213
rect 19518 20204 19524 20216
rect 19576 20204 19582 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 6546 20040 6552 20052
rect 6507 20012 6552 20040
rect 6546 20000 6552 20012
rect 6604 20000 6610 20052
rect 16206 20000 16212 20052
rect 16264 20040 16270 20052
rect 19245 20043 19303 20049
rect 19245 20040 19257 20043
rect 16264 20012 19257 20040
rect 16264 20000 16270 20012
rect 19245 20009 19257 20012
rect 19291 20009 19303 20043
rect 19245 20003 19303 20009
rect 5166 19972 5172 19984
rect 5127 19944 5172 19972
rect 5166 19932 5172 19944
rect 5224 19932 5230 19984
rect 10962 19972 10968 19984
rect 5368 19944 10968 19972
rect 5368 19845 5396 19944
rect 10962 19932 10968 19944
rect 11020 19932 11026 19984
rect 11425 19907 11483 19913
rect 11425 19904 11437 19907
rect 5552 19876 11437 19904
rect 4249 19839 4307 19845
rect 4249 19805 4261 19839
rect 4295 19805 4307 19839
rect 4249 19799 4307 19805
rect 5353 19839 5411 19845
rect 5353 19805 5365 19839
rect 5399 19805 5411 19839
rect 5353 19799 5411 19805
rect 4264 19768 4292 19799
rect 5552 19768 5580 19876
rect 11425 19873 11437 19876
rect 11471 19873 11483 19907
rect 11425 19867 11483 19873
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19805 6239 19839
rect 6181 19799 6239 19805
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 9309 19839 9367 19845
rect 9309 19836 9321 19839
rect 6779 19808 9321 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 9309 19805 9321 19808
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 9585 19839 9643 19845
rect 9585 19805 9597 19839
rect 9631 19836 9643 19839
rect 9858 19836 9864 19848
rect 9631 19808 9720 19836
rect 9819 19808 9864 19836
rect 9631 19805 9643 19808
rect 9585 19799 9643 19805
rect 5902 19768 5908 19780
rect 4264 19740 5580 19768
rect 5863 19740 5908 19768
rect 5902 19728 5908 19740
rect 5960 19728 5966 19780
rect 6196 19768 6224 19799
rect 6196 19740 6914 19768
rect 4062 19700 4068 19712
rect 4023 19672 4068 19700
rect 4062 19660 4068 19672
rect 4120 19660 4126 19712
rect 6886 19700 6914 19740
rect 9582 19700 9588 19712
rect 6886 19672 9588 19700
rect 9582 19660 9588 19672
rect 9640 19660 9646 19712
rect 9692 19700 9720 19808
rect 9858 19796 9864 19808
rect 9916 19796 9922 19848
rect 11698 19836 11704 19848
rect 11659 19808 11704 19836
rect 11698 19796 11704 19808
rect 11756 19796 11762 19848
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19836 15531 19839
rect 16025 19839 16083 19845
rect 16025 19836 16037 19839
rect 15519 19808 16037 19836
rect 15519 19805 15531 19808
rect 15473 19799 15531 19805
rect 16025 19805 16037 19808
rect 16071 19836 16083 19839
rect 17494 19836 17500 19848
rect 16071 19808 17500 19836
rect 16071 19805 16083 19808
rect 16025 19799 16083 19805
rect 17494 19796 17500 19808
rect 17552 19836 17558 19848
rect 18046 19836 18052 19848
rect 17552 19808 18052 19836
rect 17552 19796 17558 19808
rect 18046 19796 18052 19808
rect 18104 19796 18110 19848
rect 18874 19836 18880 19848
rect 18835 19808 18880 19836
rect 18874 19796 18880 19808
rect 18932 19796 18938 19848
rect 20625 19839 20683 19845
rect 20625 19805 20637 19839
rect 20671 19836 20683 19839
rect 20714 19836 20720 19848
rect 20671 19808 20720 19836
rect 20671 19805 20683 19808
rect 20625 19799 20683 19805
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 20898 19836 20904 19848
rect 20859 19808 20904 19836
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 10137 19771 10195 19777
rect 10137 19737 10149 19771
rect 10183 19768 10195 19771
rect 15102 19768 15108 19780
rect 10183 19740 15108 19768
rect 10183 19737 10195 19740
rect 10137 19731 10195 19737
rect 15102 19728 15108 19740
rect 15160 19728 15166 19780
rect 15286 19777 15292 19780
rect 15228 19771 15292 19777
rect 15228 19737 15240 19771
rect 15274 19737 15292 19771
rect 15228 19731 15292 19737
rect 15286 19728 15292 19731
rect 15344 19728 15350 19780
rect 16292 19771 16350 19777
rect 16292 19737 16304 19771
rect 16338 19768 16350 19771
rect 16390 19768 16396 19780
rect 16338 19740 16396 19768
rect 16338 19737 16350 19740
rect 16292 19731 16350 19737
rect 16390 19728 16396 19740
rect 16448 19728 16454 19780
rect 18322 19768 18328 19780
rect 16546 19740 18328 19768
rect 11238 19700 11244 19712
rect 9692 19672 11244 19700
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 14093 19703 14151 19709
rect 14093 19669 14105 19703
rect 14139 19700 14151 19703
rect 14550 19700 14556 19712
rect 14139 19672 14556 19700
rect 14139 19669 14151 19672
rect 14093 19663 14151 19669
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 14918 19660 14924 19712
rect 14976 19700 14982 19712
rect 16546 19700 16574 19740
rect 18322 19728 18328 19740
rect 18380 19728 18386 19780
rect 20254 19768 20260 19780
rect 19536 19740 20260 19768
rect 14976 19672 16574 19700
rect 17405 19703 17463 19709
rect 14976 19660 14982 19672
rect 17405 19669 17417 19703
rect 17451 19700 17463 19703
rect 19536 19700 19564 19740
rect 20254 19728 20260 19740
rect 20312 19768 20318 19780
rect 20358 19771 20416 19777
rect 20358 19768 20370 19771
rect 20312 19740 20370 19768
rect 20312 19728 20318 19740
rect 20358 19737 20370 19740
rect 20404 19737 20416 19771
rect 20358 19731 20416 19737
rect 17451 19672 19564 19700
rect 17451 19669 17463 19672
rect 17405 19663 17463 19669
rect 20622 19660 20628 19712
rect 20680 19700 20686 19712
rect 21085 19703 21143 19709
rect 21085 19700 21097 19703
rect 20680 19672 21097 19700
rect 20680 19660 20686 19672
rect 21085 19669 21097 19672
rect 21131 19669 21143 19703
rect 21085 19663 21143 19669
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 10134 19496 10140 19508
rect 9732 19468 10140 19496
rect 9732 19456 9738 19468
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 10413 19499 10471 19505
rect 10413 19465 10425 19499
rect 10459 19465 10471 19499
rect 10413 19459 10471 19465
rect 9953 19431 10011 19437
rect 9953 19397 9965 19431
rect 9999 19428 10011 19431
rect 9999 19400 10364 19428
rect 9999 19397 10011 19400
rect 9953 19391 10011 19397
rect 10042 19360 10048 19372
rect 10003 19332 10048 19360
rect 10042 19320 10048 19332
rect 10100 19320 10106 19372
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19261 9919 19295
rect 10336 19292 10364 19400
rect 10428 19360 10456 19459
rect 11238 19456 11244 19508
rect 11296 19496 11302 19508
rect 11517 19499 11575 19505
rect 11517 19496 11529 19499
rect 11296 19468 11529 19496
rect 11296 19456 11302 19468
rect 11517 19465 11529 19468
rect 11563 19465 11575 19499
rect 11517 19459 11575 19465
rect 15749 19499 15807 19505
rect 15749 19465 15761 19499
rect 15795 19496 15807 19499
rect 15838 19496 15844 19508
rect 15795 19468 15844 19496
rect 15795 19465 15807 19468
rect 15749 19459 15807 19465
rect 15838 19456 15844 19468
rect 15896 19456 15902 19508
rect 16209 19499 16267 19505
rect 16209 19465 16221 19499
rect 16255 19496 16267 19499
rect 18138 19496 18144 19508
rect 16255 19468 18144 19496
rect 16255 19465 16267 19468
rect 16209 19459 16267 19465
rect 18138 19456 18144 19468
rect 18196 19456 18202 19508
rect 18322 19496 18328 19508
rect 18283 19468 18328 19496
rect 18322 19456 18328 19468
rect 18380 19456 18386 19508
rect 19702 19456 19708 19508
rect 19760 19496 19766 19508
rect 19981 19499 20039 19505
rect 19981 19496 19993 19499
rect 19760 19468 19993 19496
rect 19760 19456 19766 19468
rect 19981 19465 19993 19468
rect 20027 19465 20039 19499
rect 19981 19459 20039 19465
rect 10502 19388 10508 19440
rect 10560 19428 10566 19440
rect 11977 19431 12035 19437
rect 11977 19428 11989 19431
rect 10560 19400 11989 19428
rect 10560 19388 10566 19400
rect 11977 19397 11989 19400
rect 12023 19397 12035 19431
rect 11977 19391 12035 19397
rect 13848 19431 13906 19437
rect 13848 19397 13860 19431
rect 13894 19428 13906 19431
rect 14366 19428 14372 19440
rect 13894 19400 14372 19428
rect 13894 19397 13906 19400
rect 13848 19391 13906 19397
rect 14366 19388 14372 19400
rect 14424 19428 14430 19440
rect 14918 19428 14924 19440
rect 14424 19400 14924 19428
rect 14424 19388 14430 19400
rect 14918 19388 14924 19400
rect 14976 19388 14982 19440
rect 15856 19428 15884 19456
rect 15856 19400 17080 19428
rect 10689 19363 10747 19369
rect 10689 19360 10701 19363
rect 10428 19332 10701 19360
rect 10689 19329 10701 19332
rect 10735 19329 10747 19363
rect 10962 19360 10968 19372
rect 10923 19332 10968 19360
rect 10689 19323 10747 19329
rect 10962 19320 10968 19332
rect 11020 19320 11026 19372
rect 11882 19360 11888 19372
rect 11072 19332 11744 19360
rect 11843 19332 11888 19360
rect 11072 19292 11100 19332
rect 10336 19264 11100 19292
rect 11716 19292 11744 19332
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 12894 19360 12900 19372
rect 11992 19332 12900 19360
rect 11992 19292 12020 19332
rect 12894 19320 12900 19332
rect 12952 19320 12958 19372
rect 14642 19369 14648 19372
rect 14636 19323 14648 19369
rect 14700 19360 14706 19372
rect 14700 19332 14736 19360
rect 14642 19320 14648 19323
rect 14700 19320 14706 19332
rect 15102 19320 15108 19372
rect 15160 19360 15166 19372
rect 16942 19369 16948 19372
rect 16025 19363 16083 19369
rect 16025 19360 16037 19363
rect 15160 19332 16037 19360
rect 15160 19320 15166 19332
rect 16025 19329 16037 19332
rect 16071 19329 16083 19363
rect 16936 19360 16948 19369
rect 16903 19332 16948 19360
rect 16025 19323 16083 19329
rect 16936 19323 16948 19332
rect 16942 19320 16948 19323
rect 17000 19320 17006 19372
rect 17052 19360 17080 19400
rect 18046 19388 18052 19440
rect 18104 19428 18110 19440
rect 20714 19428 20720 19440
rect 18104 19400 20720 19428
rect 18104 19388 18110 19400
rect 19720 19369 19748 19400
rect 20714 19388 20720 19400
rect 20772 19428 20778 19440
rect 20772 19400 21404 19428
rect 20772 19388 20778 19400
rect 19438 19363 19496 19369
rect 19438 19360 19450 19363
rect 17052 19332 19450 19360
rect 19438 19329 19450 19332
rect 19484 19329 19496 19363
rect 19438 19323 19496 19329
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19329 19763 19363
rect 21082 19360 21088 19372
rect 21140 19369 21146 19372
rect 21376 19369 21404 19400
rect 21052 19332 21088 19360
rect 19705 19323 19763 19329
rect 21082 19320 21088 19332
rect 21140 19323 21152 19369
rect 21361 19363 21419 19369
rect 21361 19329 21373 19363
rect 21407 19329 21419 19363
rect 21361 19323 21419 19329
rect 21140 19320 21146 19323
rect 11716 19264 12020 19292
rect 12161 19295 12219 19301
rect 9861 19255 9919 19261
rect 12161 19261 12173 19295
rect 12207 19292 12219 19295
rect 14093 19295 14151 19301
rect 12207 19264 13124 19292
rect 12207 19261 12219 19264
rect 12161 19255 12219 19261
rect 9876 19224 9904 19255
rect 12434 19224 12440 19236
rect 9876 19196 12440 19224
rect 12434 19184 12440 19196
rect 12492 19184 12498 19236
rect 12526 19116 12532 19168
rect 12584 19156 12590 19168
rect 12713 19159 12771 19165
rect 12713 19156 12725 19159
rect 12584 19128 12725 19156
rect 12584 19116 12590 19128
rect 12713 19125 12725 19128
rect 12759 19125 12771 19159
rect 13096 19156 13124 19264
rect 14093 19261 14105 19295
rect 14139 19292 14151 19295
rect 14274 19292 14280 19304
rect 14139 19264 14280 19292
rect 14139 19261 14151 19264
rect 14093 19255 14151 19261
rect 14274 19252 14280 19264
rect 14332 19292 14338 19304
rect 14369 19295 14427 19301
rect 14369 19292 14381 19295
rect 14332 19264 14381 19292
rect 14332 19252 14338 19264
rect 14369 19261 14381 19264
rect 14415 19261 14427 19295
rect 14369 19255 14427 19261
rect 16574 19252 16580 19304
rect 16632 19292 16638 19304
rect 16669 19295 16727 19301
rect 16669 19292 16681 19295
rect 16632 19264 16681 19292
rect 16632 19252 16638 19264
rect 16669 19261 16681 19264
rect 16715 19261 16727 19295
rect 16669 19255 16727 19261
rect 15378 19156 15384 19168
rect 13096 19128 15384 19156
rect 12713 19119 12771 19125
rect 15378 19116 15384 19128
rect 15436 19116 15442 19168
rect 18049 19159 18107 19165
rect 18049 19125 18061 19159
rect 18095 19156 18107 19159
rect 18230 19156 18236 19168
rect 18095 19128 18236 19156
rect 18095 19125 18107 19128
rect 18049 19119 18107 19125
rect 18230 19116 18236 19128
rect 18288 19116 18294 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 10042 18816 10048 18828
rect 10003 18788 10048 18816
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 11241 18819 11299 18825
rect 11241 18785 11253 18819
rect 11287 18816 11299 18819
rect 11882 18816 11888 18828
rect 11287 18788 11888 18816
rect 11287 18785 11299 18788
rect 11241 18779 11299 18785
rect 11882 18776 11888 18788
rect 11940 18776 11946 18828
rect 12618 18757 12624 18760
rect 12345 18751 12403 18757
rect 12345 18717 12357 18751
rect 12391 18717 12403 18751
rect 12345 18711 12403 18717
rect 12601 18751 12624 18757
rect 12601 18717 12613 18751
rect 12601 18711 12624 18717
rect 12360 18612 12388 18711
rect 12618 18708 12624 18711
rect 12676 18708 12682 18760
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 12728 18720 14105 18748
rect 12728 18612 12756 18720
rect 14093 18717 14105 18720
rect 14139 18748 14151 18751
rect 14182 18748 14188 18760
rect 14139 18720 14188 18748
rect 14139 18717 14151 18720
rect 14093 18711 14151 18717
rect 14182 18708 14188 18720
rect 14240 18748 14246 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 14240 18720 15761 18748
rect 14240 18708 14246 18720
rect 15749 18717 15761 18720
rect 15795 18748 15807 18751
rect 16574 18748 16580 18760
rect 15795 18720 16580 18748
rect 15795 18717 15807 18720
rect 15749 18711 15807 18717
rect 16574 18708 16580 18720
rect 16632 18748 16638 18760
rect 17402 18748 17408 18760
rect 16632 18720 17408 18748
rect 16632 18708 16638 18720
rect 17402 18708 17408 18720
rect 17460 18748 17466 18760
rect 18785 18751 18843 18757
rect 18785 18748 18797 18751
rect 17460 18720 18797 18748
rect 17460 18708 17466 18720
rect 18785 18717 18797 18720
rect 18831 18748 18843 18751
rect 19058 18748 19064 18760
rect 18831 18720 19064 18748
rect 18831 18717 18843 18720
rect 18785 18711 18843 18717
rect 19058 18708 19064 18720
rect 19116 18748 19122 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 19116 18720 19257 18748
rect 19116 18708 19122 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 12802 18640 12808 18692
rect 12860 18680 12866 18692
rect 14338 18683 14396 18689
rect 14338 18680 14350 18683
rect 12860 18652 14350 18680
rect 12860 18640 12866 18652
rect 14338 18649 14350 18652
rect 14384 18649 14396 18683
rect 14338 18643 14396 18649
rect 15194 18640 15200 18692
rect 15252 18680 15258 18692
rect 15994 18683 16052 18689
rect 15994 18680 16006 18683
rect 15252 18652 16006 18680
rect 15252 18640 15258 18652
rect 15994 18649 16006 18652
rect 16040 18649 16052 18683
rect 15994 18643 16052 18649
rect 17678 18640 17684 18692
rect 17736 18680 17742 18692
rect 18518 18683 18576 18689
rect 18518 18680 18530 18683
rect 17736 18652 18530 18680
rect 17736 18640 17742 18652
rect 18518 18649 18530 18652
rect 18564 18649 18576 18683
rect 18518 18643 18576 18649
rect 18690 18640 18696 18692
rect 18748 18680 18754 18692
rect 19490 18683 19548 18689
rect 19490 18680 19502 18683
rect 18748 18652 19502 18680
rect 18748 18640 18754 18652
rect 19490 18649 19502 18652
rect 19536 18649 19548 18683
rect 19490 18643 19548 18649
rect 12360 18584 12756 18612
rect 13725 18615 13783 18621
rect 13725 18581 13737 18615
rect 13771 18612 13783 18615
rect 13814 18612 13820 18624
rect 13771 18584 13820 18612
rect 13771 18581 13783 18584
rect 13725 18575 13783 18581
rect 13814 18572 13820 18584
rect 13872 18572 13878 18624
rect 15286 18572 15292 18624
rect 15344 18612 15350 18624
rect 15473 18615 15531 18621
rect 15473 18612 15485 18615
rect 15344 18584 15485 18612
rect 15344 18572 15350 18584
rect 15473 18581 15485 18584
rect 15519 18581 15531 18615
rect 17126 18612 17132 18624
rect 17087 18584 17132 18612
rect 15473 18575 15531 18581
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 17405 18615 17463 18621
rect 17405 18581 17417 18615
rect 17451 18612 17463 18615
rect 17494 18612 17500 18624
rect 17451 18584 17500 18612
rect 17451 18581 17463 18584
rect 17405 18575 17463 18581
rect 17494 18572 17500 18584
rect 17552 18572 17558 18624
rect 20438 18572 20444 18624
rect 20496 18612 20502 18624
rect 20625 18615 20683 18621
rect 20625 18612 20637 18615
rect 20496 18584 20637 18612
rect 20496 18572 20502 18584
rect 20625 18581 20637 18584
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 13814 18300 13820 18352
rect 13872 18340 13878 18352
rect 13940 18343 13998 18349
rect 13940 18340 13952 18343
rect 13872 18312 13952 18340
rect 13872 18300 13878 18312
rect 13940 18309 13952 18312
rect 13986 18340 13998 18343
rect 14458 18340 14464 18352
rect 13986 18312 14464 18340
rect 13986 18309 13998 18312
rect 13940 18303 13998 18309
rect 14458 18300 14464 18312
rect 14516 18300 14522 18352
rect 14182 18272 14188 18284
rect 14143 18244 14188 18272
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 17402 18272 17408 18284
rect 17363 18244 17408 18272
rect 17402 18232 17408 18244
rect 17460 18232 17466 18284
rect 17661 18275 17719 18281
rect 17661 18272 17673 18275
rect 17503 18244 17673 18272
rect 15378 18164 15384 18216
rect 15436 18204 15442 18216
rect 16298 18204 16304 18216
rect 15436 18176 16304 18204
rect 15436 18164 15442 18176
rect 16298 18164 16304 18176
rect 16356 18204 16362 18216
rect 17503 18204 17531 18244
rect 17661 18241 17673 18244
rect 17707 18241 17719 18275
rect 17661 18235 17719 18241
rect 20438 18232 20444 18284
rect 20496 18281 20502 18284
rect 20496 18272 20508 18281
rect 20714 18272 20720 18284
rect 20496 18244 20541 18272
rect 20675 18244 20720 18272
rect 20496 18235 20508 18244
rect 20496 18232 20502 18235
rect 20714 18232 20720 18244
rect 20772 18232 20778 18284
rect 16356 18176 17531 18204
rect 16356 18164 16362 18176
rect 10594 18028 10600 18080
rect 10652 18068 10658 18080
rect 12802 18068 12808 18080
rect 10652 18040 12808 18068
rect 10652 18028 10658 18040
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 18782 18068 18788 18080
rect 18743 18040 18788 18068
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 19337 18071 19395 18077
rect 19337 18037 19349 18071
rect 19383 18068 19395 18071
rect 19610 18068 19616 18080
rect 19383 18040 19616 18068
rect 19383 18037 19395 18040
rect 19337 18031 19395 18037
rect 19610 18028 19616 18040
rect 19668 18028 19674 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 16390 17864 16396 17876
rect 16351 17836 16396 17864
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 17402 17824 17408 17876
rect 17460 17864 17466 17876
rect 17460 17836 17816 17864
rect 17460 17824 17466 17836
rect 17788 17737 17816 17836
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17728 17831 17731
rect 17954 17728 17960 17740
rect 17819 17700 17960 17728
rect 17819 17697 17831 17700
rect 17773 17691 17831 17697
rect 17954 17688 17960 17700
rect 18012 17688 18018 17740
rect 17494 17620 17500 17672
rect 17552 17669 17558 17672
rect 17552 17660 17564 17669
rect 17552 17632 17597 17660
rect 17552 17623 17564 17632
rect 17552 17620 17558 17623
rect 19518 17620 19524 17672
rect 19576 17660 19582 17672
rect 19889 17663 19947 17669
rect 19889 17660 19901 17663
rect 19576 17632 19901 17660
rect 19576 17620 19582 17632
rect 19889 17629 19901 17632
rect 19935 17660 19947 17663
rect 20714 17660 20720 17672
rect 19935 17632 20720 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 16942 17552 16948 17604
rect 17000 17592 17006 17604
rect 18141 17595 18199 17601
rect 18141 17592 18153 17595
rect 17000 17564 18153 17592
rect 17000 17552 17006 17564
rect 18141 17561 18153 17564
rect 18187 17561 18199 17595
rect 18141 17555 18199 17561
rect 18414 17552 18420 17604
rect 18472 17592 18478 17604
rect 18966 17592 18972 17604
rect 18472 17564 18972 17592
rect 18472 17552 18478 17564
rect 18966 17552 18972 17564
rect 19024 17592 19030 17604
rect 20134 17595 20192 17601
rect 20134 17592 20146 17595
rect 19024 17564 20146 17592
rect 19024 17552 19030 17564
rect 20134 17561 20146 17564
rect 20180 17561 20192 17595
rect 20134 17555 20192 17561
rect 21269 17527 21327 17533
rect 21269 17493 21281 17527
rect 21315 17524 21327 17527
rect 21358 17524 21364 17536
rect 21315 17496 21364 17524
rect 21315 17493 21327 17496
rect 21269 17487 21327 17493
rect 21358 17484 21364 17496
rect 21416 17484 21422 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 11517 17323 11575 17329
rect 11517 17289 11529 17323
rect 11563 17320 11575 17323
rect 11698 17320 11704 17332
rect 11563 17292 11704 17320
rect 11563 17289 11575 17292
rect 11517 17283 11575 17289
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 14001 17323 14059 17329
rect 14001 17289 14013 17323
rect 14047 17320 14059 17323
rect 14642 17320 14648 17332
rect 14047 17292 14648 17320
rect 14047 17289 14059 17292
rect 14001 17283 14059 17289
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 17678 17320 17684 17332
rect 17639 17292 17684 17320
rect 17678 17280 17684 17292
rect 17736 17280 17742 17332
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 19521 17323 19579 17329
rect 19521 17320 19533 17323
rect 19484 17292 19533 17320
rect 19484 17280 19490 17292
rect 19521 17289 19533 17292
rect 19567 17320 19579 17323
rect 19886 17320 19892 17332
rect 19567 17292 19892 17320
rect 19567 17289 19579 17292
rect 19521 17283 19579 17289
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 14550 17261 14556 17264
rect 14544 17252 14556 17261
rect 12636 17224 14320 17252
rect 14511 17224 14556 17252
rect 11882 17184 11888 17196
rect 11843 17156 11888 17184
rect 11882 17144 11888 17156
rect 11940 17144 11946 17196
rect 12342 17144 12348 17196
rect 12400 17184 12406 17196
rect 12636 17193 12664 17224
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 12400 17156 12633 17184
rect 12400 17144 12406 17156
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 12888 17187 12946 17193
rect 12888 17153 12900 17187
rect 12934 17184 12946 17187
rect 13814 17184 13820 17196
rect 12934 17156 13820 17184
rect 12934 17153 12946 17156
rect 12888 17147 12946 17153
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 14292 17193 14320 17224
rect 14544 17215 14556 17224
rect 14550 17212 14556 17215
rect 14608 17212 14614 17264
rect 18322 17212 18328 17264
rect 18380 17252 18386 17264
rect 18782 17252 18788 17264
rect 18840 17261 18846 17264
rect 18380 17224 18788 17252
rect 18380 17212 18386 17224
rect 18782 17212 18788 17224
rect 18840 17252 18852 17261
rect 18840 17224 18885 17252
rect 18840 17215 18852 17224
rect 18840 17212 18846 17215
rect 20714 17212 20720 17264
rect 20772 17252 20778 17264
rect 20772 17224 21312 17252
rect 20772 17212 20778 17224
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17184 14335 17187
rect 14366 17184 14372 17196
rect 14323 17156 14372 17184
rect 14323 17153 14335 17156
rect 14277 17147 14335 17153
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 19058 17184 19064 17196
rect 19019 17156 19064 17184
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 21013 17187 21071 17193
rect 21013 17153 21025 17187
rect 21059 17184 21071 17187
rect 21174 17184 21180 17196
rect 21059 17156 21180 17184
rect 21059 17153 21071 17156
rect 21013 17147 21071 17153
rect 21174 17144 21180 17156
rect 21232 17144 21238 17196
rect 21284 17193 21312 17224
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17153 21327 17187
rect 21269 17147 21327 17153
rect 11974 17116 11980 17128
rect 11935 17088 11980 17116
rect 11974 17076 11980 17088
rect 12032 17076 12038 17128
rect 12161 17119 12219 17125
rect 12161 17085 12173 17119
rect 12207 17116 12219 17119
rect 12207 17088 12664 17116
rect 12207 17085 12219 17088
rect 12161 17079 12219 17085
rect 12636 16980 12664 17088
rect 14550 16980 14556 16992
rect 12636 16952 14556 16980
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 15657 16983 15715 16989
rect 15657 16980 15669 16983
rect 15436 16952 15669 16980
rect 15436 16940 15442 16952
rect 15657 16949 15669 16952
rect 15703 16949 15715 16983
rect 15657 16943 15715 16949
rect 19889 16983 19947 16989
rect 19889 16949 19901 16983
rect 19935 16980 19947 16983
rect 20898 16980 20904 16992
rect 19935 16952 20904 16980
rect 19935 16949 19947 16952
rect 19889 16943 19947 16949
rect 20898 16940 20904 16952
rect 20956 16980 20962 16992
rect 21082 16980 21088 16992
rect 20956 16952 21088 16980
rect 20956 16940 20962 16952
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 17954 16776 17960 16788
rect 17236 16748 17960 16776
rect 11882 16640 11888 16652
rect 11843 16612 11888 16640
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 12342 16640 12348 16652
rect 12303 16612 12348 16640
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 17236 16649 17264 16748
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 18230 16736 18236 16788
rect 18288 16776 18294 16788
rect 19337 16779 19395 16785
rect 19337 16776 19349 16779
rect 18288 16748 19349 16776
rect 18288 16736 18294 16748
rect 19337 16745 19349 16748
rect 19383 16776 19395 16779
rect 22462 16776 22468 16788
rect 19383 16748 22468 16776
rect 19383 16745 19395 16748
rect 19337 16739 19395 16745
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 17221 16643 17279 16649
rect 17221 16640 17233 16643
rect 16500 16612 17233 16640
rect 12434 16532 12440 16584
rect 12492 16572 12498 16584
rect 12492 16544 14320 16572
rect 12492 16532 12498 16544
rect 12612 16507 12670 16513
rect 12612 16473 12624 16507
rect 12658 16504 12670 16507
rect 12710 16504 12716 16516
rect 12658 16476 12716 16504
rect 12658 16473 12670 16476
rect 12612 16467 12670 16473
rect 12710 16464 12716 16476
rect 12768 16464 12774 16516
rect 13725 16439 13783 16445
rect 13725 16405 13737 16439
rect 13771 16436 13783 16439
rect 13814 16436 13820 16448
rect 13771 16408 13820 16436
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 14292 16436 14320 16544
rect 14366 16532 14372 16584
rect 14424 16572 14430 16584
rect 15105 16575 15163 16581
rect 15105 16572 15117 16575
rect 14424 16544 15117 16572
rect 14424 16532 14430 16544
rect 15105 16541 15117 16544
rect 15151 16572 15163 16575
rect 16500 16572 16528 16612
rect 17221 16609 17233 16612
rect 17267 16609 17279 16643
rect 17221 16603 17279 16609
rect 15151 16544 16528 16572
rect 17488 16575 17546 16581
rect 15151 16541 15163 16544
rect 15105 16535 15163 16541
rect 17488 16541 17500 16575
rect 17534 16572 17546 16575
rect 18230 16572 18236 16584
rect 17534 16544 18236 16572
rect 17534 16541 17546 16544
rect 17488 16535 17546 16541
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 19058 16532 19064 16584
rect 19116 16572 19122 16584
rect 19518 16572 19524 16584
rect 19116 16544 19524 16572
rect 19116 16532 19122 16544
rect 19518 16532 19524 16544
rect 19576 16572 19582 16584
rect 19889 16575 19947 16581
rect 19889 16572 19901 16575
rect 19576 16544 19901 16572
rect 19576 16532 19582 16544
rect 19889 16541 19901 16544
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 19978 16532 19984 16584
rect 20036 16572 20042 16584
rect 20145 16575 20203 16581
rect 20145 16572 20157 16575
rect 20036 16544 20157 16572
rect 20036 16532 20042 16544
rect 20145 16541 20157 16544
rect 20191 16541 20203 16575
rect 20145 16535 20203 16541
rect 15378 16513 15384 16516
rect 15372 16504 15384 16513
rect 15339 16476 15384 16504
rect 15372 16467 15384 16476
rect 15378 16464 15384 16467
rect 15436 16464 15442 16516
rect 16942 16464 16948 16516
rect 17000 16504 17006 16516
rect 17000 16476 21312 16504
rect 17000 16464 17006 16476
rect 16114 16436 16120 16448
rect 14292 16408 16120 16436
rect 16114 16396 16120 16408
rect 16172 16436 16178 16448
rect 16485 16439 16543 16445
rect 16485 16436 16497 16439
rect 16172 16408 16497 16436
rect 16172 16396 16178 16408
rect 16485 16405 16497 16408
rect 16531 16405 16543 16439
rect 16485 16399 16543 16405
rect 18601 16439 18659 16445
rect 18601 16405 18613 16439
rect 18647 16436 18659 16439
rect 18690 16436 18696 16448
rect 18647 16408 18696 16436
rect 18647 16405 18659 16408
rect 18601 16399 18659 16405
rect 18690 16396 18696 16408
rect 18748 16396 18754 16448
rect 21284 16445 21312 16476
rect 21269 16439 21327 16445
rect 21269 16405 21281 16439
rect 21315 16405 21327 16439
rect 21269 16399 21327 16405
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 9858 16232 9864 16244
rect 9819 16204 9864 16232
rect 9858 16192 9864 16204
rect 9916 16192 9922 16244
rect 10321 16235 10379 16241
rect 10321 16201 10333 16235
rect 10367 16232 10379 16235
rect 13722 16232 13728 16244
rect 10367 16204 13728 16232
rect 10367 16201 10379 16204
rect 10321 16195 10379 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 14918 16232 14924 16244
rect 13872 16204 14924 16232
rect 13872 16192 13878 16204
rect 14918 16192 14924 16204
rect 14976 16192 14982 16244
rect 15749 16235 15807 16241
rect 15749 16201 15761 16235
rect 15795 16232 15807 16235
rect 16298 16232 16304 16244
rect 15795 16204 16304 16232
rect 15795 16201 15807 16204
rect 15749 16195 15807 16201
rect 16298 16192 16304 16204
rect 16356 16192 16362 16244
rect 12728 16136 14412 16164
rect 12728 16105 12756 16136
rect 14384 16108 14412 16136
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 15562 16164 15568 16176
rect 15344 16136 15568 16164
rect 15344 16124 15350 16136
rect 15562 16124 15568 16136
rect 15620 16124 15626 16176
rect 17804 16167 17862 16173
rect 17804 16133 17816 16167
rect 17850 16164 17862 16167
rect 19518 16164 19524 16176
rect 17850 16136 19524 16164
rect 17850 16133 17862 16136
rect 17804 16127 17862 16133
rect 19518 16124 19524 16136
rect 19576 16124 19582 16176
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16096 10287 16099
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 10275 16068 10885 16096
rect 10275 16065 10287 16068
rect 10229 16059 10287 16065
rect 10873 16065 10885 16068
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 12713 16099 12771 16105
rect 12713 16065 12725 16099
rect 12759 16065 12771 16099
rect 12713 16059 12771 16065
rect 12980 16099 13038 16105
rect 12980 16065 12992 16099
rect 13026 16096 13038 16099
rect 13814 16096 13820 16108
rect 13026 16068 13820 16096
rect 13026 16065 13038 16068
rect 12980 16059 13038 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 14366 16096 14372 16108
rect 14327 16068 14372 16096
rect 14366 16056 14372 16068
rect 14424 16056 14430 16108
rect 14636 16099 14694 16105
rect 14636 16065 14648 16099
rect 14682 16096 14694 16099
rect 15102 16096 15108 16108
rect 14682 16068 15108 16096
rect 14682 16065 14694 16068
rect 14636 16059 14694 16065
rect 15102 16056 15108 16068
rect 15160 16056 15166 16108
rect 17954 16056 17960 16108
rect 18012 16056 18018 16108
rect 20064 16099 20122 16105
rect 20064 16065 20076 16099
rect 20110 16096 20122 16099
rect 20438 16096 20444 16108
rect 20110 16068 20444 16096
rect 20110 16065 20122 16068
rect 20064 16059 20122 16065
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 16028 10563 16031
rect 10594 16028 10600 16040
rect 10551 16000 10600 16028
rect 10551 15997 10563 16000
rect 10505 15991 10563 15997
rect 10594 15988 10600 16000
rect 10652 15988 10658 16040
rect 17972 16028 18000 16056
rect 18049 16031 18107 16037
rect 18049 16028 18061 16031
rect 17972 16000 18061 16028
rect 18049 15997 18061 16000
rect 18095 16028 18107 16031
rect 19058 16028 19064 16040
rect 18095 16000 19064 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 19058 15988 19064 16000
rect 19116 16028 19122 16040
rect 19797 16031 19855 16037
rect 19797 16028 19809 16031
rect 19116 16000 19809 16028
rect 19116 15988 19122 16000
rect 19797 15997 19809 16000
rect 19843 15997 19855 16031
rect 19797 15991 19855 15997
rect 14093 15895 14151 15901
rect 14093 15861 14105 15895
rect 14139 15892 14151 15895
rect 15286 15892 15292 15904
rect 14139 15864 15292 15892
rect 14139 15861 14151 15864
rect 14093 15855 14151 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 15712 15864 16681 15892
rect 15712 15852 15718 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 21174 15892 21180 15904
rect 21087 15864 21180 15892
rect 16669 15855 16727 15861
rect 21174 15852 21180 15864
rect 21232 15892 21238 15904
rect 21542 15892 21548 15904
rect 21232 15864 21548 15892
rect 21232 15852 21238 15864
rect 21542 15852 21548 15864
rect 21600 15852 21606 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15552 16543 15555
rect 17954 15552 17960 15564
rect 16531 15524 17960 15552
rect 16531 15521 16543 15524
rect 16485 15515 16543 15521
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 19058 15444 19064 15496
rect 19116 15484 19122 15496
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 19116 15456 19533 15484
rect 19116 15444 19122 15456
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19610 15444 19616 15496
rect 19668 15484 19674 15496
rect 19777 15487 19835 15493
rect 19777 15484 19789 15487
rect 19668 15456 19789 15484
rect 19668 15444 19674 15456
rect 19777 15453 19789 15456
rect 19823 15453 19835 15487
rect 19777 15447 19835 15453
rect 16114 15376 16120 15428
rect 16172 15416 16178 15428
rect 16218 15419 16276 15425
rect 16218 15416 16230 15419
rect 16172 15388 16230 15416
rect 16172 15376 16178 15388
rect 16218 15385 16230 15388
rect 16264 15385 16276 15419
rect 16218 15379 16276 15385
rect 15102 15348 15108 15360
rect 15063 15320 15108 15348
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 19610 15308 19616 15360
rect 19668 15348 19674 15360
rect 19886 15348 19892 15360
rect 19668 15320 19892 15348
rect 19668 15308 19674 15320
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 20901 15351 20959 15357
rect 20901 15317 20913 15351
rect 20947 15348 20959 15351
rect 21266 15348 21272 15360
rect 20947 15320 21272 15348
rect 20947 15317 20959 15320
rect 20901 15311 20959 15317
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 10134 15144 10140 15156
rect 10095 15116 10140 15144
rect 10134 15104 10140 15116
rect 10192 15104 10198 15156
rect 10502 15008 10508 15020
rect 10463 14980 10508 15008
rect 10502 14968 10508 14980
rect 10560 14968 10566 15020
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 12250 15008 12256 15020
rect 10643 14980 12256 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 12250 14968 12256 14980
rect 12308 14968 12314 15020
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 14102 15011 14160 15017
rect 14102 15008 14114 15011
rect 12492 14980 14114 15008
rect 12492 14968 12498 14980
rect 14102 14977 14114 14980
rect 14148 14977 14160 15011
rect 14366 15008 14372 15020
rect 14327 14980 14372 15008
rect 14102 14971 14160 14977
rect 14366 14968 14372 14980
rect 14424 15008 14430 15020
rect 15470 15008 15476 15020
rect 14424 14980 15476 15008
rect 14424 14968 14430 14980
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 20553 15011 20611 15017
rect 20553 14977 20565 15011
rect 20599 15008 20611 15011
rect 20714 15008 20720 15020
rect 20599 14980 20720 15008
rect 20599 14977 20611 14980
rect 20553 14971 20611 14977
rect 20714 14968 20720 14980
rect 20772 15008 20778 15020
rect 21358 15008 21364 15020
rect 20772 14980 21364 15008
rect 20772 14968 20778 14980
rect 21358 14968 21364 14980
rect 21416 14968 21422 15020
rect 10781 14943 10839 14949
rect 10781 14909 10793 14943
rect 10827 14940 10839 14943
rect 12526 14940 12532 14952
rect 10827 14912 12532 14940
rect 10827 14909 10839 14912
rect 10781 14903 10839 14909
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 20806 14940 20812 14952
rect 20767 14912 20812 14940
rect 20806 14900 20812 14912
rect 20864 14900 20870 14952
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 12989 14807 13047 14813
rect 12989 14804 13001 14807
rect 12768 14776 13001 14804
rect 12768 14764 12774 14776
rect 12989 14773 13001 14776
rect 13035 14773 13047 14807
rect 12989 14767 13047 14773
rect 17862 14764 17868 14816
rect 17920 14804 17926 14816
rect 19429 14807 19487 14813
rect 19429 14804 19441 14807
rect 17920 14776 19441 14804
rect 17920 14764 17926 14776
rect 19429 14773 19441 14776
rect 19475 14773 19487 14807
rect 19429 14767 19487 14773
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 10226 14600 10232 14612
rect 10187 14572 10232 14600
rect 10226 14560 10232 14572
rect 10284 14560 10290 14612
rect 15102 14600 15108 14612
rect 12360 14572 15108 14600
rect 12360 14532 12388 14572
rect 15102 14560 15108 14572
rect 15160 14560 15166 14612
rect 16298 14532 16304 14544
rect 9692 14504 12388 14532
rect 16259 14504 16304 14532
rect 9692 14473 9720 14504
rect 16298 14492 16304 14504
rect 16356 14492 16362 14544
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14433 9735 14467
rect 10502 14464 10508 14476
rect 10463 14436 10508 14464
rect 9677 14427 9735 14433
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 15470 14464 15476 14476
rect 15431 14436 15476 14464
rect 15470 14424 15476 14436
rect 15528 14424 15534 14476
rect 12345 14399 12403 14405
rect 12345 14365 12357 14399
rect 12391 14396 12403 14399
rect 12986 14396 12992 14408
rect 12391 14368 12992 14396
rect 12391 14365 12403 14368
rect 12345 14359 12403 14365
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 16298 14396 16304 14408
rect 14108 14368 16304 14396
rect 9861 14331 9919 14337
rect 9861 14328 9873 14331
rect 9232 14300 9873 14328
rect 9232 14272 9260 14300
rect 9861 14297 9873 14300
rect 9907 14297 9919 14331
rect 9861 14291 9919 14297
rect 12612 14331 12670 14337
rect 12612 14297 12624 14331
rect 12658 14328 12670 14331
rect 14108 14328 14136 14368
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14396 17739 14399
rect 19058 14396 19064 14408
rect 17727 14368 19064 14396
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 19058 14356 19064 14368
rect 19116 14396 19122 14408
rect 20625 14399 20683 14405
rect 20625 14396 20637 14399
rect 19116 14368 20637 14396
rect 19116 14356 19122 14368
rect 20625 14365 20637 14368
rect 20671 14396 20683 14399
rect 20806 14396 20812 14408
rect 20671 14368 20812 14396
rect 20671 14365 20683 14368
rect 20625 14359 20683 14365
rect 20806 14356 20812 14368
rect 20864 14396 20870 14408
rect 21358 14396 21364 14408
rect 20864 14368 21364 14396
rect 20864 14356 20870 14368
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 12658 14300 14136 14328
rect 12658 14297 12670 14300
rect 12612 14291 12670 14297
rect 9214 14260 9220 14272
rect 9175 14232 9220 14260
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 9769 14263 9827 14269
rect 9769 14229 9781 14263
rect 9815 14260 9827 14263
rect 11054 14260 11060 14272
rect 9815 14232 11060 14260
rect 9815 14229 9827 14232
rect 9769 14223 9827 14229
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 14108 14269 14136 14300
rect 15194 14288 15200 14340
rect 15252 14337 15258 14340
rect 15252 14328 15264 14337
rect 15654 14328 15660 14340
rect 15252 14300 15660 14328
rect 15252 14291 15264 14300
rect 15252 14288 15258 14291
rect 15654 14288 15660 14300
rect 15712 14288 15718 14340
rect 17436 14331 17494 14337
rect 17436 14297 17448 14331
rect 17482 14328 17494 14331
rect 17862 14328 17868 14340
rect 17482 14300 17868 14328
rect 17482 14297 17494 14300
rect 17436 14291 17494 14297
rect 17862 14288 17868 14300
rect 17920 14288 17926 14340
rect 18138 14288 18144 14340
rect 18196 14328 18202 14340
rect 20358 14331 20416 14337
rect 20358 14328 20370 14331
rect 18196 14300 20370 14328
rect 18196 14288 18202 14300
rect 20358 14297 20370 14300
rect 20404 14297 20416 14331
rect 20358 14291 20416 14297
rect 13725 14263 13783 14269
rect 13725 14260 13737 14263
rect 13320 14232 13737 14260
rect 13320 14220 13326 14232
rect 13725 14229 13737 14232
rect 13771 14229 13783 14263
rect 13725 14223 13783 14229
rect 14093 14263 14151 14269
rect 14093 14229 14105 14263
rect 14139 14229 14151 14263
rect 14093 14223 14151 14229
rect 18598 14220 18604 14272
rect 18656 14260 18662 14272
rect 19245 14263 19303 14269
rect 19245 14260 19257 14263
rect 18656 14232 19257 14260
rect 18656 14220 18662 14232
rect 19245 14229 19257 14232
rect 19291 14229 19303 14263
rect 19245 14223 19303 14229
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 12434 14056 12440 14068
rect 12395 14028 12440 14056
rect 12434 14016 12440 14028
rect 12492 14016 12498 14068
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 14093 14059 14151 14065
rect 14093 14056 14105 14059
rect 13872 14028 14105 14056
rect 13872 14016 13878 14028
rect 14093 14025 14105 14028
rect 14139 14056 14151 14059
rect 14366 14056 14372 14068
rect 14139 14028 14372 14056
rect 14139 14025 14151 14028
rect 14093 14019 14151 14025
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 14826 14016 14832 14068
rect 14884 14056 14890 14068
rect 17126 14056 17132 14068
rect 14884 14028 17132 14056
rect 14884 14016 14890 14028
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14056 18107 14059
rect 18138 14056 18144 14068
rect 18095 14028 18144 14056
rect 18095 14025 18107 14028
rect 18049 14019 18107 14025
rect 18138 14016 18144 14028
rect 18196 14016 18202 14068
rect 19981 14059 20039 14065
rect 19981 14025 19993 14059
rect 20027 14056 20039 14059
rect 20438 14056 20444 14068
rect 20027 14028 20444 14056
rect 20027 14025 20039 14028
rect 19981 14019 20039 14025
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 12986 13948 12992 14000
rect 13044 13988 13050 14000
rect 16942 13997 16948 14000
rect 16936 13988 16948 13997
rect 13044 13960 15516 13988
rect 16903 13960 16948 13988
rect 13044 13948 13050 13960
rect 13832 13929 13860 13960
rect 15488 13932 15516 13960
rect 16936 13951 16948 13960
rect 16942 13948 16948 13951
rect 17000 13948 17006 14000
rect 19058 13988 19064 14000
rect 18340 13960 19064 13988
rect 13561 13923 13619 13929
rect 13561 13889 13573 13923
rect 13607 13920 13619 13923
rect 13817 13923 13875 13929
rect 13607 13892 13768 13920
rect 13607 13889 13619 13892
rect 13561 13883 13619 13889
rect 13740 13852 13768 13892
rect 13817 13889 13829 13923
rect 13863 13889 13875 13923
rect 13817 13883 13875 13889
rect 14826 13880 14832 13932
rect 14884 13920 14890 13932
rect 15206 13923 15264 13929
rect 15206 13920 15218 13923
rect 14884 13892 15218 13920
rect 14884 13880 14890 13892
rect 15206 13889 15218 13892
rect 15252 13889 15264 13923
rect 15470 13920 15476 13932
rect 15431 13892 15476 13920
rect 15206 13883 15264 13889
rect 15470 13880 15476 13892
rect 15528 13920 15534 13932
rect 15654 13920 15660 13932
rect 15528 13892 15660 13920
rect 15528 13880 15534 13892
rect 15654 13880 15660 13892
rect 15712 13920 15718 13932
rect 18340 13929 18368 13960
rect 19058 13948 19064 13960
rect 19116 13948 19122 14000
rect 18598 13929 18604 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 15712 13892 16681 13920
rect 15712 13880 15718 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 18325 13923 18383 13929
rect 18325 13889 18337 13923
rect 18371 13889 18383 13923
rect 18592 13920 18604 13929
rect 18559 13892 18604 13920
rect 18325 13883 18383 13889
rect 18592 13883 18604 13892
rect 18598 13880 18604 13883
rect 18656 13880 18662 13932
rect 21105 13923 21163 13929
rect 21105 13889 21117 13923
rect 21151 13920 21163 13923
rect 21266 13920 21272 13932
rect 21151 13892 21272 13920
rect 21151 13889 21163 13892
rect 21105 13883 21163 13889
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 21358 13852 21364 13864
rect 13740 13824 13860 13852
rect 21319 13824 21364 13852
rect 13832 13796 13860 13824
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 22002 13812 22008 13864
rect 22060 13852 22066 13864
rect 22554 13852 22560 13864
rect 22060 13824 22560 13852
rect 22060 13812 22066 13824
rect 22554 13812 22560 13824
rect 22612 13812 22618 13864
rect 13814 13744 13820 13796
rect 13872 13744 13878 13796
rect 19702 13716 19708 13728
rect 19663 13688 19708 13716
rect 19702 13676 19708 13688
rect 19760 13676 19766 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14277 13515 14335 13521
rect 14277 13512 14289 13515
rect 13872 13484 14289 13512
rect 13872 13472 13878 13484
rect 14277 13481 14289 13484
rect 14323 13481 14335 13515
rect 14277 13475 14335 13481
rect 14734 13472 14740 13524
rect 14792 13512 14798 13524
rect 21082 13512 21088 13524
rect 14792 13484 16896 13512
rect 21043 13484 21088 13512
rect 14792 13472 14798 13484
rect 16761 13447 16819 13453
rect 16761 13413 16773 13447
rect 16807 13413 16819 13447
rect 16761 13407 16819 13413
rect 15654 13376 15660 13388
rect 15615 13348 15660 13376
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 15194 13200 15200 13252
rect 15252 13240 15258 13252
rect 15390 13243 15448 13249
rect 15390 13240 15402 13243
rect 15252 13212 15402 13240
rect 15252 13200 15258 13212
rect 15390 13209 15402 13212
rect 15436 13240 15448 13243
rect 16776 13240 16804 13407
rect 16868 13308 16896 13484
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 18141 13379 18199 13385
rect 18141 13345 18153 13379
rect 18187 13376 18199 13379
rect 19058 13376 19064 13388
rect 18187 13348 19064 13376
rect 18187 13345 18199 13348
rect 18141 13339 18199 13345
rect 19058 13336 19064 13348
rect 19116 13376 19122 13388
rect 19245 13379 19303 13385
rect 19245 13376 19257 13379
rect 19116 13348 19257 13376
rect 19116 13336 19122 13348
rect 19245 13345 19257 13348
rect 19291 13345 19303 13379
rect 19245 13339 19303 13345
rect 17874 13311 17932 13317
rect 17874 13308 17886 13311
rect 16868 13280 17886 13308
rect 17874 13277 17886 13280
rect 17920 13277 17932 13311
rect 20898 13308 20904 13320
rect 20859 13280 20904 13308
rect 17874 13271 17932 13277
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 15436 13212 16804 13240
rect 15436 13209 15448 13212
rect 15390 13203 15448 13209
rect 17218 13200 17224 13252
rect 17276 13240 17282 13252
rect 19512 13243 19570 13249
rect 17276 13212 19472 13240
rect 17276 13200 17282 13212
rect 12802 13132 12808 13184
rect 12860 13172 12866 13184
rect 17310 13172 17316 13184
rect 12860 13144 17316 13172
rect 12860 13132 12866 13144
rect 17310 13132 17316 13144
rect 17368 13132 17374 13184
rect 19444 13172 19472 13212
rect 19512 13209 19524 13243
rect 19558 13240 19570 13243
rect 19702 13240 19708 13252
rect 19558 13212 19708 13240
rect 19558 13209 19570 13212
rect 19512 13203 19570 13209
rect 19702 13200 19708 13212
rect 19760 13240 19766 13252
rect 20070 13240 20076 13252
rect 19760 13212 20076 13240
rect 19760 13200 19766 13212
rect 20070 13200 20076 13212
rect 20128 13200 20134 13252
rect 20625 13175 20683 13181
rect 20625 13172 20637 13175
rect 19444 13144 20637 13172
rect 20625 13141 20637 13144
rect 20671 13172 20683 13175
rect 21082 13172 21088 13184
rect 20671 13144 21088 13172
rect 20671 13141 20683 13144
rect 20625 13135 20683 13141
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11885 12971 11943 12977
rect 11885 12968 11897 12971
rect 11112 12940 11897 12968
rect 11112 12928 11118 12940
rect 11885 12937 11897 12940
rect 11931 12968 11943 12971
rect 12713 12971 12771 12977
rect 12713 12968 12725 12971
rect 11931 12940 12725 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 12713 12937 12725 12940
rect 12759 12968 12771 12971
rect 12802 12968 12808 12980
rect 12759 12940 12808 12968
rect 12759 12937 12771 12940
rect 12713 12931 12771 12937
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 14550 12928 14556 12980
rect 14608 12968 14614 12980
rect 14734 12968 14740 12980
rect 14608 12940 14740 12968
rect 14608 12928 14614 12940
rect 14734 12928 14740 12940
rect 14792 12928 14798 12980
rect 17221 12971 17279 12977
rect 17221 12968 17233 12971
rect 15580 12940 17233 12968
rect 12434 12900 12440 12912
rect 11808 12872 12440 12900
rect 11808 12773 11836 12872
rect 12434 12860 12440 12872
rect 12492 12860 12498 12912
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12801 12035 12835
rect 12986 12832 12992 12844
rect 12947 12804 12992 12832
rect 11977 12795 12035 12801
rect 11793 12767 11851 12773
rect 11793 12733 11805 12767
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 5534 12656 5540 12708
rect 5592 12696 5598 12708
rect 11057 12699 11115 12705
rect 11057 12696 11069 12699
rect 5592 12668 11069 12696
rect 5592 12656 5598 12668
rect 11057 12665 11069 12668
rect 11103 12696 11115 12699
rect 11992 12696 12020 12795
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13262 12841 13268 12844
rect 13256 12832 13268 12841
rect 13223 12804 13268 12832
rect 13256 12795 13268 12804
rect 13262 12792 13268 12795
rect 13320 12792 13326 12844
rect 13538 12792 13544 12844
rect 13596 12832 13602 12844
rect 15580 12832 15608 12940
rect 17221 12937 17233 12940
rect 17267 12937 17279 12971
rect 17221 12931 17279 12937
rect 19518 12928 19524 12980
rect 19576 12968 19582 12980
rect 19886 12968 19892 12980
rect 19576 12940 19892 12968
rect 19576 12928 19582 12940
rect 19886 12928 19892 12940
rect 19944 12968 19950 12980
rect 19981 12971 20039 12977
rect 19981 12968 19993 12971
rect 19944 12940 19993 12968
rect 19944 12928 19950 12940
rect 19981 12937 19993 12940
rect 20027 12937 20039 12971
rect 19981 12931 20039 12937
rect 15654 12860 15660 12912
rect 15712 12900 15718 12912
rect 15712 12872 16160 12900
rect 15712 12860 15718 12872
rect 16132 12841 16160 12872
rect 21082 12860 21088 12912
rect 21140 12909 21146 12912
rect 21140 12900 21152 12909
rect 21140 12872 21185 12900
rect 21140 12863 21152 12872
rect 21140 12860 21146 12863
rect 15850 12835 15908 12841
rect 15850 12832 15862 12835
rect 13596 12804 15862 12832
rect 13596 12792 13602 12804
rect 15850 12801 15862 12804
rect 15896 12801 15908 12835
rect 15850 12795 15908 12801
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12801 16175 12835
rect 18334 12835 18392 12841
rect 18334 12832 18346 12835
rect 16117 12795 16175 12801
rect 16546 12804 18346 12832
rect 11103 12668 12020 12696
rect 11103 12665 11115 12668
rect 11057 12659 11115 12665
rect 12345 12631 12403 12637
rect 12345 12597 12357 12631
rect 12391 12628 12403 12631
rect 12526 12628 12532 12640
rect 12391 12600 12532 12628
rect 12391 12597 12403 12600
rect 12345 12591 12403 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 14369 12631 14427 12637
rect 14369 12597 14381 12631
rect 14415 12628 14427 12631
rect 15010 12628 15016 12640
rect 14415 12600 15016 12628
rect 14415 12597 14427 12600
rect 14369 12591 14427 12597
rect 15010 12588 15016 12600
rect 15068 12628 15074 12640
rect 16546 12628 16574 12804
rect 18334 12801 18346 12804
rect 18380 12801 18392 12835
rect 18334 12795 18392 12801
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12832 18659 12835
rect 19058 12832 19064 12844
rect 18647 12804 19064 12832
rect 18647 12801 18659 12804
rect 18601 12795 18659 12801
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 21358 12832 21364 12844
rect 21319 12804 21364 12832
rect 21358 12792 21364 12804
rect 21416 12792 21422 12844
rect 15068 12600 16574 12628
rect 15068 12588 15074 12600
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 18690 12424 18696 12436
rect 18651 12396 18696 12424
rect 18690 12384 18696 12396
rect 18748 12384 18754 12436
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20530 12424 20536 12436
rect 20491 12396 20536 12424
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 21085 12427 21143 12433
rect 21085 12393 21097 12427
rect 21131 12424 21143 12427
rect 21450 12424 21456 12436
rect 21131 12396 21456 12424
rect 21131 12393 21143 12396
rect 21085 12387 21143 12393
rect 21450 12384 21456 12396
rect 21508 12384 21514 12436
rect 13906 12316 13912 12368
rect 13964 12356 13970 12368
rect 14366 12356 14372 12368
rect 13964 12328 14372 12356
rect 13964 12316 13970 12328
rect 14366 12316 14372 12328
rect 14424 12316 14430 12368
rect 14829 12359 14887 12365
rect 14829 12325 14841 12359
rect 14875 12325 14887 12359
rect 14829 12319 14887 12325
rect 16485 12359 16543 12365
rect 16485 12325 16497 12359
rect 16531 12356 16543 12359
rect 16531 12328 17264 12356
rect 16531 12325 16543 12328
rect 16485 12319 16543 12325
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 13872 12260 14197 12288
rect 13872 12248 13878 12260
rect 14185 12257 14197 12260
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 14844 12220 14872 12319
rect 15838 12288 15844 12300
rect 15799 12260 15844 12288
rect 15838 12248 15844 12260
rect 15896 12248 15902 12300
rect 17037 12223 17095 12229
rect 17037 12220 17049 12223
rect 14844 12192 17049 12220
rect 17037 12189 17049 12192
rect 17083 12189 17095 12223
rect 17236 12220 17264 12328
rect 17313 12291 17371 12297
rect 17313 12257 17325 12291
rect 17359 12288 17371 12291
rect 17359 12260 20392 12288
rect 17359 12257 17371 12260
rect 17313 12251 17371 12257
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 17236 12192 17785 12220
rect 17037 12183 17095 12189
rect 17773 12189 17785 12192
rect 17819 12189 17831 12223
rect 18509 12223 18567 12229
rect 18509 12220 18521 12223
rect 17773 12183 17831 12189
rect 17880 12192 18521 12220
rect 12158 12044 12164 12096
rect 12216 12084 12222 12096
rect 14369 12087 14427 12093
rect 14369 12084 14381 12087
rect 12216 12056 14381 12084
rect 12216 12044 12222 12056
rect 14369 12053 14381 12056
rect 14415 12053 14427 12087
rect 14369 12047 14427 12053
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 15473 12087 15531 12093
rect 14516 12056 14561 12084
rect 14516 12044 14522 12056
rect 15473 12053 15485 12087
rect 15519 12084 15531 12087
rect 15562 12084 15568 12096
rect 15519 12056 15568 12084
rect 15519 12053 15531 12056
rect 15473 12047 15531 12053
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 15746 12044 15752 12096
rect 15804 12084 15810 12096
rect 16025 12087 16083 12093
rect 16025 12084 16037 12087
rect 15804 12056 16037 12084
rect 15804 12044 15810 12056
rect 16025 12053 16037 12056
rect 16071 12053 16083 12087
rect 16025 12047 16083 12053
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 16172 12056 16217 12084
rect 16172 12044 16178 12056
rect 17126 12044 17132 12096
rect 17184 12084 17190 12096
rect 17880 12084 17908 12192
rect 18509 12189 18521 12192
rect 18555 12189 18567 12223
rect 18509 12183 18567 12189
rect 19518 12180 19524 12232
rect 19576 12220 19582 12232
rect 20364 12229 20392 12260
rect 21266 12248 21272 12300
rect 21324 12288 21330 12300
rect 22186 12288 22192 12300
rect 21324 12260 22192 12288
rect 21324 12248 21330 12260
rect 22186 12248 22192 12260
rect 22244 12248 22250 12300
rect 19797 12223 19855 12229
rect 19797 12220 19809 12223
rect 19576 12192 19809 12220
rect 19576 12180 19582 12192
rect 19797 12189 19809 12192
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 20349 12223 20407 12229
rect 20349 12189 20361 12223
rect 20395 12189 20407 12223
rect 20349 12183 20407 12189
rect 20438 12180 20444 12232
rect 20496 12220 20502 12232
rect 20901 12223 20959 12229
rect 20901 12220 20913 12223
rect 20496 12192 20913 12220
rect 20496 12180 20502 12192
rect 20901 12189 20913 12192
rect 20947 12189 20959 12223
rect 20901 12183 20959 12189
rect 18049 12155 18107 12161
rect 18049 12121 18061 12155
rect 18095 12152 18107 12155
rect 21266 12152 21272 12164
rect 18095 12124 21272 12152
rect 18095 12121 18107 12124
rect 18049 12115 18107 12121
rect 21266 12112 21272 12124
rect 21324 12112 21330 12164
rect 17184 12056 17908 12084
rect 17184 12044 17190 12056
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 12526 11840 12532 11892
rect 12584 11880 12590 11892
rect 12805 11883 12863 11889
rect 12805 11880 12817 11883
rect 12584 11852 12817 11880
rect 12584 11840 12590 11852
rect 12805 11849 12817 11852
rect 12851 11849 12863 11883
rect 12805 11843 12863 11849
rect 13265 11883 13323 11889
rect 13265 11849 13277 11883
rect 13311 11849 13323 11883
rect 13265 11843 13323 11849
rect 14185 11883 14243 11889
rect 14185 11849 14197 11883
rect 14231 11880 14243 11883
rect 14458 11880 14464 11892
rect 14231 11852 14464 11880
rect 14231 11849 14243 11852
rect 14185 11843 14243 11849
rect 13280 11812 13308 11843
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 15562 11880 15568 11892
rect 15523 11852 15568 11880
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 16114 11840 16120 11892
rect 16172 11880 16178 11892
rect 16669 11883 16727 11889
rect 16669 11880 16681 11883
rect 16172 11852 16681 11880
rect 16172 11840 16178 11852
rect 16669 11849 16681 11852
rect 16715 11849 16727 11883
rect 16669 11843 16727 11849
rect 17034 11840 17040 11892
rect 17092 11880 17098 11892
rect 17129 11883 17187 11889
rect 17129 11880 17141 11883
rect 17092 11852 17141 11880
rect 17092 11840 17098 11852
rect 17129 11849 17141 11852
rect 17175 11849 17187 11883
rect 18506 11880 18512 11892
rect 18467 11852 18512 11880
rect 17129 11843 17187 11849
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 20622 11840 20628 11892
rect 20680 11880 20686 11892
rect 20993 11883 21051 11889
rect 20993 11880 21005 11883
rect 20680 11852 21005 11880
rect 20680 11840 20686 11852
rect 20993 11849 21005 11852
rect 21039 11849 21051 11883
rect 20993 11843 21051 11849
rect 13280 11784 19656 11812
rect 12897 11747 12955 11753
rect 12897 11713 12909 11747
rect 12943 11744 12955 11747
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 12943 11716 13553 11744
rect 12943 11713 12955 11716
rect 12897 11707 12955 11713
rect 13541 11713 13553 11716
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 14461 11747 14519 11753
rect 14461 11713 14473 11747
rect 14507 11744 14519 11747
rect 14826 11744 14832 11756
rect 14507 11716 14832 11744
rect 14507 11713 14519 11716
rect 14461 11707 14519 11713
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 17497 11747 17555 11753
rect 17497 11713 17509 11747
rect 17543 11744 17555 11747
rect 17954 11744 17960 11756
rect 17543 11716 17960 11744
rect 17543 11713 17555 11716
rect 17497 11707 17555 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 18046 11704 18052 11756
rect 18104 11744 18110 11756
rect 19628 11753 19656 11784
rect 18325 11747 18383 11753
rect 18325 11744 18337 11747
rect 18104 11716 18337 11744
rect 18104 11704 18110 11716
rect 18325 11713 18337 11716
rect 18371 11713 18383 11747
rect 18325 11707 18383 11713
rect 18877 11747 18935 11753
rect 18877 11713 18889 11747
rect 18923 11713 18935 11747
rect 18877 11707 18935 11713
rect 19613 11747 19671 11753
rect 19613 11713 19625 11747
rect 19659 11713 19671 11747
rect 20806 11744 20812 11756
rect 20767 11716 20812 11744
rect 19613 11707 19671 11713
rect 12710 11676 12716 11688
rect 12671 11648 12716 11676
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 14734 11676 14740 11688
rect 14695 11648 14740 11676
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 15286 11676 15292 11688
rect 15247 11648 15292 11676
rect 15286 11636 15292 11648
rect 15344 11636 15350 11688
rect 15378 11636 15384 11688
rect 15436 11676 15442 11688
rect 15473 11679 15531 11685
rect 15473 11676 15485 11679
rect 15436 11648 15485 11676
rect 15436 11636 15442 11648
rect 15473 11645 15485 11648
rect 15519 11645 15531 11679
rect 17586 11676 17592 11688
rect 17547 11648 17592 11676
rect 15473 11639 15531 11645
rect 17586 11636 17592 11648
rect 17644 11636 17650 11688
rect 17678 11636 17684 11688
rect 17736 11676 17742 11688
rect 17736 11648 17781 11676
rect 17736 11636 17742 11648
rect 15933 11611 15991 11617
rect 15933 11577 15945 11611
rect 15979 11608 15991 11611
rect 18892 11608 18920 11707
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 19153 11679 19211 11685
rect 19153 11645 19165 11679
rect 19199 11645 19211 11679
rect 19153 11639 19211 11645
rect 19889 11679 19947 11685
rect 19889 11645 19901 11679
rect 19935 11676 19947 11679
rect 20714 11676 20720 11688
rect 19935 11648 20720 11676
rect 19935 11645 19947 11648
rect 19889 11639 19947 11645
rect 15979 11580 18920 11608
rect 19168 11608 19196 11639
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 21450 11608 21456 11620
rect 19168 11580 21456 11608
rect 15979 11577 15991 11580
rect 15933 11571 15991 11577
rect 21450 11568 21456 11580
rect 21508 11568 21514 11620
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 15194 11540 15200 11552
rect 11664 11512 15200 11540
rect 11664 11500 11670 11512
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 15838 11500 15844 11552
rect 15896 11540 15902 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 15896 11512 16313 11540
rect 15896 11500 15902 11512
rect 16301 11509 16313 11512
rect 16347 11540 16359 11543
rect 18690 11540 18696 11552
rect 16347 11512 18696 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 12158 11336 12164 11348
rect 12119 11308 12164 11336
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 12437 11339 12495 11345
rect 12437 11305 12449 11339
rect 12483 11336 12495 11339
rect 12894 11336 12900 11348
rect 12483 11308 12900 11336
rect 12483 11305 12495 11308
rect 12437 11299 12495 11305
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 14826 11336 14832 11348
rect 14787 11308 14832 11336
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 15378 11336 15384 11348
rect 15339 11308 15384 11336
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 18782 11296 18788 11348
rect 18840 11336 18846 11348
rect 19429 11339 19487 11345
rect 19429 11336 19441 11339
rect 18840 11308 19441 11336
rect 18840 11296 18846 11308
rect 19429 11305 19441 11308
rect 19475 11305 19487 11339
rect 19429 11299 19487 11305
rect 20993 11339 21051 11345
rect 20993 11305 21005 11339
rect 21039 11336 21051 11339
rect 21174 11336 21180 11348
rect 21039 11308 21180 11336
rect 21039 11305 21051 11308
rect 20993 11299 21051 11305
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 15470 11268 15476 11280
rect 13096 11240 15476 11268
rect 11606 11200 11612 11212
rect 11567 11172 11612 11200
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 13096 11209 13124 11240
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 16942 11228 16948 11280
rect 17000 11268 17006 11280
rect 17402 11268 17408 11280
rect 17000 11240 17408 11268
rect 17000 11228 17006 11240
rect 17402 11228 17408 11240
rect 17460 11228 17466 11280
rect 18874 11268 18880 11280
rect 18835 11240 18880 11268
rect 18874 11228 18880 11240
rect 18932 11228 18938 11280
rect 13081 11203 13139 11209
rect 13081 11169 13093 11203
rect 13127 11169 13139 11203
rect 13081 11163 13139 11169
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11200 14335 11203
rect 14550 11200 14556 11212
rect 14323 11172 14556 11200
rect 14323 11169 14335 11172
rect 14277 11163 14335 11169
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 14918 11160 14924 11212
rect 14976 11200 14982 11212
rect 15933 11203 15991 11209
rect 15933 11200 15945 11203
rect 14976 11172 15945 11200
rect 14976 11160 14982 11172
rect 15933 11169 15945 11172
rect 15979 11169 15991 11203
rect 17494 11200 17500 11212
rect 17455 11172 17500 11200
rect 15933 11163 15991 11169
rect 17494 11160 17500 11172
rect 17552 11160 17558 11212
rect 17954 11200 17960 11212
rect 17915 11172 17960 11200
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 18138 11160 18144 11212
rect 18196 11200 18202 11212
rect 18782 11200 18788 11212
rect 18196 11172 18788 11200
rect 18196 11160 18202 11172
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 12860 11104 14381 11132
rect 12860 11092 12866 11104
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 14734 11092 14740 11144
rect 14792 11132 14798 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 14792 11104 19257 11132
rect 14792 11092 14798 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 20809 11135 20867 11141
rect 20809 11101 20821 11135
rect 20855 11132 20867 11135
rect 20990 11132 20996 11144
rect 20855 11104 20996 11132
rect 20855 11101 20867 11104
rect 20809 11095 20867 11101
rect 20990 11092 20996 11104
rect 21048 11092 21054 11144
rect 6638 11024 6644 11076
rect 6696 11064 6702 11076
rect 11057 11067 11115 11073
rect 11057 11064 11069 11067
rect 6696 11036 11069 11064
rect 6696 11024 6702 11036
rect 11057 11033 11069 11036
rect 11103 11064 11115 11067
rect 11793 11067 11851 11073
rect 11793 11064 11805 11067
rect 11103 11036 11805 11064
rect 11103 11033 11115 11036
rect 11057 11027 11115 11033
rect 11793 11033 11805 11036
rect 11839 11033 11851 11067
rect 11793 11027 11851 11033
rect 12342 11024 12348 11076
rect 12400 11064 12406 11076
rect 12897 11067 12955 11073
rect 12897 11064 12909 11067
rect 12400 11036 12909 11064
rect 12400 11024 12406 11036
rect 12897 11033 12909 11036
rect 12943 11033 12955 11067
rect 12897 11027 12955 11033
rect 13725 11067 13783 11073
rect 13725 11033 13737 11067
rect 13771 11064 13783 11067
rect 14461 11067 14519 11073
rect 14461 11064 14473 11067
rect 13771 11036 14473 11064
rect 13771 11033 13783 11036
rect 13725 11027 13783 11033
rect 14461 11033 14473 11036
rect 14507 11033 14519 11067
rect 15838 11064 15844 11076
rect 15799 11036 15844 11064
rect 14461 11027 14519 11033
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 16577 11067 16635 11073
rect 16577 11033 16589 11067
rect 16623 11064 16635 11067
rect 17034 11064 17040 11076
rect 16623 11036 17040 11064
rect 16623 11033 16635 11036
rect 16577 11027 16635 11033
rect 17034 11024 17040 11036
rect 17092 11024 17098 11076
rect 17313 11067 17371 11073
rect 17313 11033 17325 11067
rect 17359 11033 17371 11067
rect 17313 11027 17371 11033
rect 17405 11067 17463 11073
rect 17405 11033 17417 11067
rect 17451 11064 17463 11067
rect 18874 11064 18880 11076
rect 17451 11036 18880 11064
rect 17451 11033 17463 11036
rect 17405 11027 17463 11033
rect 11701 10999 11759 11005
rect 11701 10965 11713 10999
rect 11747 10996 11759 10999
rect 12360 10996 12388 11024
rect 11747 10968 12388 10996
rect 11747 10965 11759 10968
rect 11701 10959 11759 10965
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 12805 10999 12863 11005
rect 12805 10996 12817 10999
rect 12768 10968 12817 10996
rect 12768 10956 12774 10968
rect 12805 10965 12817 10968
rect 12851 10965 12863 10999
rect 12805 10959 12863 10965
rect 15562 10956 15568 11008
rect 15620 10996 15626 11008
rect 15749 10999 15807 11005
rect 15749 10996 15761 10999
rect 15620 10968 15761 10996
rect 15620 10956 15626 10968
rect 15749 10965 15761 10968
rect 15795 10965 15807 10999
rect 16942 10996 16948 11008
rect 16903 10968 16948 10996
rect 15749 10959 15807 10965
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 17328 10996 17356 11027
rect 18874 11024 18880 11036
rect 18932 11024 18938 11076
rect 19150 11024 19156 11076
rect 19208 11064 19214 11076
rect 19797 11067 19855 11073
rect 19797 11064 19809 11067
rect 19208 11036 19809 11064
rect 19208 11024 19214 11036
rect 19797 11033 19809 11036
rect 19843 11033 19855 11067
rect 19797 11027 19855 11033
rect 20257 11067 20315 11073
rect 20257 11033 20269 11067
rect 20303 11064 20315 11067
rect 20346 11064 20352 11076
rect 20303 11036 20352 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 20346 11024 20352 11036
rect 20404 11024 20410 11076
rect 21082 11024 21088 11076
rect 21140 11064 21146 11076
rect 21450 11064 21456 11076
rect 21140 11036 21456 11064
rect 21140 11024 21146 11036
rect 21450 11024 21456 11036
rect 21508 11024 21514 11076
rect 18506 10996 18512 11008
rect 17328 10968 18512 10996
rect 18506 10956 18512 10968
rect 18564 10956 18570 11008
rect 18690 10956 18696 11008
rect 18748 10996 18754 11008
rect 19168 10996 19196 11024
rect 18748 10968 19196 10996
rect 18748 10956 18754 10968
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 12250 10752 12256 10804
rect 12308 10792 12314 10804
rect 13725 10795 13783 10801
rect 13725 10792 13737 10795
rect 12308 10764 13737 10792
rect 12308 10752 12314 10764
rect 13725 10761 13737 10764
rect 13771 10761 13783 10795
rect 13725 10755 13783 10761
rect 14734 10752 14740 10804
rect 14792 10792 14798 10804
rect 16669 10795 16727 10801
rect 16669 10792 16681 10795
rect 14792 10764 16681 10792
rect 14792 10752 14798 10764
rect 16669 10761 16681 10764
rect 16715 10761 16727 10795
rect 16669 10755 16727 10761
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 17000 10764 17141 10792
rect 17000 10752 17006 10764
rect 17129 10761 17141 10764
rect 17175 10761 17187 10795
rect 17129 10755 17187 10761
rect 17586 10752 17592 10804
rect 17644 10792 17650 10804
rect 17681 10795 17739 10801
rect 17681 10792 17693 10795
rect 17644 10764 17693 10792
rect 17644 10752 17650 10764
rect 17681 10761 17693 10764
rect 17727 10761 17739 10795
rect 20162 10792 20168 10804
rect 20123 10764 20168 10792
rect 17681 10755 17739 10761
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 20993 10795 21051 10801
rect 20993 10761 21005 10795
rect 21039 10792 21051 10795
rect 22094 10792 22100 10804
rect 21039 10764 22100 10792
rect 21039 10761 21051 10764
rect 20993 10755 21051 10761
rect 22094 10752 22100 10764
rect 22152 10752 22158 10804
rect 5810 10684 5816 10736
rect 5868 10724 5874 10736
rect 12342 10724 12348 10736
rect 5868 10696 6914 10724
rect 12255 10696 12348 10724
rect 5868 10684 5874 10696
rect 6886 10656 6914 10696
rect 12342 10684 12348 10696
rect 12400 10724 12406 10736
rect 13357 10727 13415 10733
rect 12400 10696 12664 10724
rect 12400 10684 12406 10696
rect 12434 10656 12440 10668
rect 6886 10628 12440 10656
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 12636 10656 12664 10696
rect 13357 10693 13369 10727
rect 13403 10724 13415 10727
rect 16574 10724 16580 10736
rect 13403 10696 16580 10724
rect 13403 10693 13415 10696
rect 13357 10687 13415 10693
rect 13372 10656 13400 10687
rect 16574 10684 16580 10696
rect 16632 10684 16638 10736
rect 17034 10724 17040 10736
rect 16995 10696 17040 10724
rect 17034 10684 17040 10696
rect 17092 10684 17098 10736
rect 18049 10727 18107 10733
rect 18049 10693 18061 10727
rect 18095 10724 18107 10727
rect 18138 10724 18144 10736
rect 18095 10696 18144 10724
rect 18095 10693 18107 10696
rect 18049 10687 18107 10693
rect 18138 10684 18144 10696
rect 18196 10684 18202 10736
rect 19153 10727 19211 10733
rect 19153 10693 19165 10727
rect 19199 10724 19211 10727
rect 20346 10724 20352 10736
rect 19199 10696 20352 10724
rect 19199 10693 19211 10696
rect 19153 10687 19211 10693
rect 20346 10684 20352 10696
rect 20404 10684 20410 10736
rect 12636 10628 13400 10656
rect 13722 10616 13728 10668
rect 13780 10656 13786 10668
rect 14093 10659 14151 10665
rect 14093 10656 14105 10659
rect 13780 10628 14105 10656
rect 13780 10616 13786 10628
rect 14093 10625 14105 10628
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10656 14795 10659
rect 14826 10656 14832 10668
rect 14783 10628 14832 10656
rect 14783 10625 14795 10628
rect 14737 10619 14795 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 15841 10659 15899 10665
rect 15841 10625 15853 10659
rect 15887 10656 15899 10659
rect 15930 10656 15936 10668
rect 15887 10628 15936 10656
rect 15887 10625 15899 10628
rect 15841 10619 15899 10625
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 16117 10659 16175 10665
rect 16117 10625 16129 10659
rect 16163 10656 16175 10659
rect 17126 10656 17132 10668
rect 16163 10628 17132 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 17126 10616 17132 10628
rect 17184 10616 17190 10668
rect 18506 10616 18512 10668
rect 18564 10656 18570 10668
rect 19061 10659 19119 10665
rect 19061 10656 19073 10659
rect 18564 10628 19073 10656
rect 18564 10616 18570 10628
rect 19061 10625 19073 10628
rect 19107 10656 19119 10659
rect 20073 10659 20131 10665
rect 20073 10656 20085 10659
rect 19107 10628 20085 10656
rect 19107 10625 19119 10628
rect 19061 10619 19119 10625
rect 20073 10625 20085 10628
rect 20119 10625 20131 10659
rect 20073 10619 20131 10625
rect 20714 10616 20720 10668
rect 20772 10656 20778 10668
rect 20809 10659 20867 10665
rect 20809 10656 20821 10659
rect 20772 10628 20821 10656
rect 20772 10616 20778 10628
rect 20809 10625 20821 10628
rect 20855 10625 20867 10659
rect 20809 10619 20867 10625
rect 12710 10588 12716 10600
rect 12671 10560 12716 10588
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10557 14243 10591
rect 14185 10551 14243 10557
rect 14200 10452 14228 10551
rect 14274 10548 14280 10600
rect 14332 10588 14338 10600
rect 15013 10591 15071 10597
rect 14332 10560 14377 10588
rect 14332 10548 14338 10560
rect 15013 10557 15025 10591
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 15028 10520 15056 10551
rect 16390 10548 16396 10600
rect 16448 10588 16454 10600
rect 17221 10591 17279 10597
rect 17221 10588 17233 10591
rect 16448 10560 17233 10588
rect 16448 10548 16454 10560
rect 17221 10557 17233 10560
rect 17267 10557 17279 10591
rect 17221 10551 17279 10557
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18141 10591 18199 10597
rect 18141 10588 18153 10591
rect 18012 10560 18153 10588
rect 18012 10548 18018 10560
rect 18141 10557 18153 10560
rect 18187 10557 18199 10591
rect 18322 10588 18328 10600
rect 18283 10560 18328 10588
rect 18141 10551 18199 10557
rect 18046 10520 18052 10532
rect 15028 10492 18052 10520
rect 18046 10480 18052 10492
rect 18104 10480 18110 10532
rect 18156 10520 18184 10551
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 18414 10548 18420 10600
rect 18472 10588 18478 10600
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 18472 10560 19257 10588
rect 18472 10548 18478 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 20254 10548 20260 10600
rect 20312 10588 20318 10600
rect 20312 10560 20357 10588
rect 20312 10548 20318 10560
rect 19150 10520 19156 10532
rect 18156 10492 19156 10520
rect 19150 10480 19156 10492
rect 19208 10480 19214 10532
rect 15470 10452 15476 10464
rect 14200 10424 15476 10452
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 17494 10412 17500 10464
rect 17552 10452 17558 10464
rect 18693 10455 18751 10461
rect 18693 10452 18705 10455
rect 17552 10424 18705 10452
rect 17552 10412 17558 10424
rect 18693 10421 18705 10424
rect 18739 10421 18751 10455
rect 19702 10452 19708 10464
rect 19663 10424 19708 10452
rect 18693 10415 18751 10421
rect 19702 10412 19708 10424
rect 19760 10412 19766 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 2958 10208 2964 10260
rect 3016 10248 3022 10260
rect 12710 10248 12716 10260
rect 3016 10220 12716 10248
rect 3016 10208 3022 10220
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 13722 10248 13728 10260
rect 13679 10220 13728 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 13722 10208 13728 10220
rect 13780 10208 13786 10260
rect 14826 10248 14832 10260
rect 14787 10220 14832 10248
rect 14826 10208 14832 10220
rect 14884 10208 14890 10260
rect 15930 10248 15936 10260
rect 15891 10220 15936 10248
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16114 10208 16120 10260
rect 16172 10248 16178 10260
rect 19702 10248 19708 10260
rect 16172 10220 19708 10248
rect 16172 10208 16178 10220
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 20162 10208 20168 10260
rect 20220 10248 20226 10260
rect 20441 10251 20499 10257
rect 20441 10248 20453 10251
rect 20220 10220 20453 10248
rect 20220 10208 20226 10220
rect 20441 10217 20453 10220
rect 20487 10217 20499 10251
rect 20441 10211 20499 10217
rect 20993 10251 21051 10257
rect 20993 10217 21005 10251
rect 21039 10248 21051 10251
rect 22554 10248 22560 10260
rect 21039 10220 22560 10248
rect 21039 10217 21051 10220
rect 20993 10211 21051 10217
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 11974 10140 11980 10192
rect 12032 10180 12038 10192
rect 12437 10183 12495 10189
rect 12437 10180 12449 10183
rect 12032 10152 12449 10180
rect 12032 10140 12038 10152
rect 12437 10149 12449 10152
rect 12483 10149 12495 10183
rect 15654 10180 15660 10192
rect 12437 10143 12495 10149
rect 13096 10152 15660 10180
rect 13096 10121 13124 10152
rect 15654 10140 15660 10152
rect 15712 10140 15718 10192
rect 16574 10140 16580 10192
rect 16632 10180 16638 10192
rect 17586 10180 17592 10192
rect 16632 10152 17592 10180
rect 16632 10140 16638 10152
rect 17586 10140 17592 10152
rect 17644 10140 17650 10192
rect 20622 10180 20628 10192
rect 17696 10152 20628 10180
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 14277 10115 14335 10121
rect 14277 10081 14289 10115
rect 14323 10112 14335 10115
rect 15010 10112 15016 10124
rect 14323 10084 15016 10112
rect 14323 10081 14335 10084
rect 14277 10075 14335 10081
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 16298 10072 16304 10124
rect 16356 10112 16362 10124
rect 16485 10115 16543 10121
rect 16485 10112 16497 10115
rect 16356 10084 16497 10112
rect 16356 10072 16362 10084
rect 16485 10081 16497 10084
rect 16531 10081 16543 10115
rect 17494 10112 17500 10124
rect 17455 10084 17500 10112
rect 16485 10075 16543 10081
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 17696 10121 17724 10152
rect 20622 10140 20628 10152
rect 20680 10140 20686 10192
rect 17681 10115 17739 10121
rect 17681 10081 17693 10115
rect 17727 10081 17739 10115
rect 17681 10075 17739 10081
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18414 10112 18420 10124
rect 18012 10084 18420 10112
rect 18012 10072 18018 10084
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 19521 10115 19579 10121
rect 19521 10081 19533 10115
rect 19567 10112 19579 10115
rect 20438 10112 20444 10124
rect 19567 10084 20444 10112
rect 19567 10081 19579 10084
rect 19521 10075 19579 10081
rect 20438 10072 20444 10084
rect 20496 10072 20502 10124
rect 22002 10072 22008 10124
rect 22060 10112 22066 10124
rect 22370 10112 22376 10124
rect 22060 10084 22376 10112
rect 22060 10072 22066 10084
rect 22370 10072 22376 10084
rect 22428 10072 22434 10124
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 19242 10044 19248 10056
rect 12492 10016 13308 10044
rect 19203 10016 19248 10044
rect 12492 10004 12498 10016
rect 12805 9979 12863 9985
rect 12805 9976 12817 9979
rect 12084 9948 12817 9976
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 12084 9917 12112 9948
rect 12805 9945 12817 9948
rect 12851 9945 12863 9979
rect 13280 9976 13308 10016
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 20809 10047 20867 10053
rect 20809 10044 20821 10047
rect 19352 10016 20821 10044
rect 15562 9976 15568 9988
rect 13280 9948 15568 9976
rect 12805 9939 12863 9945
rect 15562 9936 15568 9948
rect 15620 9936 15626 9988
rect 17405 9979 17463 9985
rect 17405 9945 17417 9979
rect 17451 9976 17463 9979
rect 18049 9979 18107 9985
rect 18049 9976 18061 9979
rect 17451 9948 18061 9976
rect 17451 9945 17463 9948
rect 17405 9939 17463 9945
rect 18049 9945 18061 9948
rect 18095 9945 18107 9979
rect 18049 9939 18107 9945
rect 18322 9936 18328 9988
rect 18380 9976 18386 9988
rect 19352 9976 19380 10016
rect 20809 10013 20821 10016
rect 20855 10013 20867 10047
rect 20809 10007 20867 10013
rect 18380 9948 19380 9976
rect 18380 9936 18386 9948
rect 12069 9911 12127 9917
rect 12069 9908 12081 9911
rect 2832 9880 12081 9908
rect 2832 9868 2838 9880
rect 12069 9877 12081 9880
rect 12115 9877 12127 9911
rect 12069 9871 12127 9877
rect 12897 9911 12955 9917
rect 12897 9877 12909 9911
rect 12943 9908 12955 9911
rect 13354 9908 13360 9920
rect 12943 9880 13360 9908
rect 12943 9877 12955 9880
rect 12897 9871 12955 9877
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 14366 9908 14372 9920
rect 14327 9880 14372 9908
rect 14366 9868 14372 9880
rect 14424 9868 14430 9920
rect 14461 9911 14519 9917
rect 14461 9877 14473 9911
rect 14507 9908 14519 9911
rect 15105 9911 15163 9917
rect 15105 9908 15117 9911
rect 14507 9880 15117 9908
rect 14507 9877 14519 9880
rect 14461 9871 14519 9877
rect 15105 9877 15117 9880
rect 15151 9877 15163 9911
rect 16298 9908 16304 9920
rect 16259 9880 16304 9908
rect 15105 9871 15163 9877
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 16390 9868 16396 9920
rect 16448 9908 16454 9920
rect 17034 9908 17040 9920
rect 16448 9880 16493 9908
rect 16995 9880 17040 9908
rect 16448 9868 16454 9880
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 18506 9908 18512 9920
rect 18467 9880 18512 9908
rect 18506 9868 18512 9880
rect 18564 9908 18570 9920
rect 19981 9911 20039 9917
rect 19981 9908 19993 9911
rect 18564 9880 19993 9908
rect 18564 9868 18570 9880
rect 19981 9877 19993 9880
rect 20027 9877 20039 9911
rect 19981 9871 20039 9877
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 13722 9704 13728 9716
rect 4396 9676 13728 9704
rect 4396 9664 4402 9676
rect 13722 9664 13728 9676
rect 13780 9664 13786 9716
rect 14369 9707 14427 9713
rect 14369 9673 14381 9707
rect 14415 9704 14427 9707
rect 15470 9704 15476 9716
rect 14415 9676 15476 9704
rect 14415 9673 14427 9676
rect 14369 9667 14427 9673
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 12345 9639 12403 9645
rect 12345 9605 12357 9639
rect 12391 9636 12403 9639
rect 13354 9636 13360 9648
rect 12391 9608 13360 9636
rect 12391 9605 12403 9608
rect 12345 9599 12403 9605
rect 13354 9596 13360 9608
rect 13412 9596 13418 9648
rect 15194 9636 15200 9648
rect 14292 9608 15200 9636
rect 12437 9571 12495 9577
rect 12437 9568 12449 9571
rect 11716 9540 12449 9568
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 11716 9373 11744 9540
rect 12437 9537 12449 9540
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 13538 9500 13544 9512
rect 12299 9472 13544 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 14292 9509 14320 9608
rect 15194 9596 15200 9608
rect 15252 9596 15258 9648
rect 16298 9596 16304 9648
rect 16356 9636 16362 9648
rect 16669 9639 16727 9645
rect 16669 9636 16681 9639
rect 16356 9608 16681 9636
rect 16356 9596 16362 9608
rect 16669 9605 16681 9608
rect 16715 9605 16727 9639
rect 16669 9599 16727 9605
rect 18233 9639 18291 9645
rect 18233 9605 18245 9639
rect 18279 9636 18291 9639
rect 18322 9636 18328 9648
rect 18279 9608 18328 9636
rect 18279 9605 18291 9608
rect 18233 9599 18291 9605
rect 18322 9596 18328 9608
rect 18380 9596 18386 9648
rect 20809 9639 20867 9645
rect 20809 9605 20821 9639
rect 20855 9636 20867 9639
rect 20898 9636 20904 9648
rect 20855 9608 20904 9636
rect 20855 9605 20867 9608
rect 20809 9599 20867 9605
rect 20898 9596 20904 9608
rect 20956 9596 20962 9648
rect 21358 9636 21364 9648
rect 21319 9608 21364 9636
rect 21358 9596 21364 9608
rect 21416 9596 21422 9648
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9537 14519 9571
rect 14461 9531 14519 9537
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9469 14335 9503
rect 14277 9463 14335 9469
rect 14476 9500 14504 9531
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 17957 9571 18015 9577
rect 17957 9568 17969 9571
rect 17736 9540 17969 9568
rect 17736 9528 17742 9540
rect 17957 9537 17969 9540
rect 18003 9537 18015 9571
rect 17957 9531 18015 9537
rect 19061 9571 19119 9577
rect 19061 9537 19073 9571
rect 19107 9568 19119 9571
rect 19705 9571 19763 9577
rect 19705 9568 19717 9571
rect 19107 9540 19717 9568
rect 19107 9537 19119 9540
rect 19061 9531 19119 9537
rect 19705 9537 19717 9540
rect 19751 9537 19763 9571
rect 19705 9531 19763 9537
rect 20438 9528 20444 9580
rect 20496 9568 20502 9580
rect 20533 9571 20591 9577
rect 20533 9568 20545 9571
rect 20496 9540 20545 9568
rect 20496 9528 20502 9540
rect 20533 9537 20545 9540
rect 20579 9537 20591 9571
rect 20533 9531 20591 9537
rect 15105 9503 15163 9509
rect 15105 9500 15117 9503
rect 14476 9472 15117 9500
rect 12802 9432 12808 9444
rect 12763 9404 12808 9432
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 14476 9432 14504 9472
rect 15105 9469 15117 9472
rect 15151 9469 15163 9503
rect 15105 9463 15163 9469
rect 15470 9460 15476 9512
rect 15528 9500 15534 9512
rect 15565 9503 15623 9509
rect 15565 9500 15577 9503
rect 15528 9472 15577 9500
rect 15528 9460 15534 9472
rect 15565 9469 15577 9472
rect 15611 9500 15623 9503
rect 18874 9500 18880 9512
rect 15611 9472 18880 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 18874 9460 18880 9472
rect 18932 9460 18938 9512
rect 19797 9503 19855 9509
rect 19797 9469 19809 9503
rect 19843 9469 19855 9503
rect 19797 9463 19855 9469
rect 13780 9404 14504 9432
rect 14829 9435 14887 9441
rect 13780 9392 13786 9404
rect 14829 9401 14841 9435
rect 14875 9432 14887 9435
rect 16390 9432 16396 9444
rect 14875 9404 16396 9432
rect 14875 9401 14887 9404
rect 14829 9395 14887 9401
rect 16390 9392 16396 9404
rect 16448 9392 16454 9444
rect 19242 9392 19248 9444
rect 19300 9432 19306 9444
rect 19337 9435 19395 9441
rect 19337 9432 19349 9435
rect 19300 9404 19349 9432
rect 19300 9392 19306 9404
rect 19337 9401 19349 9404
rect 19383 9401 19395 9435
rect 19337 9395 19395 9401
rect 11701 9367 11759 9373
rect 11701 9364 11713 9367
rect 7156 9336 11713 9364
rect 7156 9324 7162 9336
rect 11701 9333 11713 9336
rect 11747 9333 11759 9367
rect 13354 9364 13360 9376
rect 13315 9336 13360 9364
rect 11701 9327 11759 9333
rect 13354 9324 13360 9336
rect 13412 9364 13418 9376
rect 13633 9367 13691 9373
rect 13633 9364 13645 9367
rect 13412 9336 13645 9364
rect 13412 9324 13418 9336
rect 13633 9333 13645 9336
rect 13679 9333 13691 9367
rect 17494 9364 17500 9376
rect 17455 9336 17500 9364
rect 13633 9327 13691 9333
rect 17494 9324 17500 9336
rect 17552 9364 17558 9376
rect 18138 9364 18144 9376
rect 17552 9336 18144 9364
rect 17552 9324 17558 9336
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 19812 9364 19840 9463
rect 19886 9460 19892 9512
rect 19944 9500 19950 9512
rect 19944 9472 19989 9500
rect 19944 9460 19950 9472
rect 19886 9364 19892 9376
rect 19812 9336 19892 9364
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 11238 9120 11244 9172
rect 11296 9160 11302 9172
rect 17494 9160 17500 9172
rect 11296 9132 17500 9160
rect 11296 9120 11302 9132
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 20070 9092 20076 9104
rect 18064 9064 20076 9092
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 18064 9033 18092 9064
rect 20070 9052 20076 9064
rect 20128 9052 20134 9104
rect 16393 9027 16451 9033
rect 16393 9024 16405 9027
rect 16264 8996 16405 9024
rect 16264 8984 16270 8996
rect 16393 8993 16405 8996
rect 16439 8993 16451 9027
rect 16393 8987 16451 8993
rect 18049 9027 18107 9033
rect 18049 8993 18061 9027
rect 18095 8993 18107 9027
rect 18049 8987 18107 8993
rect 20257 9027 20315 9033
rect 20257 8993 20269 9027
rect 20303 9024 20315 9027
rect 20806 9024 20812 9036
rect 20303 8996 20812 9024
rect 20303 8993 20315 8996
rect 20257 8987 20315 8993
rect 20806 8984 20812 8996
rect 20864 8984 20870 9036
rect 16114 8916 16120 8968
rect 16172 8956 16178 8968
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 16172 8928 16313 8956
rect 16172 8916 16178 8928
rect 16301 8925 16313 8928
rect 16347 8925 16359 8959
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 16301 8919 16359 8925
rect 18616 8928 19257 8956
rect 16209 8891 16267 8897
rect 16209 8857 16221 8891
rect 16255 8888 16267 8891
rect 16853 8891 16911 8897
rect 16853 8888 16865 8891
rect 16255 8860 16865 8888
rect 16255 8857 16267 8860
rect 16209 8851 16267 8857
rect 16853 8857 16865 8860
rect 16899 8857 16911 8891
rect 16853 8851 16911 8857
rect 16942 8848 16948 8900
rect 17000 8888 17006 8900
rect 18233 8891 18291 8897
rect 18233 8888 18245 8891
rect 17000 8860 18245 8888
rect 17000 8848 17006 8860
rect 18233 8857 18245 8860
rect 18279 8857 18291 8891
rect 18233 8851 18291 8857
rect 14550 8820 14556 8832
rect 14511 8792 14556 8820
rect 14550 8780 14556 8792
rect 14608 8780 14614 8832
rect 15194 8780 15200 8832
rect 15252 8820 15258 8832
rect 15841 8823 15899 8829
rect 15841 8820 15853 8823
rect 15252 8792 15853 8820
rect 15252 8780 15258 8792
rect 15841 8789 15853 8792
rect 15887 8789 15899 8823
rect 15841 8783 15899 8789
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 17589 8823 17647 8829
rect 17589 8820 17601 8823
rect 17368 8792 17601 8820
rect 17368 8780 17374 8792
rect 17589 8789 17601 8792
rect 17635 8820 17647 8823
rect 17862 8820 17868 8832
rect 17635 8792 17868 8820
rect 17635 8789 17647 8792
rect 17589 8783 17647 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 18138 8820 18144 8832
rect 18099 8792 18144 8820
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 18616 8829 18644 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 19981 8959 20039 8965
rect 19981 8925 19993 8959
rect 20027 8956 20039 8959
rect 20070 8956 20076 8968
rect 20027 8928 20076 8956
rect 20027 8925 20039 8928
rect 19981 8919 20039 8925
rect 20070 8916 20076 8928
rect 20128 8916 20134 8968
rect 21085 8959 21143 8965
rect 21085 8925 21097 8959
rect 21131 8956 21143 8959
rect 21358 8956 21364 8968
rect 21131 8928 21364 8956
rect 21131 8925 21143 8928
rect 21085 8919 21143 8925
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 19521 8891 19579 8897
rect 19521 8857 19533 8891
rect 19567 8888 19579 8891
rect 20990 8888 20996 8900
rect 19567 8860 20996 8888
rect 19567 8857 19579 8860
rect 19521 8851 19579 8857
rect 20990 8848 20996 8860
rect 21048 8848 21054 8900
rect 18601 8823 18659 8829
rect 18601 8789 18613 8823
rect 18647 8789 18659 8823
rect 20898 8820 20904 8832
rect 20859 8792 20904 8820
rect 18601 8783 18659 8789
rect 20898 8780 20904 8792
rect 20956 8780 20962 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 14550 8616 14556 8628
rect 14511 8588 14556 8616
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 14921 8619 14979 8625
rect 14921 8585 14933 8619
rect 14967 8616 14979 8619
rect 17037 8619 17095 8625
rect 17037 8616 17049 8619
rect 14967 8588 17049 8616
rect 14967 8585 14979 8588
rect 14921 8579 14979 8585
rect 17037 8585 17049 8588
rect 17083 8585 17095 8619
rect 17037 8579 17095 8585
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17678 8616 17684 8628
rect 17184 8588 17229 8616
rect 17639 8588 17684 8616
rect 17184 8576 17190 8588
rect 17678 8576 17684 8588
rect 17736 8576 17742 8628
rect 17770 8576 17776 8628
rect 17828 8616 17834 8628
rect 19337 8619 19395 8625
rect 19337 8616 19349 8619
rect 17828 8588 19349 8616
rect 17828 8576 17834 8588
rect 19337 8585 19349 8588
rect 19383 8585 19395 8619
rect 20438 8616 20444 8628
rect 20399 8588 20444 8616
rect 19337 8579 19395 8585
rect 20438 8576 20444 8588
rect 20496 8576 20502 8628
rect 20993 8619 21051 8625
rect 20993 8585 21005 8619
rect 21039 8616 21051 8619
rect 21634 8616 21640 8628
rect 21039 8588 21640 8616
rect 21039 8585 21051 8588
rect 20993 8579 21051 8585
rect 21634 8576 21640 8588
rect 21692 8576 21698 8628
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 13872 8520 17264 8548
rect 13872 8508 13878 8520
rect 14461 8483 14519 8489
rect 14461 8480 14473 8483
rect 13832 8452 14473 8480
rect 5258 8372 5264 8424
rect 5316 8412 5322 8424
rect 13832 8421 13860 8452
rect 14461 8449 14473 8452
rect 14507 8449 14519 8483
rect 15841 8483 15899 8489
rect 15841 8480 15853 8483
rect 14461 8443 14519 8449
rect 15212 8452 15853 8480
rect 13817 8415 13875 8421
rect 13817 8412 13829 8415
rect 5316 8384 13829 8412
rect 5316 8372 5322 8384
rect 13817 8381 13829 8384
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 14369 8415 14427 8421
rect 14369 8381 14381 8415
rect 14415 8412 14427 8415
rect 14550 8412 14556 8424
rect 14415 8384 14556 8412
rect 14415 8381 14427 8384
rect 14369 8375 14427 8381
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 9122 8304 9128 8356
rect 9180 8344 9186 8356
rect 15212 8353 15240 8452
rect 15841 8449 15853 8452
rect 15887 8449 15899 8483
rect 15841 8443 15899 8449
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8480 15991 8483
rect 16022 8480 16028 8492
rect 15979 8452 16028 8480
rect 15979 8449 15991 8452
rect 15933 8443 15991 8449
rect 16022 8440 16028 8452
rect 16080 8440 16086 8492
rect 17236 8421 17264 8520
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 18049 8483 18107 8489
rect 18049 8480 18061 8483
rect 17368 8452 18061 8480
rect 17368 8440 17374 8452
rect 18049 8449 18061 8452
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 18322 8440 18328 8492
rect 18380 8480 18386 8492
rect 19153 8483 19211 8489
rect 19153 8480 19165 8483
rect 18380 8452 19165 8480
rect 18380 8440 18386 8452
rect 19153 8449 19165 8452
rect 19199 8449 19211 8483
rect 19153 8443 19211 8449
rect 20073 8483 20131 8489
rect 20073 8449 20085 8483
rect 20119 8480 20131 8483
rect 20162 8480 20168 8492
rect 20119 8452 20168 8480
rect 20119 8449 20131 8452
rect 20073 8443 20131 8449
rect 20162 8440 20168 8452
rect 20220 8440 20226 8492
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8480 20867 8483
rect 21082 8480 21088 8492
rect 20855 8452 21088 8480
rect 20855 8449 20867 8452
rect 20809 8443 20867 8449
rect 21082 8440 21088 8452
rect 21140 8440 21146 8492
rect 15749 8415 15807 8421
rect 15749 8381 15761 8415
rect 15795 8381 15807 8415
rect 17221 8415 17279 8421
rect 15749 8375 15807 8381
rect 15948 8384 17172 8412
rect 15197 8347 15255 8353
rect 15197 8344 15209 8347
rect 9180 8316 15209 8344
rect 9180 8304 9186 8316
rect 15197 8313 15209 8316
rect 15243 8313 15255 8347
rect 15764 8344 15792 8375
rect 15948 8344 15976 8384
rect 15764 8316 15976 8344
rect 16301 8347 16359 8353
rect 15197 8307 15255 8313
rect 16301 8313 16313 8347
rect 16347 8344 16359 8347
rect 16942 8344 16948 8356
rect 16347 8316 16948 8344
rect 16347 8313 16359 8316
rect 16301 8307 16359 8313
rect 16942 8304 16948 8316
rect 17000 8304 17006 8356
rect 17144 8344 17172 8384
rect 17221 8381 17233 8415
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 18012 8384 18153 8412
rect 18012 8372 18018 8384
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 18230 8372 18236 8424
rect 18288 8412 18294 8424
rect 19794 8412 19800 8424
rect 18288 8384 18333 8412
rect 19755 8384 19800 8412
rect 18288 8372 18294 8384
rect 19794 8372 19800 8384
rect 19852 8372 19858 8424
rect 19978 8412 19984 8424
rect 19939 8384 19984 8412
rect 19978 8372 19984 8384
rect 20036 8372 20042 8424
rect 18598 8344 18604 8356
rect 17144 8316 18604 8344
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 18874 8304 18880 8356
rect 18932 8344 18938 8356
rect 18932 8316 19288 8344
rect 18932 8304 18938 8316
rect 16669 8279 16727 8285
rect 16669 8245 16681 8279
rect 16715 8276 16727 8279
rect 16758 8276 16764 8288
rect 16715 8248 16764 8276
rect 16715 8245 16727 8248
rect 16669 8239 16727 8245
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 18690 8276 18696 8288
rect 18651 8248 18696 8276
rect 18690 8236 18696 8248
rect 18748 8236 18754 8288
rect 19260 8276 19288 8316
rect 20990 8276 20996 8288
rect 19260 8248 20996 8276
rect 20990 8236 20996 8248
rect 21048 8236 21054 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 14366 8032 14372 8084
rect 14424 8072 14430 8084
rect 14829 8075 14887 8081
rect 14829 8072 14841 8075
rect 14424 8044 14841 8072
rect 14424 8032 14430 8044
rect 14829 8041 14841 8044
rect 14875 8041 14887 8075
rect 14829 8035 14887 8041
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18417 8075 18475 8081
rect 18417 8072 18429 8075
rect 18196 8044 18429 8072
rect 18196 8032 18202 8044
rect 18417 8041 18429 8044
rect 18463 8041 18475 8075
rect 18417 8035 18475 8041
rect 19978 8032 19984 8084
rect 20036 8072 20042 8084
rect 20349 8075 20407 8081
rect 20349 8072 20361 8075
rect 20036 8044 20361 8072
rect 20036 8032 20042 8044
rect 20349 8041 20361 8044
rect 20395 8041 20407 8075
rect 20349 8035 20407 8041
rect 13262 7896 13268 7948
rect 13320 7936 13326 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 13320 7908 14197 7936
rect 13320 7896 13326 7908
rect 14185 7905 14197 7908
rect 14231 7905 14243 7939
rect 14185 7899 14243 7905
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7936 15899 7939
rect 16022 7936 16028 7948
rect 15887 7908 16028 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 17865 7939 17923 7945
rect 17865 7905 17877 7939
rect 17911 7936 17923 7939
rect 18598 7936 18604 7948
rect 17911 7908 18604 7936
rect 17911 7905 17923 7908
rect 17865 7899 17923 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 19518 7936 19524 7948
rect 19479 7908 19524 7936
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 20993 7939 21051 7945
rect 20993 7905 21005 7939
rect 21039 7936 21051 7939
rect 21174 7936 21180 7948
rect 21039 7908 21180 7936
rect 21039 7905 21051 7908
rect 20993 7899 21051 7905
rect 21174 7896 21180 7908
rect 21232 7896 21238 7948
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5776 7840 5825 7868
rect 5776 7828 5782 7840
rect 5813 7837 5825 7840
rect 5859 7868 5871 7871
rect 6089 7871 6147 7877
rect 6089 7868 6101 7871
rect 5859 7840 6101 7868
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 6089 7837 6101 7840
rect 6135 7837 6147 7871
rect 16758 7868 16764 7880
rect 16719 7840 16764 7868
rect 6089 7831 6147 7837
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7868 17095 7871
rect 18322 7868 18328 7880
rect 17083 7840 18328 7868
rect 17083 7837 17095 7840
rect 17037 7831 17095 7837
rect 18322 7828 18328 7840
rect 18380 7828 18386 7880
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 19116 7840 19257 7868
rect 19116 7828 19122 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 14461 7803 14519 7809
rect 14461 7800 14473 7803
rect 13648 7772 14473 7800
rect 5626 7732 5632 7744
rect 5587 7704 5632 7732
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 13648 7741 13676 7772
rect 14461 7769 14473 7772
rect 14507 7769 14519 7803
rect 14461 7763 14519 7769
rect 16485 7803 16543 7809
rect 16485 7769 16497 7803
rect 16531 7800 16543 7803
rect 17957 7803 18015 7809
rect 17957 7800 17969 7803
rect 16531 7772 17969 7800
rect 16531 7769 16543 7772
rect 16485 7763 16543 7769
rect 17957 7769 17969 7772
rect 18003 7800 18015 7803
rect 18230 7800 18236 7812
rect 18003 7772 18236 7800
rect 18003 7769 18015 7772
rect 17957 7763 18015 7769
rect 18230 7760 18236 7772
rect 18288 7800 18294 7812
rect 18782 7800 18788 7812
rect 18288 7772 18788 7800
rect 18288 7760 18294 7772
rect 18782 7760 18788 7772
rect 18840 7800 18846 7812
rect 19981 7803 20039 7809
rect 19981 7800 19993 7803
rect 18840 7772 19993 7800
rect 18840 7760 18846 7772
rect 19981 7769 19993 7772
rect 20027 7800 20039 7803
rect 21082 7800 21088 7812
rect 20027 7772 21088 7800
rect 20027 7769 20039 7772
rect 19981 7763 20039 7769
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 13633 7735 13691 7741
rect 13633 7732 13645 7735
rect 13596 7704 13645 7732
rect 13596 7692 13602 7704
rect 13633 7701 13645 7704
rect 13679 7701 13691 7735
rect 13633 7695 13691 7701
rect 14369 7735 14427 7741
rect 14369 7701 14381 7735
rect 14415 7732 14427 7735
rect 15197 7735 15255 7741
rect 15197 7732 15209 7735
rect 14415 7704 15209 7732
rect 14415 7701 14427 7704
rect 14369 7695 14427 7701
rect 15197 7701 15209 7704
rect 15243 7732 15255 7735
rect 15286 7732 15292 7744
rect 15243 7704 15292 7732
rect 15243 7701 15255 7704
rect 15197 7695 15255 7701
rect 15286 7692 15292 7704
rect 15344 7692 15350 7744
rect 15562 7732 15568 7744
rect 15523 7704 15568 7732
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 18049 7735 18107 7741
rect 18049 7701 18061 7735
rect 18095 7732 18107 7735
rect 18138 7732 18144 7744
rect 18095 7704 18144 7732
rect 18095 7701 18107 7704
rect 18049 7695 18107 7701
rect 18138 7692 18144 7704
rect 18196 7732 18202 7744
rect 18690 7732 18696 7744
rect 18196 7704 18696 7732
rect 18196 7692 18202 7704
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 20714 7732 20720 7744
rect 20675 7704 20720 7732
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 20864 7704 20909 7732
rect 20864 7692 20870 7704
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 13446 7528 13452 7540
rect 5684 7500 13452 7528
rect 5684 7488 5690 7500
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 13630 7528 13636 7540
rect 13591 7500 13636 7528
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 14093 7531 14151 7537
rect 14093 7497 14105 7531
rect 14139 7528 14151 7531
rect 14737 7531 14795 7537
rect 14737 7528 14749 7531
rect 14139 7500 14749 7528
rect 14139 7497 14151 7500
rect 14093 7491 14151 7497
rect 14737 7497 14749 7500
rect 14783 7528 14795 7531
rect 15286 7528 15292 7540
rect 14783 7500 15292 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 15286 7488 15292 7500
rect 15344 7528 15350 7540
rect 16022 7528 16028 7540
rect 15344 7500 16028 7528
rect 15344 7488 15350 7500
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 17126 7488 17132 7540
rect 17184 7528 17190 7540
rect 17313 7531 17371 7537
rect 17313 7528 17325 7531
rect 17184 7500 17325 7528
rect 17184 7488 17190 7500
rect 17313 7497 17325 7500
rect 17359 7497 17371 7531
rect 17313 7491 17371 7497
rect 17773 7531 17831 7537
rect 17773 7497 17785 7531
rect 17819 7528 17831 7531
rect 18230 7528 18236 7540
rect 17819 7500 18236 7528
rect 17819 7497 17831 7500
rect 17773 7491 17831 7497
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 19058 7528 19064 7540
rect 19019 7500 19064 7528
rect 19058 7488 19064 7500
rect 19116 7488 19122 7540
rect 20070 7528 20076 7540
rect 20031 7500 20076 7528
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 20625 7531 20683 7537
rect 20625 7497 20637 7531
rect 20671 7528 20683 7531
rect 20806 7528 20812 7540
rect 20671 7500 20812 7528
rect 20671 7497 20683 7500
rect 20625 7491 20683 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 21082 7528 21088 7540
rect 21043 7500 21088 7528
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 14608 7432 16804 7460
rect 14608 7420 14614 7432
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 12406 7364 13369 7392
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 12406 7188 12434 7364
rect 13357 7361 13369 7364
rect 13403 7392 13415 7395
rect 14001 7395 14059 7401
rect 14001 7392 14013 7395
rect 13403 7364 14013 7392
rect 13403 7361 13415 7364
rect 13357 7355 13415 7361
rect 14001 7361 14013 7364
rect 14047 7361 14059 7395
rect 15654 7392 15660 7404
rect 15615 7364 15660 7392
rect 14001 7355 14059 7361
rect 15654 7352 15660 7364
rect 15712 7352 15718 7404
rect 14274 7324 14280 7336
rect 14235 7296 14280 7324
rect 14274 7284 14280 7296
rect 14332 7284 14338 7336
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7293 15439 7327
rect 15562 7324 15568 7336
rect 15523 7296 15568 7324
rect 15381 7287 15439 7293
rect 11020 7160 12434 7188
rect 15396 7188 15424 7287
rect 15562 7284 15568 7296
rect 15620 7284 15626 7336
rect 16666 7324 16672 7336
rect 16627 7296 16672 7324
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 16776 7324 16804 7432
rect 16942 7420 16948 7472
rect 17000 7460 17006 7472
rect 18693 7463 18751 7469
rect 18693 7460 18705 7463
rect 17000 7432 18705 7460
rect 17000 7420 17006 7432
rect 18693 7429 18705 7432
rect 18739 7429 18751 7463
rect 20530 7460 20536 7472
rect 18693 7423 18751 7429
rect 18800 7432 20536 7460
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 18138 7392 18144 7404
rect 17727 7364 18144 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 18800 7392 18828 7432
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 18432 7364 18828 7392
rect 18432 7333 18460 7364
rect 18874 7352 18880 7404
rect 18932 7392 18938 7404
rect 19705 7395 19763 7401
rect 19705 7392 19717 7395
rect 18932 7364 19717 7392
rect 18932 7352 18938 7364
rect 19705 7361 19717 7364
rect 19751 7361 19763 7395
rect 20990 7392 20996 7404
rect 20951 7364 20996 7392
rect 19705 7355 19763 7361
rect 20990 7352 20996 7364
rect 21048 7352 21054 7404
rect 17865 7327 17923 7333
rect 17865 7324 17877 7327
rect 16776 7296 17877 7324
rect 17865 7293 17877 7296
rect 17911 7293 17923 7327
rect 17865 7287 17923 7293
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7293 18475 7327
rect 18598 7324 18604 7336
rect 18559 7296 18604 7324
rect 18417 7287 18475 7293
rect 18598 7284 18604 7296
rect 18656 7284 18662 7336
rect 19518 7324 19524 7336
rect 19479 7296 19524 7324
rect 19518 7284 19524 7296
rect 19576 7284 19582 7336
rect 19613 7327 19671 7333
rect 19613 7293 19625 7327
rect 19659 7293 19671 7327
rect 19613 7287 19671 7293
rect 21269 7327 21327 7333
rect 21269 7293 21281 7327
rect 21315 7324 21327 7327
rect 21542 7324 21548 7336
rect 21315 7296 21548 7324
rect 21315 7293 21327 7296
rect 21269 7287 21327 7293
rect 16025 7259 16083 7265
rect 16025 7225 16037 7259
rect 16071 7256 16083 7259
rect 17310 7256 17316 7268
rect 16071 7228 17316 7256
rect 16071 7225 16083 7228
rect 16025 7219 16083 7225
rect 17310 7216 17316 7228
rect 17368 7216 17374 7268
rect 19628 7256 19656 7287
rect 21542 7284 21548 7296
rect 21600 7284 21606 7336
rect 19702 7256 19708 7268
rect 19628 7228 19708 7256
rect 19702 7216 19708 7228
rect 19760 7216 19766 7268
rect 17402 7188 17408 7200
rect 15396 7160 17408 7188
rect 11020 7148 11026 7160
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 20070 6984 20076 6996
rect 13504 6956 20076 6984
rect 13504 6944 13510 6956
rect 20070 6944 20076 6956
rect 20128 6944 20134 6996
rect 20625 6987 20683 6993
rect 20625 6953 20637 6987
rect 20671 6984 20683 6987
rect 20714 6984 20720 6996
rect 20671 6956 20720 6984
rect 20671 6953 20683 6956
rect 20625 6947 20683 6953
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 17497 6919 17555 6925
rect 17497 6885 17509 6919
rect 17543 6885 17555 6919
rect 17497 6879 17555 6885
rect 15013 6851 15071 6857
rect 15013 6817 15025 6851
rect 15059 6848 15071 6851
rect 15286 6848 15292 6860
rect 15059 6820 15292 6848
rect 15059 6817 15071 6820
rect 15013 6811 15071 6817
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 15473 6851 15531 6857
rect 15473 6817 15485 6851
rect 15519 6848 15531 6851
rect 15654 6848 15660 6860
rect 15519 6820 15660 6848
rect 15519 6817 15531 6820
rect 15473 6811 15531 6817
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 15764 6820 16313 6848
rect 15304 6780 15332 6808
rect 15764 6780 15792 6820
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16301 6811 16359 6817
rect 16390 6808 16396 6860
rect 16448 6848 16454 6860
rect 16945 6851 17003 6857
rect 16448 6820 16896 6848
rect 16448 6808 16454 6820
rect 15304 6752 15792 6780
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6780 16175 6783
rect 16666 6780 16672 6792
rect 16163 6752 16672 6780
rect 16163 6749 16175 6752
rect 16117 6743 16175 6749
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 16868 6780 16896 6820
rect 16945 6817 16957 6851
rect 16991 6848 17003 6851
rect 17402 6848 17408 6860
rect 16991 6820 17408 6848
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 17512 6848 17540 6879
rect 17862 6876 17868 6928
rect 17920 6916 17926 6928
rect 17920 6888 18460 6916
rect 17920 6876 17926 6888
rect 17954 6848 17960 6860
rect 17512 6820 17960 6848
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 18046 6808 18052 6860
rect 18104 6848 18110 6860
rect 18325 6851 18383 6857
rect 18325 6848 18337 6851
rect 18104 6820 18337 6848
rect 18104 6808 18110 6820
rect 18325 6817 18337 6820
rect 18371 6817 18383 6851
rect 18325 6811 18383 6817
rect 18230 6780 18236 6792
rect 16868 6752 18092 6780
rect 18191 6752 18236 6780
rect 16209 6715 16267 6721
rect 16209 6681 16221 6715
rect 16255 6712 16267 6715
rect 18064 6712 18092 6752
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 18432 6780 18460 6888
rect 18782 6876 18788 6928
rect 18840 6916 18846 6928
rect 20257 6919 20315 6925
rect 20257 6916 20269 6919
rect 18840 6888 20269 6916
rect 18840 6876 18846 6888
rect 20257 6885 20269 6888
rect 20303 6885 20315 6919
rect 21174 6916 21180 6928
rect 20257 6879 20315 6885
rect 20640 6888 21180 6916
rect 19429 6851 19487 6857
rect 19429 6817 19441 6851
rect 19475 6848 19487 6851
rect 20640 6848 20668 6888
rect 21174 6876 21180 6888
rect 21232 6876 21238 6928
rect 19475 6820 20668 6848
rect 19475 6817 19487 6820
rect 19429 6811 19487 6817
rect 20714 6808 20720 6860
rect 20772 6848 20778 6860
rect 21269 6851 21327 6857
rect 21269 6848 21281 6851
rect 20772 6820 21281 6848
rect 20772 6808 20778 6820
rect 21269 6817 21281 6820
rect 21315 6848 21327 6851
rect 21542 6848 21548 6860
rect 21315 6820 21548 6848
rect 21315 6817 21327 6820
rect 21269 6811 21327 6817
rect 21542 6808 21548 6820
rect 21600 6808 21606 6860
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 18432 6752 21005 6780
rect 20993 6749 21005 6752
rect 21039 6780 21051 6783
rect 21634 6780 21640 6792
rect 21039 6752 21640 6780
rect 21039 6749 21051 6752
rect 20993 6743 21051 6749
rect 21634 6740 21640 6752
rect 21692 6740 21698 6792
rect 18141 6715 18199 6721
rect 18141 6712 18153 6715
rect 16255 6684 17816 6712
rect 18064 6684 18153 6712
rect 16255 6681 16267 6684
rect 16209 6675 16267 6681
rect 13354 6604 13360 6656
rect 13412 6644 13418 6656
rect 14645 6647 14703 6653
rect 14645 6644 14657 6647
rect 13412 6616 14657 6644
rect 13412 6604 13418 6616
rect 14645 6613 14657 6616
rect 14691 6644 14703 6647
rect 15654 6644 15660 6656
rect 14691 6616 15660 6644
rect 14691 6613 14703 6616
rect 14645 6607 14703 6613
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 15749 6647 15807 6653
rect 15749 6613 15761 6647
rect 15795 6644 15807 6647
rect 16114 6644 16120 6656
rect 15795 6616 16120 6644
rect 15795 6613 15807 6616
rect 15749 6607 15807 6613
rect 16114 6604 16120 6616
rect 16172 6604 16178 6656
rect 16298 6604 16304 6656
rect 16356 6644 16362 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 16356 6616 17049 6644
rect 16356 6604 16362 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 17037 6607 17095 6613
rect 17129 6647 17187 6653
rect 17129 6613 17141 6647
rect 17175 6644 17187 6647
rect 17402 6644 17408 6656
rect 17175 6616 17408 6644
rect 17175 6613 17187 6616
rect 17129 6607 17187 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 17788 6653 17816 6684
rect 18141 6681 18153 6684
rect 18187 6712 18199 6715
rect 18506 6712 18512 6724
rect 18187 6684 18512 6712
rect 18187 6681 18199 6684
rect 18141 6675 18199 6681
rect 18506 6672 18512 6684
rect 18564 6712 18570 6724
rect 18785 6715 18843 6721
rect 18785 6712 18797 6715
rect 18564 6684 18797 6712
rect 18564 6672 18570 6684
rect 18785 6681 18797 6684
rect 18831 6681 18843 6715
rect 22186 6712 22192 6724
rect 18785 6675 18843 6681
rect 18892 6684 22192 6712
rect 17773 6647 17831 6653
rect 17773 6613 17785 6647
rect 17819 6613 17831 6647
rect 17773 6607 17831 6613
rect 17862 6604 17868 6656
rect 17920 6644 17926 6656
rect 18892 6644 18920 6684
rect 22186 6672 22192 6684
rect 22244 6672 22250 6724
rect 19518 6644 19524 6656
rect 17920 6616 18920 6644
rect 19479 6616 19524 6644
rect 17920 6604 17926 6616
rect 19518 6604 19524 6616
rect 19576 6604 19582 6656
rect 19610 6604 19616 6656
rect 19668 6644 19674 6656
rect 19981 6647 20039 6653
rect 19668 6616 19713 6644
rect 19668 6604 19674 6616
rect 19981 6613 19993 6647
rect 20027 6644 20039 6647
rect 20162 6644 20168 6656
rect 20027 6616 20168 6644
rect 20027 6613 20039 6616
rect 19981 6607 20039 6613
rect 20162 6604 20168 6616
rect 20220 6604 20226 6656
rect 21085 6647 21143 6653
rect 21085 6613 21097 6647
rect 21131 6644 21143 6647
rect 21542 6644 21548 6656
rect 21131 6616 21548 6644
rect 21131 6613 21143 6616
rect 21085 6607 21143 6613
rect 21542 6604 21548 6616
rect 21600 6604 21606 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 15841 6443 15899 6449
rect 15841 6409 15853 6443
rect 15887 6440 15899 6443
rect 15930 6440 15936 6452
rect 15887 6412 15936 6440
rect 15887 6409 15899 6412
rect 15841 6403 15899 6409
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 16298 6440 16304 6452
rect 16259 6412 16304 6440
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 17402 6440 17408 6452
rect 17363 6412 17408 6440
rect 17402 6400 17408 6412
rect 17460 6400 17466 6452
rect 18417 6443 18475 6449
rect 18417 6409 18429 6443
rect 18463 6440 18475 6443
rect 18598 6440 18604 6452
rect 18463 6412 18604 6440
rect 18463 6409 18475 6412
rect 18417 6403 18475 6409
rect 18598 6400 18604 6412
rect 18656 6400 18662 6452
rect 19245 6443 19303 6449
rect 19245 6409 19257 6443
rect 19291 6440 19303 6443
rect 19610 6440 19616 6452
rect 19291 6412 19616 6440
rect 19291 6409 19303 6412
rect 19245 6403 19303 6409
rect 19610 6400 19616 6412
rect 19668 6400 19674 6452
rect 19981 6443 20039 6449
rect 19981 6409 19993 6443
rect 20027 6440 20039 6443
rect 20533 6443 20591 6449
rect 20533 6440 20545 6443
rect 20027 6412 20545 6440
rect 20027 6409 20039 6412
rect 19981 6403 20039 6409
rect 20533 6409 20545 6412
rect 20579 6409 20591 6443
rect 20533 6403 20591 6409
rect 20993 6443 21051 6449
rect 20993 6409 21005 6443
rect 21039 6440 21051 6443
rect 21082 6440 21088 6452
rect 21039 6412 21088 6440
rect 21039 6409 21051 6412
rect 20993 6403 21051 6409
rect 21082 6400 21088 6412
rect 21140 6400 21146 6452
rect 16390 6372 16396 6384
rect 12406 6344 16396 6372
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 12406 6100 12434 6344
rect 16390 6332 16396 6344
rect 16448 6332 16454 6384
rect 19426 6372 19432 6384
rect 16960 6344 19432 6372
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6304 14795 6307
rect 15194 6304 15200 6316
rect 14783 6276 15200 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16022 6304 16028 6316
rect 15979 6276 16028 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16022 6264 16028 6276
rect 16080 6264 16086 6316
rect 16960 6304 16988 6344
rect 19426 6332 19432 6344
rect 19484 6332 19490 6384
rect 16868 6276 16988 6304
rect 17037 6307 17095 6313
rect 12894 6196 12900 6248
rect 12952 6236 12958 6248
rect 14461 6239 14519 6245
rect 14461 6236 14473 6239
rect 12952 6208 14473 6236
rect 12952 6196 12958 6208
rect 14461 6205 14473 6208
rect 14507 6205 14519 6239
rect 14461 6199 14519 6205
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6236 15807 6239
rect 16298 6236 16304 6248
rect 15795 6208 16304 6236
rect 15795 6205 15807 6208
rect 15749 6199 15807 6205
rect 16298 6196 16304 6208
rect 16356 6236 16362 6248
rect 16868 6245 16896 6276
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17862 6304 17868 6316
rect 17083 6276 17724 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 16853 6239 16911 6245
rect 16853 6236 16865 6239
rect 16356 6208 16865 6236
rect 16356 6196 16362 6208
rect 16853 6205 16865 6208
rect 16899 6205 16911 6239
rect 16853 6199 16911 6205
rect 16945 6239 17003 6245
rect 16945 6205 16957 6239
rect 16991 6236 17003 6239
rect 17402 6236 17408 6248
rect 16991 6208 17408 6236
rect 16991 6205 17003 6208
rect 16945 6199 17003 6205
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 9824 6072 12434 6100
rect 15289 6103 15347 6109
rect 9824 6060 9830 6072
rect 15289 6069 15301 6103
rect 15335 6100 15347 6103
rect 15930 6100 15936 6112
rect 15335 6072 15936 6100
rect 15335 6069 15347 6072
rect 15289 6063 15347 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 17696 6100 17724 6276
rect 17788 6276 17868 6304
rect 17788 6245 17816 6276
rect 17862 6264 17868 6276
rect 17920 6264 17926 6316
rect 18046 6304 18052 6316
rect 18007 6276 18052 6304
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6304 19947 6307
rect 20530 6304 20536 6316
rect 19935 6276 20536 6304
rect 19935 6273 19947 6276
rect 19889 6267 19947 6273
rect 20530 6264 20536 6276
rect 20588 6264 20594 6316
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6304 20959 6307
rect 20990 6304 20996 6316
rect 20947 6276 20996 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 20990 6264 20996 6276
rect 21048 6304 21054 6316
rect 21358 6304 21364 6316
rect 21048 6276 21364 6304
rect 21048 6264 21054 6276
rect 21358 6264 21364 6276
rect 21416 6264 21422 6316
rect 17773 6239 17831 6245
rect 17773 6205 17785 6239
rect 17819 6205 17831 6239
rect 17954 6236 17960 6248
rect 17915 6208 17960 6236
rect 17773 6199 17831 6205
rect 17954 6196 17960 6208
rect 18012 6196 18018 6248
rect 18966 6196 18972 6248
rect 19024 6236 19030 6248
rect 20073 6239 20131 6245
rect 20073 6236 20085 6239
rect 19024 6208 20085 6236
rect 19024 6196 19030 6208
rect 20073 6205 20085 6208
rect 20119 6205 20131 6239
rect 20073 6199 20131 6205
rect 21174 6196 21180 6248
rect 21232 6236 21238 6248
rect 22462 6236 22468 6248
rect 21232 6208 22468 6236
rect 21232 6196 21238 6208
rect 22462 6196 22468 6208
rect 22520 6196 22526 6248
rect 19521 6171 19579 6177
rect 19521 6137 19533 6171
rect 19567 6168 19579 6171
rect 19702 6168 19708 6180
rect 19567 6140 19708 6168
rect 19567 6137 19579 6140
rect 19521 6131 19579 6137
rect 19702 6128 19708 6140
rect 19760 6128 19766 6180
rect 18322 6100 18328 6112
rect 17696 6072 18328 6100
rect 18322 6060 18328 6072
rect 18380 6060 18386 6112
rect 18782 6100 18788 6112
rect 18743 6072 18788 6100
rect 18782 6060 18788 6072
rect 18840 6060 18846 6112
rect 19426 6060 19432 6112
rect 19484 6100 19490 6112
rect 19610 6100 19616 6112
rect 19484 6072 19616 6100
rect 19484 6060 19490 6072
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 20070 6060 20076 6112
rect 20128 6100 20134 6112
rect 20806 6100 20812 6112
rect 20128 6072 20812 6100
rect 20128 6060 20134 6072
rect 20806 6060 20812 6072
rect 20864 6060 20870 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 16209 5899 16267 5905
rect 16209 5865 16221 5899
rect 16255 5896 16267 5899
rect 16942 5896 16948 5908
rect 16255 5868 16948 5896
rect 16255 5865 16267 5868
rect 16209 5859 16267 5865
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 17862 5896 17868 5908
rect 17052 5868 17868 5896
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 17052 5760 17080 5868
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 18874 5896 18880 5908
rect 18835 5868 18880 5896
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 19518 5896 19524 5908
rect 19479 5868 19524 5896
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 20530 5896 20536 5908
rect 20491 5868 20536 5896
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 17773 5831 17831 5837
rect 17773 5797 17785 5831
rect 17819 5828 17831 5831
rect 19886 5828 19892 5840
rect 17819 5800 19892 5828
rect 17819 5797 17831 5800
rect 17773 5791 17831 5797
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 17218 5760 17224 5772
rect 15703 5732 17080 5760
rect 17179 5732 17224 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 17218 5720 17224 5732
rect 17276 5720 17282 5772
rect 18325 5763 18383 5769
rect 18325 5729 18337 5763
rect 18371 5760 18383 5763
rect 18966 5760 18972 5772
rect 18371 5732 18972 5760
rect 18371 5729 18383 5732
rect 18325 5723 18383 5729
rect 18966 5720 18972 5732
rect 19024 5720 19030 5772
rect 20165 5763 20223 5769
rect 20165 5729 20177 5763
rect 20211 5760 20223 5763
rect 20714 5760 20720 5772
rect 20211 5732 20720 5760
rect 20211 5729 20223 5732
rect 20165 5723 20223 5729
rect 20714 5720 20720 5732
rect 20772 5720 20778 5772
rect 21174 5760 21180 5772
rect 21135 5732 21180 5760
rect 21174 5720 21180 5732
rect 21232 5720 21238 5772
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5692 14611 5695
rect 14734 5692 14740 5704
rect 14599 5664 14740 5692
rect 14599 5661 14611 5664
rect 14553 5655 14611 5661
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 16022 5652 16028 5704
rect 16080 5692 16086 5704
rect 18874 5692 18880 5704
rect 16080 5664 18880 5692
rect 16080 5652 16086 5664
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 13446 5584 13452 5636
rect 13504 5624 13510 5636
rect 14277 5627 14335 5633
rect 14277 5624 14289 5627
rect 13504 5596 14289 5624
rect 13504 5584 13510 5596
rect 14277 5593 14289 5596
rect 14323 5593 14335 5627
rect 14277 5587 14335 5593
rect 15841 5627 15899 5633
rect 15841 5593 15853 5627
rect 15887 5624 15899 5627
rect 16485 5627 16543 5633
rect 16485 5624 16497 5627
rect 15887 5596 16497 5624
rect 15887 5593 15899 5596
rect 15841 5587 15899 5593
rect 16485 5593 16497 5596
rect 16531 5593 16543 5627
rect 16485 5587 16543 5593
rect 17126 5584 17132 5636
rect 17184 5624 17190 5636
rect 17405 5627 17463 5633
rect 17405 5624 17417 5627
rect 17184 5596 17417 5624
rect 17184 5584 17190 5596
rect 17405 5593 17417 5596
rect 17451 5593 17463 5627
rect 17405 5587 17463 5593
rect 18690 5584 18696 5636
rect 18748 5624 18754 5636
rect 20901 5627 20959 5633
rect 18748 5596 20024 5624
rect 18748 5584 18754 5596
rect 15194 5556 15200 5568
rect 15155 5528 15200 5556
rect 15194 5516 15200 5528
rect 15252 5556 15258 5568
rect 15749 5559 15807 5565
rect 15749 5556 15761 5559
rect 15252 5528 15761 5556
rect 15252 5516 15258 5528
rect 15749 5525 15761 5528
rect 15795 5525 15807 5559
rect 15749 5519 15807 5525
rect 15930 5516 15936 5568
rect 15988 5556 15994 5568
rect 17313 5559 17371 5565
rect 17313 5556 17325 5559
rect 15988 5528 17325 5556
rect 15988 5516 15994 5528
rect 17313 5525 17325 5528
rect 17359 5556 17371 5559
rect 17770 5556 17776 5568
rect 17359 5528 17776 5556
rect 17359 5525 17371 5528
rect 17313 5519 17371 5525
rect 17770 5516 17776 5528
rect 17828 5516 17834 5568
rect 18414 5556 18420 5568
rect 18375 5528 18420 5556
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 18506 5516 18512 5568
rect 18564 5556 18570 5568
rect 18564 5528 18609 5556
rect 18564 5516 18570 5528
rect 19610 5516 19616 5568
rect 19668 5556 19674 5568
rect 19996 5565 20024 5596
rect 20901 5593 20913 5627
rect 20947 5624 20959 5627
rect 21634 5624 21640 5636
rect 20947 5596 21640 5624
rect 20947 5593 20959 5596
rect 20901 5587 20959 5593
rect 21634 5584 21640 5596
rect 21692 5584 21698 5636
rect 19889 5559 19947 5565
rect 19889 5556 19901 5559
rect 19668 5528 19901 5556
rect 19668 5516 19674 5528
rect 19889 5525 19901 5528
rect 19935 5525 19947 5559
rect 19889 5519 19947 5525
rect 19981 5559 20039 5565
rect 19981 5525 19993 5559
rect 20027 5556 20039 5559
rect 20714 5556 20720 5568
rect 20027 5528 20720 5556
rect 20027 5525 20039 5528
rect 19981 5519 20039 5525
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 20990 5516 20996 5568
rect 21048 5556 21054 5568
rect 21542 5556 21548 5568
rect 21048 5528 21548 5556
rect 21048 5516 21054 5528
rect 21542 5516 21548 5528
rect 21600 5516 21606 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 15565 5355 15623 5361
rect 15565 5321 15577 5355
rect 15611 5352 15623 5355
rect 15654 5352 15660 5364
rect 15611 5324 15660 5352
rect 15611 5321 15623 5324
rect 15565 5315 15623 5321
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 16298 5352 16304 5364
rect 16259 5324 16304 5352
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 17678 5312 17684 5364
rect 17736 5312 17742 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18233 5355 18291 5361
rect 18233 5352 18245 5355
rect 18012 5324 18245 5352
rect 18012 5312 18018 5324
rect 18233 5321 18245 5324
rect 18279 5321 18291 5355
rect 18233 5315 18291 5321
rect 18506 5312 18512 5364
rect 18564 5352 18570 5364
rect 18693 5355 18751 5361
rect 18693 5352 18705 5355
rect 18564 5324 18705 5352
rect 18564 5312 18570 5324
rect 18693 5321 18705 5324
rect 18739 5321 18751 5355
rect 18693 5315 18751 5321
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19521 5355 19579 5361
rect 19521 5352 19533 5355
rect 19484 5324 19533 5352
rect 19484 5312 19490 5324
rect 19521 5321 19533 5324
rect 19567 5321 19579 5355
rect 20990 5352 20996 5364
rect 20951 5324 20996 5352
rect 19521 5315 19579 5321
rect 20990 5312 20996 5324
rect 21048 5312 21054 5364
rect 15197 5287 15255 5293
rect 15197 5253 15209 5287
rect 15243 5284 15255 5287
rect 17696 5284 17724 5312
rect 15243 5256 17724 5284
rect 17865 5287 17923 5293
rect 15243 5253 15255 5256
rect 15197 5247 15255 5253
rect 17865 5253 17877 5287
rect 17911 5284 17923 5287
rect 18874 5284 18880 5296
rect 17911 5256 18880 5284
rect 17911 5253 17923 5256
rect 17865 5247 17923 5253
rect 18874 5244 18880 5256
rect 18932 5284 18938 5296
rect 20257 5287 20315 5293
rect 20257 5284 20269 5287
rect 18932 5256 20269 5284
rect 18932 5244 18938 5256
rect 20257 5253 20269 5256
rect 20303 5253 20315 5287
rect 20257 5247 20315 5253
rect 17034 5176 17040 5228
rect 17092 5216 17098 5228
rect 17129 5219 17187 5225
rect 17129 5216 17141 5219
rect 17092 5188 17141 5216
rect 17092 5176 17098 5188
rect 17129 5185 17141 5188
rect 17175 5185 17187 5219
rect 17129 5179 17187 5185
rect 20809 5219 20867 5225
rect 20809 5185 20821 5219
rect 20855 5216 20867 5219
rect 21266 5216 21272 5228
rect 20855 5188 21272 5216
rect 20855 5185 20867 5188
rect 20809 5179 20867 5185
rect 21266 5176 21272 5188
rect 21324 5176 21330 5228
rect 16022 5108 16028 5160
rect 16080 5148 16086 5160
rect 16853 5151 16911 5157
rect 16853 5148 16865 5151
rect 16080 5120 16865 5148
rect 16080 5108 16086 5120
rect 16853 5117 16865 5120
rect 16899 5117 16911 5151
rect 17678 5148 17684 5160
rect 17639 5120 17684 5148
rect 16853 5111 16911 5117
rect 17678 5108 17684 5120
rect 17736 5108 17742 5160
rect 17770 5108 17776 5160
rect 17828 5148 17834 5160
rect 17828 5120 19748 5148
rect 17828 5108 17834 5120
rect 15933 5083 15991 5089
rect 15933 5049 15945 5083
rect 15979 5080 15991 5083
rect 18690 5080 18696 5092
rect 15979 5052 18696 5080
rect 15979 5049 15991 5052
rect 15933 5043 15991 5049
rect 18690 5040 18696 5052
rect 18748 5040 18754 5092
rect 19720 5024 19748 5120
rect 18966 4972 18972 5024
rect 19024 5012 19030 5024
rect 19153 5015 19211 5021
rect 19153 5012 19165 5015
rect 19024 4984 19165 5012
rect 19024 4972 19030 4984
rect 19153 4981 19165 4984
rect 19199 4981 19211 5015
rect 19153 4975 19211 4981
rect 19702 4972 19708 5024
rect 19760 5012 19766 5024
rect 19889 5015 19947 5021
rect 19889 5012 19901 5015
rect 19760 4984 19901 5012
rect 19760 4972 19766 4984
rect 19889 4981 19901 4984
rect 19935 4981 19947 5015
rect 19889 4975 19947 4981
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 15746 4808 15752 4820
rect 15707 4780 15752 4808
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 18046 4768 18052 4820
rect 18104 4808 18110 4820
rect 18141 4811 18199 4817
rect 18141 4808 18153 4811
rect 18104 4780 18153 4808
rect 18104 4768 18110 4780
rect 18141 4777 18153 4780
rect 18187 4777 18199 4811
rect 18141 4771 18199 4777
rect 18230 4768 18236 4820
rect 18288 4808 18294 4820
rect 18785 4811 18843 4817
rect 18785 4808 18797 4811
rect 18288 4780 18797 4808
rect 18288 4768 18294 4780
rect 18785 4777 18797 4780
rect 18831 4777 18843 4811
rect 18785 4771 18843 4777
rect 19337 4811 19395 4817
rect 19337 4777 19349 4811
rect 19383 4808 19395 4811
rect 19702 4808 19708 4820
rect 19383 4780 19708 4808
rect 19383 4777 19395 4780
rect 19337 4771 19395 4777
rect 19702 4768 19708 4780
rect 19760 4768 19766 4820
rect 20993 4811 21051 4817
rect 20993 4777 21005 4811
rect 21039 4808 21051 4811
rect 21174 4808 21180 4820
rect 21039 4780 21180 4808
rect 21039 4777 21051 4780
rect 20993 4771 21051 4777
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 14918 4700 14924 4752
rect 14976 4740 14982 4752
rect 20441 4743 20499 4749
rect 20441 4740 20453 4743
rect 14976 4712 20453 4740
rect 14976 4700 14982 4712
rect 20441 4709 20453 4712
rect 20487 4709 20499 4743
rect 20441 4703 20499 4709
rect 14642 4632 14648 4684
rect 14700 4672 14706 4684
rect 15105 4675 15163 4681
rect 15105 4672 15117 4675
rect 14700 4644 15117 4672
rect 14700 4632 14706 4644
rect 15105 4641 15117 4644
rect 15151 4641 15163 4675
rect 15105 4635 15163 4641
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 15930 4672 15936 4684
rect 15335 4644 15936 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 17589 4675 17647 4681
rect 17589 4641 17601 4675
rect 17635 4672 17647 4675
rect 17678 4672 17684 4684
rect 17635 4644 17684 4672
rect 17635 4641 17647 4644
rect 17589 4635 17647 4641
rect 17678 4632 17684 4644
rect 17736 4632 17742 4684
rect 16114 4604 16120 4616
rect 16075 4576 16120 4604
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 18046 4564 18052 4616
rect 18104 4604 18110 4616
rect 20530 4604 20536 4616
rect 18104 4576 20536 4604
rect 18104 4564 18110 4576
rect 20530 4564 20536 4576
rect 20588 4604 20594 4616
rect 20625 4607 20683 4613
rect 20625 4604 20637 4607
rect 20588 4576 20637 4604
rect 20588 4564 20594 4576
rect 20625 4573 20637 4576
rect 20671 4573 20683 4607
rect 20625 4567 20683 4573
rect 15381 4539 15439 4545
rect 15381 4536 15393 4539
rect 14660 4508 15393 4536
rect 12342 4428 12348 4480
rect 12400 4468 12406 4480
rect 14660 4477 14688 4508
rect 15381 4505 15393 4508
rect 15427 4505 15439 4539
rect 15381 4499 15439 4505
rect 16393 4539 16451 4545
rect 16393 4505 16405 4539
rect 16439 4536 16451 4539
rect 17310 4536 17316 4548
rect 16439 4508 17316 4536
rect 16439 4505 16451 4508
rect 16393 4499 16451 4505
rect 17310 4496 17316 4508
rect 17368 4496 17374 4548
rect 17773 4539 17831 4545
rect 17773 4505 17785 4539
rect 17819 4536 17831 4539
rect 18322 4536 18328 4548
rect 17819 4508 18328 4536
rect 17819 4505 17831 4508
rect 17773 4499 17831 4505
rect 18322 4496 18328 4508
rect 18380 4536 18386 4548
rect 18509 4539 18567 4545
rect 18509 4536 18521 4539
rect 18380 4508 18521 4536
rect 18380 4496 18386 4508
rect 18509 4505 18521 4508
rect 18555 4536 18567 4539
rect 18555 4508 20116 4536
rect 18555 4505 18567 4508
rect 18509 4499 18567 4505
rect 14645 4471 14703 4477
rect 14645 4468 14657 4471
rect 12400 4440 14657 4468
rect 12400 4428 12406 4440
rect 14645 4437 14657 4440
rect 14691 4437 14703 4471
rect 14645 4431 14703 4437
rect 16945 4471 17003 4477
rect 16945 4437 16957 4471
rect 16991 4468 17003 4471
rect 17034 4468 17040 4480
rect 16991 4440 17040 4468
rect 16991 4437 17003 4440
rect 16945 4431 17003 4437
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 17402 4428 17408 4480
rect 17460 4468 17466 4480
rect 17681 4471 17739 4477
rect 17681 4468 17693 4471
rect 17460 4440 17693 4468
rect 17460 4428 17466 4440
rect 17681 4437 17693 4440
rect 17727 4468 17739 4471
rect 18966 4468 18972 4480
rect 17727 4440 18972 4468
rect 17727 4437 17739 4440
rect 17681 4431 17739 4437
rect 18966 4428 18972 4440
rect 19024 4428 19030 4480
rect 19610 4468 19616 4480
rect 19571 4440 19616 4468
rect 19610 4428 19616 4440
rect 19668 4428 19674 4480
rect 20088 4477 20116 4508
rect 20073 4471 20131 4477
rect 20073 4437 20085 4471
rect 20119 4468 20131 4471
rect 20162 4468 20168 4480
rect 20119 4440 20168 4468
rect 20119 4437 20131 4440
rect 20073 4431 20131 4437
rect 20162 4428 20168 4440
rect 20220 4428 20226 4480
rect 21358 4468 21364 4480
rect 21319 4440 21364 4468
rect 21358 4428 21364 4440
rect 21416 4428 21422 4480
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 15930 4264 15936 4276
rect 15891 4236 15936 4264
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 17402 4156 17408 4208
rect 17460 4196 17466 4208
rect 18141 4199 18199 4205
rect 18141 4196 18153 4199
rect 17460 4168 18153 4196
rect 17460 4156 17466 4168
rect 18141 4165 18153 4168
rect 18187 4165 18199 4199
rect 18141 4159 18199 4165
rect 19058 4156 19064 4208
rect 19116 4196 19122 4208
rect 19116 4168 19564 4196
rect 19116 4156 19122 4168
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 15194 4128 15200 4140
rect 10376 4100 15200 4128
rect 10376 4088 10382 4100
rect 15194 4088 15200 4100
rect 15252 4088 15258 4140
rect 15378 4088 15384 4140
rect 15436 4128 15442 4140
rect 15436 4100 19288 4128
rect 15436 4088 15442 4100
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 17402 4060 17408 4072
rect 10836 4032 17408 4060
rect 10836 4020 10842 4032
rect 17402 4020 17408 4032
rect 17460 4020 17466 4072
rect 17954 4060 17960 4072
rect 17915 4032 17960 4060
rect 17954 4020 17960 4032
rect 18012 4020 18018 4072
rect 18049 4063 18107 4069
rect 18049 4029 18061 4063
rect 18095 4060 18107 4063
rect 18690 4060 18696 4072
rect 18095 4032 18696 4060
rect 18095 4029 18107 4032
rect 18049 4023 18107 4029
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 19260 4060 19288 4100
rect 19334 4088 19340 4140
rect 19392 4128 19398 4140
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19392 4100 19441 4128
rect 19392 4088 19398 4100
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 19536 4128 19564 4168
rect 19981 4131 20039 4137
rect 19981 4128 19993 4131
rect 19536 4100 19993 4128
rect 19429 4091 19487 4097
rect 19981 4097 19993 4100
rect 20027 4097 20039 4131
rect 20530 4128 20536 4140
rect 20491 4100 20536 4128
rect 19981 4091 20039 4097
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 21085 4131 21143 4137
rect 21085 4097 21097 4131
rect 21131 4128 21143 4131
rect 21450 4128 21456 4140
rect 21131 4100 21456 4128
rect 21131 4097 21143 4100
rect 21085 4091 21143 4097
rect 19260 4032 20392 4060
rect 2498 3952 2504 4004
rect 2556 3992 2562 4004
rect 9214 3992 9220 4004
rect 2556 3964 9220 3992
rect 2556 3952 2562 3964
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 15988 3964 17264 3992
rect 15988 3952 15994 3964
rect 16761 3927 16819 3933
rect 16761 3893 16773 3927
rect 16807 3924 16819 3927
rect 16942 3924 16948 3936
rect 16807 3896 16948 3924
rect 16807 3893 16819 3896
rect 16761 3887 16819 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17126 3924 17132 3936
rect 17087 3896 17132 3924
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17236 3924 17264 3964
rect 18414 3952 18420 4004
rect 18472 3992 18478 4004
rect 20364 4001 20392 4032
rect 20438 4020 20444 4072
rect 20496 4060 20502 4072
rect 20898 4060 20904 4072
rect 20496 4032 20904 4060
rect 20496 4020 20502 4032
rect 20898 4020 20904 4032
rect 20956 4020 20962 4072
rect 18509 3995 18567 4001
rect 18509 3992 18521 3995
rect 18472 3964 18521 3992
rect 18472 3952 18478 3964
rect 18509 3961 18521 3964
rect 18555 3961 18567 3995
rect 19245 3995 19303 4001
rect 19245 3992 19257 3995
rect 18509 3955 18567 3961
rect 18616 3964 19257 3992
rect 18616 3924 18644 3964
rect 19245 3961 19257 3964
rect 19291 3961 19303 3995
rect 19245 3955 19303 3961
rect 20349 3995 20407 4001
rect 20349 3961 20361 3995
rect 20395 3961 20407 3995
rect 20349 3955 20407 3961
rect 20530 3952 20536 4004
rect 20588 3992 20594 4004
rect 21100 3992 21128 4091
rect 21450 4088 21456 4100
rect 21508 4088 21514 4140
rect 20588 3964 21128 3992
rect 20588 3952 20594 3964
rect 17236 3896 18644 3924
rect 18877 3927 18935 3933
rect 18877 3893 18889 3927
rect 18923 3924 18935 3927
rect 18966 3924 18972 3936
rect 18923 3896 18972 3924
rect 18923 3893 18935 3896
rect 18877 3887 18935 3893
rect 18966 3884 18972 3896
rect 19024 3924 19030 3936
rect 19518 3924 19524 3936
rect 19024 3896 19524 3924
rect 19024 3884 19030 3896
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 19794 3924 19800 3936
rect 19755 3896 19800 3924
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 19886 3884 19892 3936
rect 19944 3924 19950 3936
rect 20901 3927 20959 3933
rect 20901 3924 20913 3927
rect 19944 3896 20913 3924
rect 19944 3884 19950 3896
rect 20901 3893 20913 3896
rect 20947 3893 20959 3927
rect 20901 3887 20959 3893
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 10962 3720 10968 3732
rect 3936 3692 10968 3720
rect 3936 3680 3942 3692
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 19337 3723 19395 3729
rect 19337 3720 19349 3723
rect 17000 3692 19349 3720
rect 17000 3680 17006 3692
rect 19337 3689 19349 3692
rect 19383 3689 19395 3723
rect 21174 3720 21180 3732
rect 21135 3692 21180 3720
rect 19337 3683 19395 3689
rect 21174 3680 21180 3692
rect 21232 3680 21238 3732
rect 4798 3612 4804 3664
rect 4856 3652 4862 3664
rect 12342 3652 12348 3664
rect 4856 3624 12348 3652
rect 4856 3612 4862 3624
rect 12342 3612 12348 3624
rect 12400 3612 12406 3664
rect 17957 3655 18015 3661
rect 17957 3621 17969 3655
rect 18003 3652 18015 3655
rect 18138 3652 18144 3664
rect 18003 3624 18144 3652
rect 18003 3621 18015 3624
rect 17957 3615 18015 3621
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 18598 3612 18604 3664
rect 18656 3652 18662 3664
rect 19889 3655 19947 3661
rect 19889 3652 19901 3655
rect 18656 3624 19901 3652
rect 18656 3612 18662 3624
rect 19889 3621 19901 3624
rect 19935 3621 19947 3655
rect 19889 3615 19947 3621
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 17034 3584 17040 3596
rect 8536 3556 17040 3584
rect 8536 3544 8542 3556
rect 17034 3544 17040 3556
rect 17092 3544 17098 3596
rect 18690 3584 18696 3596
rect 18651 3556 18696 3584
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 20254 3584 20260 3596
rect 19536 3556 20260 3584
rect 19536 3528 19564 3556
rect 20254 3544 20260 3556
rect 20312 3544 20318 3596
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3418 3516 3424 3528
rect 2832 3488 3424 3516
rect 2832 3476 2838 3488
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 15562 3516 15568 3528
rect 9456 3488 15568 3516
rect 9456 3476 9462 3488
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 16666 3516 16672 3528
rect 16627 3488 16672 3516
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3516 17003 3519
rect 17126 3516 17132 3528
rect 16991 3488 17132 3516
rect 16991 3485 17003 3488
rect 16945 3479 17003 3485
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 17310 3516 17316 3528
rect 17271 3488 17316 3516
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 19334 3516 19340 3528
rect 17460 3488 19340 3516
rect 17460 3476 17466 3488
rect 19334 3476 19340 3488
rect 19392 3476 19398 3528
rect 19518 3516 19524 3528
rect 19431 3488 19524 3516
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 19610 3476 19616 3528
rect 19668 3516 19674 3528
rect 20070 3516 20076 3528
rect 19668 3488 20076 3516
rect 19668 3476 19674 3488
rect 20070 3476 20076 3488
rect 20128 3476 20134 3528
rect 20162 3476 20168 3528
rect 20220 3516 20226 3528
rect 20901 3519 20959 3525
rect 20901 3516 20913 3519
rect 20220 3488 20913 3516
rect 20220 3476 20226 3488
rect 20901 3485 20913 3488
rect 20947 3516 20959 3519
rect 22094 3516 22100 3528
rect 20947 3488 22100 3516
rect 20947 3485 20959 3488
rect 20901 3479 20959 3485
rect 22094 3476 22100 3488
rect 22152 3476 22158 3528
rect 2038 3408 2044 3460
rect 2096 3448 2102 3460
rect 2096 3420 6914 3448
rect 2096 3408 2102 3420
rect 6886 3380 6914 3420
rect 7558 3408 7564 3460
rect 7616 3448 7622 3460
rect 13538 3448 13544 3460
rect 7616 3420 13544 3448
rect 7616 3408 7622 3420
rect 13538 3408 13544 3420
rect 13596 3408 13602 3460
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 19794 3448 19800 3460
rect 16356 3420 19800 3448
rect 16356 3408 16362 3420
rect 19794 3408 19800 3420
rect 19852 3408 19858 3460
rect 9766 3380 9772 3392
rect 6886 3352 9772 3380
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 9858 3340 9864 3392
rect 9916 3380 9922 3392
rect 15102 3380 15108 3392
rect 9916 3352 15108 3380
rect 9916 3340 9922 3352
rect 15102 3340 15108 3352
rect 15160 3340 15166 3392
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 17497 3383 17555 3389
rect 17497 3380 17509 3383
rect 17276 3352 17509 3380
rect 17276 3340 17282 3352
rect 17497 3349 17509 3352
rect 17543 3349 17555 3383
rect 17497 3343 17555 3349
rect 17954 3340 17960 3392
rect 18012 3380 18018 3392
rect 18322 3380 18328 3392
rect 18012 3352 18328 3380
rect 18012 3340 18018 3352
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 20717 3383 20775 3389
rect 20717 3380 20729 3383
rect 19392 3352 20729 3380
rect 19392 3340 19398 3352
rect 20717 3349 20729 3352
rect 20763 3349 20775 3383
rect 20717 3343 20775 3349
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 13722 3176 13728 3188
rect 8076 3148 13728 3176
rect 8076 3136 8082 3148
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 14274 3136 14280 3188
rect 14332 3176 14338 3188
rect 17034 3176 17040 3188
rect 14332 3148 17040 3176
rect 14332 3136 14338 3148
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 17313 3179 17371 3185
rect 17313 3145 17325 3179
rect 17359 3176 17371 3179
rect 17402 3176 17408 3188
rect 17359 3148 17408 3176
rect 17359 3145 17371 3148
rect 17313 3139 17371 3145
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 18046 3176 18052 3188
rect 18007 3148 18052 3176
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 18138 3136 18144 3188
rect 18196 3176 18202 3188
rect 20257 3179 20315 3185
rect 20257 3176 20269 3179
rect 18196 3148 20269 3176
rect 18196 3136 18202 3148
rect 20257 3145 20269 3148
rect 20303 3145 20315 3179
rect 20257 3139 20315 3145
rect 12158 3068 12164 3120
rect 12216 3108 12222 3120
rect 19150 3108 19156 3120
rect 12216 3080 19156 3108
rect 12216 3068 12222 3080
rect 19150 3068 19156 3080
rect 19208 3068 19214 3120
rect 19426 3068 19432 3120
rect 19484 3108 19490 3120
rect 19978 3108 19984 3120
rect 19484 3080 19984 3108
rect 19484 3068 19490 3080
rect 12894 3040 12900 3052
rect 12855 3012 12900 3040
rect 12894 3000 12900 3012
rect 12952 3000 12958 3052
rect 13446 3040 13452 3052
rect 13407 3012 13452 3040
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 16022 3040 16028 3052
rect 15983 3012 16028 3040
rect 16022 3000 16028 3012
rect 16080 3000 16086 3052
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3040 17739 3043
rect 17770 3040 17776 3052
rect 17727 3012 17776 3040
rect 17727 3009 17739 3012
rect 17681 3003 17739 3009
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3040 18475 3043
rect 19058 3040 19064 3052
rect 18463 3012 19064 3040
rect 18463 3009 18475 3012
rect 18417 3003 18475 3009
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 19334 3040 19340 3052
rect 19295 3012 19340 3040
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 19904 3049 19932 3080
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 19889 3043 19947 3049
rect 19889 3009 19901 3043
rect 19935 3009 19947 3043
rect 20346 3040 20352 3052
rect 19889 3003 19947 3009
rect 19996 3012 20352 3040
rect 14458 2932 14464 2984
rect 14516 2972 14522 2984
rect 16666 2972 16672 2984
rect 14516 2944 16672 2972
rect 14516 2932 14522 2944
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 16945 2975 17003 2981
rect 16945 2941 16957 2975
rect 16991 2972 17003 2975
rect 19996 2972 20024 3012
rect 20346 3000 20352 3012
rect 20404 3040 20410 3052
rect 20441 3043 20499 3049
rect 20441 3040 20453 3043
rect 20404 3012 20453 3040
rect 20404 3000 20410 3012
rect 20441 3009 20453 3012
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 20622 3000 20628 3052
rect 20680 3040 20686 3052
rect 21085 3043 21143 3049
rect 21085 3040 21097 3043
rect 20680 3012 21097 3040
rect 20680 3000 20686 3012
rect 21085 3009 21097 3012
rect 21131 3009 21143 3043
rect 21085 3003 21143 3009
rect 16991 2944 20024 2972
rect 16991 2941 17003 2944
rect 16945 2935 17003 2941
rect 20254 2932 20260 2984
rect 20312 2972 20318 2984
rect 20640 2972 20668 3000
rect 20312 2944 20668 2972
rect 20312 2932 20318 2944
rect 11698 2864 11704 2916
rect 11756 2904 11762 2916
rect 13265 2907 13323 2913
rect 13265 2904 13277 2907
rect 11756 2876 13277 2904
rect 11756 2864 11762 2876
rect 13265 2873 13277 2876
rect 13311 2873 13323 2907
rect 13265 2867 13323 2873
rect 13538 2864 13544 2916
rect 13596 2904 13602 2916
rect 15841 2907 15899 2913
rect 15841 2904 15853 2907
rect 13596 2876 15853 2904
rect 13596 2864 13602 2876
rect 15841 2873 15853 2876
rect 15887 2873 15899 2907
rect 15841 2867 15899 2873
rect 17678 2864 17684 2916
rect 17736 2904 17742 2916
rect 19705 2907 19763 2913
rect 19705 2904 19717 2907
rect 17736 2876 19717 2904
rect 17736 2864 17742 2876
rect 19705 2873 19717 2876
rect 19751 2873 19763 2907
rect 19705 2867 19763 2873
rect 19978 2864 19984 2916
rect 20036 2904 20042 2916
rect 20901 2907 20959 2913
rect 20901 2904 20913 2907
rect 20036 2876 20913 2904
rect 20036 2864 20042 2876
rect 20901 2873 20913 2876
rect 20947 2873 20959 2907
rect 20901 2867 20959 2873
rect 12618 2796 12624 2848
rect 12676 2836 12682 2848
rect 12713 2839 12771 2845
rect 12713 2836 12725 2839
rect 12676 2808 12725 2836
rect 12676 2796 12682 2808
rect 12713 2805 12725 2808
rect 12759 2805 12771 2839
rect 12713 2799 12771 2805
rect 13078 2796 13084 2848
rect 13136 2836 13142 2848
rect 15194 2836 15200 2848
rect 13136 2808 15200 2836
rect 13136 2796 13142 2808
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 18782 2836 18788 2848
rect 18743 2808 18788 2836
rect 18782 2796 18788 2808
rect 18840 2796 18846 2848
rect 19150 2836 19156 2848
rect 19111 2808 19156 2836
rect 19150 2796 19156 2808
rect 19208 2796 19214 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 15194 2592 15200 2644
rect 15252 2632 15258 2644
rect 19613 2635 19671 2641
rect 19613 2632 19625 2635
rect 15252 2604 19625 2632
rect 15252 2592 15258 2604
rect 19613 2601 19625 2604
rect 19659 2601 19671 2635
rect 19613 2595 19671 2601
rect 19702 2592 19708 2644
rect 19760 2632 19766 2644
rect 20901 2635 20959 2641
rect 20901 2632 20913 2635
rect 19760 2604 20913 2632
rect 19760 2592 19766 2604
rect 20901 2601 20913 2604
rect 20947 2601 20959 2635
rect 20901 2595 20959 2601
rect 19058 2524 19064 2576
rect 19116 2564 19122 2576
rect 20349 2567 20407 2573
rect 20349 2564 20361 2567
rect 19116 2536 20361 2564
rect 19116 2524 19122 2536
rect 20349 2533 20361 2536
rect 20395 2533 20407 2567
rect 20349 2527 20407 2533
rect 17405 2499 17463 2505
rect 17405 2465 17417 2499
rect 17451 2496 17463 2499
rect 20254 2496 20260 2508
rect 17451 2468 20260 2496
rect 17451 2465 17463 2468
rect 17405 2459 17463 2465
rect 20254 2456 20260 2468
rect 20312 2456 20318 2508
rect 22370 2496 22376 2508
rect 20364 2468 22376 2496
rect 18509 2431 18567 2437
rect 18509 2397 18521 2431
rect 18555 2428 18567 2431
rect 19610 2428 19616 2440
rect 18555 2400 19616 2428
rect 18555 2397 18567 2400
rect 18509 2391 18567 2397
rect 19610 2388 19616 2400
rect 19668 2388 19674 2440
rect 19794 2388 19800 2440
rect 19852 2428 19858 2440
rect 20364 2428 20392 2468
rect 22370 2456 22376 2468
rect 22428 2456 22434 2508
rect 19852 2400 20392 2428
rect 20533 2431 20591 2437
rect 19852 2388 19858 2400
rect 20533 2397 20545 2431
rect 20579 2428 20591 2431
rect 20990 2428 20996 2440
rect 20579 2400 20996 2428
rect 20579 2397 20591 2400
rect 20533 2391 20591 2397
rect 17773 2363 17831 2369
rect 17773 2329 17785 2363
rect 17819 2360 17831 2363
rect 20548 2360 20576 2391
rect 20990 2388 20996 2400
rect 21048 2388 21054 2440
rect 21082 2388 21088 2440
rect 21140 2428 21146 2440
rect 21140 2400 21185 2428
rect 21140 2388 21146 2400
rect 17819 2332 20576 2360
rect 17819 2329 17831 2332
rect 17773 2323 17831 2329
rect 17037 2295 17095 2301
rect 17037 2261 17049 2295
rect 17083 2292 17095 2295
rect 17954 2292 17960 2304
rect 17083 2264 17960 2292
rect 17083 2261 17095 2264
rect 17037 2255 17095 2261
rect 17954 2252 17960 2264
rect 18012 2252 18018 2304
rect 18141 2295 18199 2301
rect 18141 2261 18153 2295
rect 18187 2292 18199 2295
rect 18230 2292 18236 2304
rect 18187 2264 18236 2292
rect 18187 2261 18199 2264
rect 18141 2255 18199 2261
rect 18230 2252 18236 2264
rect 18288 2252 18294 2304
rect 18877 2295 18935 2301
rect 18877 2261 18889 2295
rect 18923 2292 18935 2295
rect 19334 2292 19340 2304
rect 18923 2264 19340 2292
rect 18923 2261 18935 2264
rect 18877 2255 18935 2261
rect 19334 2252 19340 2264
rect 19392 2252 19398 2304
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 5534 2048 5540 2100
rect 5592 2088 5598 2100
rect 6178 2088 6184 2100
rect 5592 2060 6184 2088
rect 5592 2048 5598 2060
rect 6178 2048 6184 2060
rect 6236 2048 6242 2100
rect 17954 2048 17960 2100
rect 18012 2088 18018 2100
rect 21082 2088 21088 2100
rect 18012 2060 21088 2088
rect 18012 2048 18018 2060
rect 21082 2048 21088 2060
rect 21140 2048 21146 2100
rect 18230 1980 18236 2032
rect 18288 2020 18294 2032
rect 19794 2020 19800 2032
rect 18288 1992 19800 2020
rect 18288 1980 18294 1992
rect 19794 1980 19800 1992
rect 19852 1980 19858 2032
<< via1 >>
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 21180 20587 21232 20596
rect 18880 20476 18932 20528
rect 17040 20408 17092 20460
rect 16212 20340 16264 20392
rect 19708 20408 19760 20460
rect 21180 20553 21189 20587
rect 21189 20553 21223 20587
rect 21223 20553 21232 20587
rect 21180 20544 21232 20553
rect 17500 20383 17552 20392
rect 17500 20349 17509 20383
rect 17509 20349 17543 20383
rect 17543 20349 17552 20383
rect 17500 20340 17552 20349
rect 20720 20383 20772 20392
rect 20720 20349 20729 20383
rect 20729 20349 20763 20383
rect 20763 20349 20772 20383
rect 20720 20340 20772 20349
rect 18972 20204 19024 20256
rect 19524 20204 19576 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 6552 20043 6604 20052
rect 6552 20009 6561 20043
rect 6561 20009 6595 20043
rect 6595 20009 6604 20043
rect 6552 20000 6604 20009
rect 16212 20000 16264 20052
rect 5172 19975 5224 19984
rect 5172 19941 5181 19975
rect 5181 19941 5215 19975
rect 5215 19941 5224 19975
rect 5172 19932 5224 19941
rect 10968 19932 11020 19984
rect 9864 19839 9916 19848
rect 5908 19771 5960 19780
rect 5908 19737 5917 19771
rect 5917 19737 5951 19771
rect 5951 19737 5960 19771
rect 5908 19728 5960 19737
rect 4068 19703 4120 19712
rect 4068 19669 4077 19703
rect 4077 19669 4111 19703
rect 4111 19669 4120 19703
rect 4068 19660 4120 19669
rect 9588 19660 9640 19712
rect 9864 19805 9873 19839
rect 9873 19805 9907 19839
rect 9907 19805 9916 19839
rect 9864 19796 9916 19805
rect 11704 19839 11756 19848
rect 11704 19805 11713 19839
rect 11713 19805 11747 19839
rect 11747 19805 11756 19839
rect 11704 19796 11756 19805
rect 17500 19796 17552 19848
rect 18052 19839 18104 19848
rect 18052 19805 18061 19839
rect 18061 19805 18095 19839
rect 18095 19805 18104 19839
rect 18052 19796 18104 19805
rect 18880 19839 18932 19848
rect 18880 19805 18889 19839
rect 18889 19805 18923 19839
rect 18923 19805 18932 19839
rect 18880 19796 18932 19805
rect 20720 19796 20772 19848
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 15108 19728 15160 19780
rect 15292 19728 15344 19780
rect 16396 19728 16448 19780
rect 11244 19660 11296 19712
rect 14556 19660 14608 19712
rect 14924 19660 14976 19712
rect 18328 19728 18380 19780
rect 20260 19728 20312 19780
rect 20628 19660 20680 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 9680 19456 9732 19508
rect 10140 19456 10192 19508
rect 10048 19363 10100 19372
rect 10048 19329 10057 19363
rect 10057 19329 10091 19363
rect 10091 19329 10100 19363
rect 10048 19320 10100 19329
rect 11244 19456 11296 19508
rect 15844 19456 15896 19508
rect 18144 19456 18196 19508
rect 18328 19499 18380 19508
rect 18328 19465 18337 19499
rect 18337 19465 18371 19499
rect 18371 19465 18380 19499
rect 18328 19456 18380 19465
rect 19708 19456 19760 19508
rect 10508 19388 10560 19440
rect 14372 19388 14424 19440
rect 14924 19388 14976 19440
rect 10968 19363 11020 19372
rect 10968 19329 10977 19363
rect 10977 19329 11011 19363
rect 11011 19329 11020 19363
rect 10968 19320 11020 19329
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 12900 19320 12952 19372
rect 14648 19363 14700 19372
rect 14648 19329 14682 19363
rect 14682 19329 14700 19363
rect 14648 19320 14700 19329
rect 15108 19320 15160 19372
rect 16948 19363 17000 19372
rect 16948 19329 16982 19363
rect 16982 19329 17000 19363
rect 16948 19320 17000 19329
rect 18052 19388 18104 19440
rect 20720 19388 20772 19440
rect 21088 19363 21140 19372
rect 21088 19329 21106 19363
rect 21106 19329 21140 19363
rect 21088 19320 21140 19329
rect 12440 19184 12492 19236
rect 12532 19116 12584 19168
rect 14280 19252 14332 19304
rect 16580 19252 16632 19304
rect 15384 19116 15436 19168
rect 18236 19116 18288 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 10048 18819 10100 18828
rect 10048 18785 10057 18819
rect 10057 18785 10091 18819
rect 10091 18785 10100 18819
rect 10048 18776 10100 18785
rect 11888 18776 11940 18828
rect 12624 18751 12676 18760
rect 12624 18717 12647 18751
rect 12647 18717 12676 18751
rect 12624 18708 12676 18717
rect 14188 18708 14240 18760
rect 16580 18708 16632 18760
rect 17408 18708 17460 18760
rect 19064 18708 19116 18760
rect 12808 18640 12860 18692
rect 15200 18640 15252 18692
rect 17684 18640 17736 18692
rect 18696 18640 18748 18692
rect 13820 18572 13872 18624
rect 15292 18572 15344 18624
rect 17132 18615 17184 18624
rect 17132 18581 17141 18615
rect 17141 18581 17175 18615
rect 17175 18581 17184 18615
rect 17132 18572 17184 18581
rect 17500 18572 17552 18624
rect 20444 18572 20496 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 13820 18300 13872 18352
rect 14464 18300 14516 18352
rect 14188 18275 14240 18284
rect 14188 18241 14197 18275
rect 14197 18241 14231 18275
rect 14231 18241 14240 18275
rect 14188 18232 14240 18241
rect 17408 18275 17460 18284
rect 17408 18241 17417 18275
rect 17417 18241 17451 18275
rect 17451 18241 17460 18275
rect 17408 18232 17460 18241
rect 15384 18164 15436 18216
rect 16304 18164 16356 18216
rect 20444 18275 20496 18284
rect 20444 18241 20462 18275
rect 20462 18241 20496 18275
rect 20720 18275 20772 18284
rect 20444 18232 20496 18241
rect 20720 18241 20729 18275
rect 20729 18241 20763 18275
rect 20763 18241 20772 18275
rect 20720 18232 20772 18241
rect 10600 18028 10652 18080
rect 12808 18071 12860 18080
rect 12808 18037 12817 18071
rect 12817 18037 12851 18071
rect 12851 18037 12860 18071
rect 12808 18028 12860 18037
rect 18788 18071 18840 18080
rect 18788 18037 18797 18071
rect 18797 18037 18831 18071
rect 18831 18037 18840 18071
rect 18788 18028 18840 18037
rect 19616 18028 19668 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 16396 17867 16448 17876
rect 16396 17833 16405 17867
rect 16405 17833 16439 17867
rect 16439 17833 16448 17867
rect 16396 17824 16448 17833
rect 17408 17824 17460 17876
rect 17960 17688 18012 17740
rect 17500 17663 17552 17672
rect 17500 17629 17518 17663
rect 17518 17629 17552 17663
rect 17500 17620 17552 17629
rect 19524 17620 19576 17672
rect 20720 17620 20772 17672
rect 16948 17552 17000 17604
rect 18420 17552 18472 17604
rect 18972 17552 19024 17604
rect 21364 17484 21416 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 11704 17280 11756 17332
rect 14648 17280 14700 17332
rect 17684 17323 17736 17332
rect 17684 17289 17693 17323
rect 17693 17289 17727 17323
rect 17727 17289 17736 17323
rect 17684 17280 17736 17289
rect 19432 17280 19484 17332
rect 19892 17280 19944 17332
rect 14556 17255 14608 17264
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 12348 17144 12400 17196
rect 13820 17144 13872 17196
rect 14556 17221 14590 17255
rect 14590 17221 14608 17255
rect 14556 17212 14608 17221
rect 18328 17212 18380 17264
rect 18788 17255 18840 17264
rect 18788 17221 18806 17255
rect 18806 17221 18840 17255
rect 18788 17212 18840 17221
rect 20720 17212 20772 17264
rect 14372 17144 14424 17196
rect 19064 17187 19116 17196
rect 19064 17153 19073 17187
rect 19073 17153 19107 17187
rect 19107 17153 19116 17187
rect 19064 17144 19116 17153
rect 21180 17144 21232 17196
rect 11980 17119 12032 17128
rect 11980 17085 11989 17119
rect 11989 17085 12023 17119
rect 12023 17085 12032 17119
rect 11980 17076 12032 17085
rect 14556 16940 14608 16992
rect 15384 16940 15436 16992
rect 20904 16940 20956 16992
rect 21088 16940 21140 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 11888 16643 11940 16652
rect 11888 16609 11897 16643
rect 11897 16609 11931 16643
rect 11931 16609 11940 16643
rect 11888 16600 11940 16609
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 17960 16736 18012 16788
rect 18236 16736 18288 16788
rect 22468 16736 22520 16788
rect 12440 16532 12492 16584
rect 12716 16464 12768 16516
rect 13820 16396 13872 16448
rect 14372 16532 14424 16584
rect 18236 16532 18288 16584
rect 19064 16532 19116 16584
rect 19524 16532 19576 16584
rect 19984 16532 20036 16584
rect 15384 16507 15436 16516
rect 15384 16473 15418 16507
rect 15418 16473 15436 16507
rect 15384 16464 15436 16473
rect 16948 16464 17000 16516
rect 16120 16396 16172 16448
rect 18696 16396 18748 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 9864 16235 9916 16244
rect 9864 16201 9873 16235
rect 9873 16201 9907 16235
rect 9907 16201 9916 16235
rect 9864 16192 9916 16201
rect 13728 16192 13780 16244
rect 13820 16192 13872 16244
rect 14924 16192 14976 16244
rect 16304 16192 16356 16244
rect 15292 16124 15344 16176
rect 15568 16124 15620 16176
rect 19524 16124 19576 16176
rect 13820 16056 13872 16108
rect 14372 16099 14424 16108
rect 14372 16065 14381 16099
rect 14381 16065 14415 16099
rect 14415 16065 14424 16099
rect 14372 16056 14424 16065
rect 15108 16056 15160 16108
rect 17960 16056 18012 16108
rect 20444 16056 20496 16108
rect 10600 15988 10652 16040
rect 19064 15988 19116 16040
rect 15292 15852 15344 15904
rect 15660 15852 15712 15904
rect 21180 15895 21232 15904
rect 21180 15861 21189 15895
rect 21189 15861 21223 15895
rect 21223 15861 21232 15895
rect 21180 15852 21232 15861
rect 21548 15852 21600 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 17960 15512 18012 15564
rect 19064 15444 19116 15496
rect 19616 15444 19668 15496
rect 16120 15376 16172 15428
rect 15108 15351 15160 15360
rect 15108 15317 15117 15351
rect 15117 15317 15151 15351
rect 15151 15317 15160 15351
rect 15108 15308 15160 15317
rect 19616 15308 19668 15360
rect 19892 15308 19944 15360
rect 21272 15308 21324 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 10140 15147 10192 15156
rect 10140 15113 10149 15147
rect 10149 15113 10183 15147
rect 10183 15113 10192 15147
rect 10140 15104 10192 15113
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 12256 14968 12308 15020
rect 12440 14968 12492 15020
rect 14372 15011 14424 15020
rect 14372 14977 14381 15011
rect 14381 14977 14415 15011
rect 14415 14977 14424 15011
rect 14372 14968 14424 14977
rect 15476 14968 15528 15020
rect 20720 14968 20772 15020
rect 21364 14968 21416 15020
rect 12532 14900 12584 14952
rect 20812 14943 20864 14952
rect 20812 14909 20821 14943
rect 20821 14909 20855 14943
rect 20855 14909 20864 14943
rect 20812 14900 20864 14909
rect 12716 14764 12768 14816
rect 17868 14764 17920 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 10232 14603 10284 14612
rect 10232 14569 10241 14603
rect 10241 14569 10275 14603
rect 10275 14569 10284 14603
rect 10232 14560 10284 14569
rect 15108 14560 15160 14612
rect 16304 14535 16356 14544
rect 16304 14501 16313 14535
rect 16313 14501 16347 14535
rect 16347 14501 16356 14535
rect 16304 14492 16356 14501
rect 10508 14467 10560 14476
rect 10508 14433 10517 14467
rect 10517 14433 10551 14467
rect 10551 14433 10560 14467
rect 10508 14424 10560 14433
rect 15476 14467 15528 14476
rect 15476 14433 15485 14467
rect 15485 14433 15519 14467
rect 15519 14433 15528 14467
rect 15476 14424 15528 14433
rect 12992 14356 13044 14408
rect 16304 14356 16356 14408
rect 19064 14356 19116 14408
rect 20812 14356 20864 14408
rect 21364 14356 21416 14408
rect 9220 14263 9272 14272
rect 9220 14229 9229 14263
rect 9229 14229 9263 14263
rect 9263 14229 9272 14263
rect 9220 14220 9272 14229
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 13268 14220 13320 14272
rect 15200 14331 15252 14340
rect 15200 14297 15218 14331
rect 15218 14297 15252 14331
rect 15200 14288 15252 14297
rect 15660 14288 15712 14340
rect 17868 14288 17920 14340
rect 18144 14288 18196 14340
rect 18604 14220 18656 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 12440 14059 12492 14068
rect 12440 14025 12449 14059
rect 12449 14025 12483 14059
rect 12483 14025 12492 14059
rect 12440 14016 12492 14025
rect 13820 14016 13872 14068
rect 14372 14016 14424 14068
rect 14832 14016 14884 14068
rect 17132 14016 17184 14068
rect 18144 14016 18196 14068
rect 20444 14016 20496 14068
rect 12992 13948 13044 14000
rect 16948 13991 17000 14000
rect 16948 13957 16982 13991
rect 16982 13957 17000 13991
rect 16948 13948 17000 13957
rect 14832 13880 14884 13932
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 15660 13880 15712 13932
rect 19064 13948 19116 14000
rect 18604 13923 18656 13932
rect 18604 13889 18638 13923
rect 18638 13889 18656 13923
rect 18604 13880 18656 13889
rect 21272 13880 21324 13932
rect 21364 13855 21416 13864
rect 21364 13821 21373 13855
rect 21373 13821 21407 13855
rect 21407 13821 21416 13855
rect 21364 13812 21416 13821
rect 22008 13812 22060 13864
rect 22560 13812 22612 13864
rect 13820 13744 13872 13796
rect 19708 13719 19760 13728
rect 19708 13685 19717 13719
rect 19717 13685 19751 13719
rect 19751 13685 19760 13719
rect 19708 13676 19760 13685
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 13820 13472 13872 13524
rect 14740 13472 14792 13524
rect 21088 13515 21140 13524
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 15200 13200 15252 13252
rect 21088 13481 21097 13515
rect 21097 13481 21131 13515
rect 21131 13481 21140 13515
rect 21088 13472 21140 13481
rect 19064 13336 19116 13388
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 17224 13200 17276 13252
rect 12808 13132 12860 13184
rect 17316 13132 17368 13184
rect 19708 13200 19760 13252
rect 20076 13200 20128 13252
rect 21088 13132 21140 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 11060 12928 11112 12980
rect 12808 12928 12860 12980
rect 14556 12928 14608 12980
rect 14740 12971 14792 12980
rect 14740 12937 14749 12971
rect 14749 12937 14783 12971
rect 14783 12937 14792 12971
rect 14740 12928 14792 12937
rect 12440 12860 12492 12912
rect 12992 12835 13044 12844
rect 5540 12656 5592 12708
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 13268 12835 13320 12844
rect 13268 12801 13302 12835
rect 13302 12801 13320 12835
rect 13268 12792 13320 12801
rect 13544 12792 13596 12844
rect 19524 12928 19576 12980
rect 19892 12928 19944 12980
rect 15660 12860 15712 12912
rect 21088 12903 21140 12912
rect 21088 12869 21106 12903
rect 21106 12869 21140 12903
rect 21088 12860 21140 12869
rect 12532 12588 12584 12640
rect 15016 12588 15068 12640
rect 19064 12792 19116 12844
rect 21364 12835 21416 12844
rect 21364 12801 21373 12835
rect 21373 12801 21407 12835
rect 21407 12801 21416 12835
rect 21364 12792 21416 12801
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 18696 12427 18748 12436
rect 18696 12393 18705 12427
rect 18705 12393 18739 12427
rect 18739 12393 18748 12427
rect 18696 12384 18748 12393
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 20536 12427 20588 12436
rect 20536 12393 20545 12427
rect 20545 12393 20579 12427
rect 20579 12393 20588 12427
rect 20536 12384 20588 12393
rect 21456 12384 21508 12436
rect 13912 12316 13964 12368
rect 14372 12316 14424 12368
rect 13820 12248 13872 12300
rect 15844 12291 15896 12300
rect 15844 12257 15853 12291
rect 15853 12257 15887 12291
rect 15887 12257 15896 12291
rect 15844 12248 15896 12257
rect 12164 12044 12216 12096
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 15568 12044 15620 12096
rect 15752 12044 15804 12096
rect 16120 12087 16172 12096
rect 16120 12053 16129 12087
rect 16129 12053 16163 12087
rect 16163 12053 16172 12087
rect 16120 12044 16172 12053
rect 17132 12044 17184 12096
rect 19524 12180 19576 12232
rect 21272 12248 21324 12300
rect 22192 12248 22244 12300
rect 20444 12180 20496 12232
rect 21272 12112 21324 12164
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 12532 11840 12584 11892
rect 14464 11840 14516 11892
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 16120 11840 16172 11892
rect 17040 11840 17092 11892
rect 18512 11883 18564 11892
rect 18512 11849 18521 11883
rect 18521 11849 18555 11883
rect 18555 11849 18564 11883
rect 18512 11840 18564 11849
rect 20628 11840 20680 11892
rect 14832 11704 14884 11756
rect 17960 11704 18012 11756
rect 18052 11704 18104 11756
rect 20812 11747 20864 11756
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 15292 11679 15344 11688
rect 15292 11645 15301 11679
rect 15301 11645 15335 11679
rect 15335 11645 15344 11679
rect 15292 11636 15344 11645
rect 15384 11636 15436 11688
rect 17592 11679 17644 11688
rect 17592 11645 17601 11679
rect 17601 11645 17635 11679
rect 17635 11645 17644 11679
rect 17592 11636 17644 11645
rect 17684 11679 17736 11688
rect 17684 11645 17693 11679
rect 17693 11645 17727 11679
rect 17727 11645 17736 11679
rect 17684 11636 17736 11645
rect 20812 11713 20821 11747
rect 20821 11713 20855 11747
rect 20855 11713 20864 11747
rect 20812 11704 20864 11713
rect 20720 11636 20772 11688
rect 21456 11568 21508 11620
rect 11612 11500 11664 11552
rect 15200 11500 15252 11552
rect 15844 11500 15896 11552
rect 18696 11500 18748 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 12164 11339 12216 11348
rect 12164 11305 12173 11339
rect 12173 11305 12207 11339
rect 12207 11305 12216 11339
rect 12164 11296 12216 11305
rect 12900 11296 12952 11348
rect 14832 11339 14884 11348
rect 14832 11305 14841 11339
rect 14841 11305 14875 11339
rect 14875 11305 14884 11339
rect 14832 11296 14884 11305
rect 15384 11339 15436 11348
rect 15384 11305 15393 11339
rect 15393 11305 15427 11339
rect 15427 11305 15436 11339
rect 15384 11296 15436 11305
rect 18788 11296 18840 11348
rect 21180 11296 21232 11348
rect 11612 11203 11664 11212
rect 11612 11169 11621 11203
rect 11621 11169 11655 11203
rect 11655 11169 11664 11203
rect 11612 11160 11664 11169
rect 15476 11228 15528 11280
rect 16948 11228 17000 11280
rect 17408 11228 17460 11280
rect 18880 11271 18932 11280
rect 18880 11237 18889 11271
rect 18889 11237 18923 11271
rect 18923 11237 18932 11271
rect 18880 11228 18932 11237
rect 14556 11160 14608 11212
rect 14924 11160 14976 11212
rect 17500 11203 17552 11212
rect 17500 11169 17509 11203
rect 17509 11169 17543 11203
rect 17543 11169 17552 11203
rect 17500 11160 17552 11169
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 18144 11160 18196 11212
rect 18788 11160 18840 11212
rect 12808 11092 12860 11144
rect 14740 11092 14792 11144
rect 20996 11092 21048 11144
rect 6644 11024 6696 11076
rect 12348 11024 12400 11076
rect 15844 11067 15896 11076
rect 15844 11033 15853 11067
rect 15853 11033 15887 11067
rect 15887 11033 15896 11067
rect 15844 11024 15896 11033
rect 17040 11024 17092 11076
rect 12716 10956 12768 11008
rect 15568 10956 15620 11008
rect 16948 10999 17000 11008
rect 16948 10965 16957 10999
rect 16957 10965 16991 10999
rect 16991 10965 17000 10999
rect 16948 10956 17000 10965
rect 18880 11024 18932 11076
rect 19156 11024 19208 11076
rect 20352 11024 20404 11076
rect 21088 11024 21140 11076
rect 21456 11024 21508 11076
rect 18512 10999 18564 11008
rect 18512 10965 18521 10999
rect 18521 10965 18555 10999
rect 18555 10965 18564 10999
rect 18512 10956 18564 10965
rect 18696 10956 18748 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 12256 10752 12308 10804
rect 14740 10752 14792 10804
rect 16948 10752 17000 10804
rect 17592 10752 17644 10804
rect 20168 10795 20220 10804
rect 20168 10761 20177 10795
rect 20177 10761 20211 10795
rect 20211 10761 20220 10795
rect 20168 10752 20220 10761
rect 22100 10752 22152 10804
rect 5816 10684 5868 10736
rect 12348 10727 12400 10736
rect 12348 10693 12357 10727
rect 12357 10693 12391 10727
rect 12391 10693 12400 10727
rect 12348 10684 12400 10693
rect 12440 10616 12492 10668
rect 16580 10684 16632 10736
rect 17040 10727 17092 10736
rect 17040 10693 17049 10727
rect 17049 10693 17083 10727
rect 17083 10693 17092 10727
rect 17040 10684 17092 10693
rect 18144 10684 18196 10736
rect 20352 10684 20404 10736
rect 13728 10616 13780 10668
rect 14832 10616 14884 10668
rect 15936 10616 15988 10668
rect 17132 10616 17184 10668
rect 18512 10616 18564 10668
rect 20720 10616 20772 10668
rect 12716 10591 12768 10600
rect 12716 10557 12725 10591
rect 12725 10557 12759 10591
rect 12759 10557 12768 10591
rect 12716 10548 12768 10557
rect 14280 10591 14332 10600
rect 14280 10557 14289 10591
rect 14289 10557 14323 10591
rect 14323 10557 14332 10591
rect 14280 10548 14332 10557
rect 16396 10548 16448 10600
rect 17960 10548 18012 10600
rect 18328 10591 18380 10600
rect 18052 10480 18104 10532
rect 18328 10557 18337 10591
rect 18337 10557 18371 10591
rect 18371 10557 18380 10591
rect 18328 10548 18380 10557
rect 18420 10548 18472 10600
rect 20260 10591 20312 10600
rect 20260 10557 20269 10591
rect 20269 10557 20303 10591
rect 20303 10557 20312 10591
rect 20260 10548 20312 10557
rect 19156 10480 19208 10532
rect 15476 10455 15528 10464
rect 15476 10421 15485 10455
rect 15485 10421 15519 10455
rect 15519 10421 15528 10455
rect 15476 10412 15528 10421
rect 17500 10412 17552 10464
rect 19708 10455 19760 10464
rect 19708 10421 19717 10455
rect 19717 10421 19751 10455
rect 19751 10421 19760 10455
rect 19708 10412 19760 10421
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 2964 10208 3016 10260
rect 12716 10208 12768 10260
rect 13728 10208 13780 10260
rect 14832 10251 14884 10260
rect 14832 10217 14841 10251
rect 14841 10217 14875 10251
rect 14875 10217 14884 10251
rect 14832 10208 14884 10217
rect 15936 10251 15988 10260
rect 15936 10217 15945 10251
rect 15945 10217 15979 10251
rect 15979 10217 15988 10251
rect 15936 10208 15988 10217
rect 16120 10208 16172 10260
rect 19708 10208 19760 10260
rect 20168 10208 20220 10260
rect 22560 10208 22612 10260
rect 11980 10140 12032 10192
rect 15660 10140 15712 10192
rect 16580 10140 16632 10192
rect 17592 10140 17644 10192
rect 15016 10072 15068 10124
rect 16304 10072 16356 10124
rect 17500 10115 17552 10124
rect 17500 10081 17509 10115
rect 17509 10081 17543 10115
rect 17543 10081 17552 10115
rect 17500 10072 17552 10081
rect 20628 10140 20680 10192
rect 17960 10072 18012 10124
rect 18420 10072 18472 10124
rect 20444 10072 20496 10124
rect 22008 10072 22060 10124
rect 22376 10072 22428 10124
rect 12440 10004 12492 10056
rect 19248 10047 19300 10056
rect 2780 9868 2832 9920
rect 19248 10013 19257 10047
rect 19257 10013 19291 10047
rect 19291 10013 19300 10047
rect 19248 10004 19300 10013
rect 15568 9979 15620 9988
rect 15568 9945 15577 9979
rect 15577 9945 15611 9979
rect 15611 9945 15620 9979
rect 15568 9936 15620 9945
rect 18328 9936 18380 9988
rect 13360 9868 13412 9920
rect 14372 9911 14424 9920
rect 14372 9877 14381 9911
rect 14381 9877 14415 9911
rect 14415 9877 14424 9911
rect 14372 9868 14424 9877
rect 16304 9911 16356 9920
rect 16304 9877 16313 9911
rect 16313 9877 16347 9911
rect 16347 9877 16356 9911
rect 16304 9868 16356 9877
rect 16396 9911 16448 9920
rect 16396 9877 16405 9911
rect 16405 9877 16439 9911
rect 16439 9877 16448 9911
rect 17040 9911 17092 9920
rect 16396 9868 16448 9877
rect 17040 9877 17049 9911
rect 17049 9877 17083 9911
rect 17083 9877 17092 9911
rect 17040 9868 17092 9877
rect 18512 9911 18564 9920
rect 18512 9877 18521 9911
rect 18521 9877 18555 9911
rect 18555 9877 18564 9911
rect 18512 9868 18564 9877
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 4344 9664 4396 9716
rect 13728 9664 13780 9716
rect 15476 9664 15528 9716
rect 13360 9596 13412 9648
rect 7104 9324 7156 9376
rect 13544 9460 13596 9512
rect 15200 9596 15252 9648
rect 16304 9596 16356 9648
rect 18328 9596 18380 9648
rect 20904 9596 20956 9648
rect 21364 9639 21416 9648
rect 21364 9605 21373 9639
rect 21373 9605 21407 9639
rect 21407 9605 21416 9639
rect 21364 9596 21416 9605
rect 17684 9528 17736 9580
rect 20444 9528 20496 9580
rect 12808 9435 12860 9444
rect 12808 9401 12817 9435
rect 12817 9401 12851 9435
rect 12851 9401 12860 9435
rect 12808 9392 12860 9401
rect 13728 9392 13780 9444
rect 15476 9460 15528 9512
rect 18880 9460 18932 9512
rect 16396 9392 16448 9444
rect 19248 9392 19300 9444
rect 13360 9367 13412 9376
rect 13360 9333 13369 9367
rect 13369 9333 13403 9367
rect 13403 9333 13412 9367
rect 13360 9324 13412 9333
rect 17500 9367 17552 9376
rect 17500 9333 17509 9367
rect 17509 9333 17543 9367
rect 17543 9333 17552 9367
rect 17500 9324 17552 9333
rect 18144 9324 18196 9376
rect 19892 9503 19944 9512
rect 19892 9469 19901 9503
rect 19901 9469 19935 9503
rect 19935 9469 19944 9503
rect 19892 9460 19944 9469
rect 19892 9324 19944 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 11244 9120 11296 9172
rect 17500 9120 17552 9172
rect 16212 8984 16264 9036
rect 20076 9052 20128 9104
rect 20812 8984 20864 9036
rect 16120 8916 16172 8968
rect 16948 8848 17000 8900
rect 14556 8823 14608 8832
rect 14556 8789 14565 8823
rect 14565 8789 14599 8823
rect 14599 8789 14608 8823
rect 14556 8780 14608 8789
rect 15200 8780 15252 8832
rect 17316 8780 17368 8832
rect 17868 8780 17920 8832
rect 18144 8823 18196 8832
rect 18144 8789 18153 8823
rect 18153 8789 18187 8823
rect 18187 8789 18196 8823
rect 18144 8780 18196 8789
rect 20076 8916 20128 8968
rect 21364 8916 21416 8968
rect 20996 8848 21048 8900
rect 20904 8823 20956 8832
rect 20904 8789 20913 8823
rect 20913 8789 20947 8823
rect 20947 8789 20956 8823
rect 20904 8780 20956 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 14556 8619 14608 8628
rect 14556 8585 14565 8619
rect 14565 8585 14599 8619
rect 14599 8585 14608 8619
rect 14556 8576 14608 8585
rect 17132 8619 17184 8628
rect 17132 8585 17141 8619
rect 17141 8585 17175 8619
rect 17175 8585 17184 8619
rect 17684 8619 17736 8628
rect 17132 8576 17184 8585
rect 17684 8585 17693 8619
rect 17693 8585 17727 8619
rect 17727 8585 17736 8619
rect 17684 8576 17736 8585
rect 17776 8576 17828 8628
rect 20444 8619 20496 8628
rect 20444 8585 20453 8619
rect 20453 8585 20487 8619
rect 20487 8585 20496 8619
rect 20444 8576 20496 8585
rect 21640 8576 21692 8628
rect 13820 8508 13872 8560
rect 5264 8372 5316 8424
rect 14556 8372 14608 8424
rect 9128 8304 9180 8356
rect 16028 8440 16080 8492
rect 17316 8440 17368 8492
rect 18328 8440 18380 8492
rect 20168 8440 20220 8492
rect 21088 8440 21140 8492
rect 16948 8304 17000 8356
rect 17960 8372 18012 8424
rect 18236 8415 18288 8424
rect 18236 8381 18245 8415
rect 18245 8381 18279 8415
rect 18279 8381 18288 8415
rect 19800 8415 19852 8424
rect 18236 8372 18288 8381
rect 19800 8381 19809 8415
rect 19809 8381 19843 8415
rect 19843 8381 19852 8415
rect 19800 8372 19852 8381
rect 19984 8415 20036 8424
rect 19984 8381 19993 8415
rect 19993 8381 20027 8415
rect 20027 8381 20036 8415
rect 19984 8372 20036 8381
rect 18604 8304 18656 8356
rect 18880 8304 18932 8356
rect 16764 8236 16816 8288
rect 18696 8279 18748 8288
rect 18696 8245 18705 8279
rect 18705 8245 18739 8279
rect 18739 8245 18748 8279
rect 18696 8236 18748 8245
rect 20996 8236 21048 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 14372 8032 14424 8084
rect 18144 8032 18196 8084
rect 19984 8032 20036 8084
rect 13268 7896 13320 7948
rect 16028 7896 16080 7948
rect 18604 7896 18656 7948
rect 19524 7939 19576 7948
rect 19524 7905 19533 7939
rect 19533 7905 19567 7939
rect 19567 7905 19576 7939
rect 19524 7896 19576 7905
rect 21180 7896 21232 7948
rect 5724 7828 5776 7880
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 18328 7828 18380 7880
rect 19064 7828 19116 7880
rect 5632 7735 5684 7744
rect 5632 7701 5641 7735
rect 5641 7701 5675 7735
rect 5675 7701 5684 7735
rect 5632 7692 5684 7701
rect 13544 7692 13596 7744
rect 18236 7760 18288 7812
rect 18788 7760 18840 7812
rect 21088 7760 21140 7812
rect 15292 7692 15344 7744
rect 15568 7735 15620 7744
rect 15568 7701 15577 7735
rect 15577 7701 15611 7735
rect 15611 7701 15620 7735
rect 15568 7692 15620 7701
rect 18144 7692 18196 7744
rect 18696 7735 18748 7744
rect 18696 7701 18705 7735
rect 18705 7701 18739 7735
rect 18739 7701 18748 7735
rect 18696 7692 18748 7701
rect 20720 7735 20772 7744
rect 20720 7701 20729 7735
rect 20729 7701 20763 7735
rect 20763 7701 20772 7735
rect 20720 7692 20772 7701
rect 20812 7735 20864 7744
rect 20812 7701 20821 7735
rect 20821 7701 20855 7735
rect 20855 7701 20864 7735
rect 20812 7692 20864 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 5632 7488 5684 7540
rect 13452 7488 13504 7540
rect 13636 7531 13688 7540
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 15292 7488 15344 7540
rect 16028 7488 16080 7540
rect 17132 7488 17184 7540
rect 18236 7488 18288 7540
rect 19064 7531 19116 7540
rect 19064 7497 19073 7531
rect 19073 7497 19107 7531
rect 19107 7497 19116 7531
rect 19064 7488 19116 7497
rect 20076 7531 20128 7540
rect 20076 7497 20085 7531
rect 20085 7497 20119 7531
rect 20119 7497 20128 7531
rect 20076 7488 20128 7497
rect 20812 7488 20864 7540
rect 21088 7531 21140 7540
rect 21088 7497 21097 7531
rect 21097 7497 21131 7531
rect 21131 7497 21140 7531
rect 21088 7488 21140 7497
rect 14556 7420 14608 7472
rect 10968 7148 11020 7200
rect 15660 7395 15712 7404
rect 15660 7361 15669 7395
rect 15669 7361 15703 7395
rect 15703 7361 15712 7395
rect 15660 7352 15712 7361
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 15568 7327 15620 7336
rect 15568 7293 15577 7327
rect 15577 7293 15611 7327
rect 15611 7293 15620 7327
rect 15568 7284 15620 7293
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 16948 7420 17000 7472
rect 18144 7352 18196 7404
rect 20536 7420 20588 7472
rect 18880 7352 18932 7404
rect 20996 7395 21048 7404
rect 20996 7361 21005 7395
rect 21005 7361 21039 7395
rect 21039 7361 21048 7395
rect 20996 7352 21048 7361
rect 18604 7327 18656 7336
rect 18604 7293 18613 7327
rect 18613 7293 18647 7327
rect 18647 7293 18656 7327
rect 18604 7284 18656 7293
rect 19524 7327 19576 7336
rect 19524 7293 19533 7327
rect 19533 7293 19567 7327
rect 19567 7293 19576 7327
rect 19524 7284 19576 7293
rect 17316 7216 17368 7268
rect 21548 7284 21600 7336
rect 19708 7216 19760 7268
rect 17408 7148 17460 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 13452 6944 13504 6996
rect 20076 6944 20128 6996
rect 20720 6944 20772 6996
rect 15292 6808 15344 6860
rect 15660 6808 15712 6860
rect 16396 6808 16448 6860
rect 16672 6740 16724 6792
rect 17408 6808 17460 6860
rect 17868 6876 17920 6928
rect 17960 6808 18012 6860
rect 18052 6808 18104 6860
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 18788 6876 18840 6928
rect 21180 6876 21232 6928
rect 20720 6808 20772 6860
rect 21548 6808 21600 6860
rect 21640 6740 21692 6792
rect 13360 6604 13412 6656
rect 15660 6604 15712 6656
rect 16120 6604 16172 6656
rect 16304 6604 16356 6656
rect 17408 6604 17460 6656
rect 18512 6672 18564 6724
rect 17868 6604 17920 6656
rect 22192 6672 22244 6724
rect 19524 6647 19576 6656
rect 19524 6613 19533 6647
rect 19533 6613 19567 6647
rect 19567 6613 19576 6647
rect 19524 6604 19576 6613
rect 19616 6647 19668 6656
rect 19616 6613 19625 6647
rect 19625 6613 19659 6647
rect 19659 6613 19668 6647
rect 19616 6604 19668 6613
rect 20168 6604 20220 6656
rect 21548 6604 21600 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 15936 6400 15988 6452
rect 16304 6443 16356 6452
rect 16304 6409 16313 6443
rect 16313 6409 16347 6443
rect 16347 6409 16356 6443
rect 16304 6400 16356 6409
rect 17408 6443 17460 6452
rect 17408 6409 17417 6443
rect 17417 6409 17451 6443
rect 17451 6409 17460 6443
rect 17408 6400 17460 6409
rect 18604 6400 18656 6452
rect 19616 6400 19668 6452
rect 21088 6400 21140 6452
rect 9772 6060 9824 6112
rect 16396 6332 16448 6384
rect 15200 6264 15252 6316
rect 16028 6264 16080 6316
rect 19432 6332 19484 6384
rect 12900 6196 12952 6248
rect 16304 6196 16356 6248
rect 17408 6196 17460 6248
rect 15936 6060 15988 6112
rect 17868 6264 17920 6316
rect 18052 6307 18104 6316
rect 18052 6273 18061 6307
rect 18061 6273 18095 6307
rect 18095 6273 18104 6307
rect 18052 6264 18104 6273
rect 20536 6264 20588 6316
rect 20996 6264 21048 6316
rect 21364 6264 21416 6316
rect 17960 6239 18012 6248
rect 17960 6205 17969 6239
rect 17969 6205 18003 6239
rect 18003 6205 18012 6239
rect 17960 6196 18012 6205
rect 18972 6196 19024 6248
rect 21180 6239 21232 6248
rect 21180 6205 21189 6239
rect 21189 6205 21223 6239
rect 21223 6205 21232 6239
rect 21180 6196 21232 6205
rect 22468 6196 22520 6248
rect 19708 6128 19760 6180
rect 18328 6060 18380 6112
rect 18788 6103 18840 6112
rect 18788 6069 18797 6103
rect 18797 6069 18831 6103
rect 18831 6069 18840 6103
rect 18788 6060 18840 6069
rect 19432 6060 19484 6112
rect 19616 6060 19668 6112
rect 20076 6060 20128 6112
rect 20812 6060 20864 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 16948 5856 17000 5908
rect 17868 5856 17920 5908
rect 18880 5899 18932 5908
rect 18880 5865 18889 5899
rect 18889 5865 18923 5899
rect 18923 5865 18932 5899
rect 18880 5856 18932 5865
rect 19524 5899 19576 5908
rect 19524 5865 19533 5899
rect 19533 5865 19567 5899
rect 19567 5865 19576 5899
rect 19524 5856 19576 5865
rect 20536 5899 20588 5908
rect 20536 5865 20545 5899
rect 20545 5865 20579 5899
rect 20579 5865 20588 5899
rect 20536 5856 20588 5865
rect 19892 5788 19944 5840
rect 17224 5763 17276 5772
rect 17224 5729 17233 5763
rect 17233 5729 17267 5763
rect 17267 5729 17276 5763
rect 17224 5720 17276 5729
rect 18972 5720 19024 5772
rect 20720 5720 20772 5772
rect 21180 5763 21232 5772
rect 21180 5729 21189 5763
rect 21189 5729 21223 5763
rect 21223 5729 21232 5763
rect 21180 5720 21232 5729
rect 14740 5652 14792 5704
rect 16028 5652 16080 5704
rect 18880 5652 18932 5704
rect 13452 5584 13504 5636
rect 17132 5584 17184 5636
rect 18696 5584 18748 5636
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 15936 5516 15988 5568
rect 17776 5516 17828 5568
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 18512 5559 18564 5568
rect 18512 5525 18521 5559
rect 18521 5525 18555 5559
rect 18555 5525 18564 5559
rect 18512 5516 18564 5525
rect 19616 5516 19668 5568
rect 21640 5584 21692 5636
rect 20720 5516 20772 5568
rect 20996 5559 21048 5568
rect 20996 5525 21005 5559
rect 21005 5525 21039 5559
rect 21039 5525 21048 5559
rect 20996 5516 21048 5525
rect 21548 5516 21600 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 15660 5312 15712 5364
rect 16304 5355 16356 5364
rect 16304 5321 16313 5355
rect 16313 5321 16347 5355
rect 16347 5321 16356 5355
rect 16304 5312 16356 5321
rect 17684 5312 17736 5364
rect 17960 5312 18012 5364
rect 18512 5312 18564 5364
rect 19432 5312 19484 5364
rect 20996 5355 21048 5364
rect 20996 5321 21005 5355
rect 21005 5321 21039 5355
rect 21039 5321 21048 5355
rect 20996 5312 21048 5321
rect 18880 5244 18932 5296
rect 17040 5176 17092 5228
rect 21272 5176 21324 5228
rect 16028 5108 16080 5160
rect 17684 5151 17736 5160
rect 17684 5117 17693 5151
rect 17693 5117 17727 5151
rect 17727 5117 17736 5151
rect 17684 5108 17736 5117
rect 17776 5151 17828 5160
rect 17776 5117 17785 5151
rect 17785 5117 17819 5151
rect 17819 5117 17828 5151
rect 17776 5108 17828 5117
rect 18696 5040 18748 5092
rect 18972 4972 19024 5024
rect 19708 4972 19760 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 18052 4768 18104 4820
rect 18236 4768 18288 4820
rect 19708 4768 19760 4820
rect 21180 4768 21232 4820
rect 14924 4700 14976 4752
rect 14648 4632 14700 4684
rect 15936 4632 15988 4684
rect 17684 4632 17736 4684
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 18052 4564 18104 4616
rect 20536 4564 20588 4616
rect 12348 4428 12400 4480
rect 17316 4496 17368 4548
rect 18328 4496 18380 4548
rect 17040 4428 17092 4480
rect 17408 4428 17460 4480
rect 18972 4428 19024 4480
rect 19616 4471 19668 4480
rect 19616 4437 19625 4471
rect 19625 4437 19659 4471
rect 19659 4437 19668 4471
rect 19616 4428 19668 4437
rect 20168 4428 20220 4480
rect 21364 4471 21416 4480
rect 21364 4437 21373 4471
rect 21373 4437 21407 4471
rect 21407 4437 21416 4471
rect 21364 4428 21416 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 15936 4267 15988 4276
rect 15936 4233 15945 4267
rect 15945 4233 15979 4267
rect 15979 4233 15988 4267
rect 15936 4224 15988 4233
rect 17408 4156 17460 4208
rect 19064 4156 19116 4208
rect 10324 4088 10376 4140
rect 15200 4088 15252 4140
rect 15384 4088 15436 4140
rect 10784 4020 10836 4072
rect 17408 4063 17460 4072
rect 17408 4029 17417 4063
rect 17417 4029 17451 4063
rect 17451 4029 17460 4063
rect 17408 4020 17460 4029
rect 17960 4063 18012 4072
rect 17960 4029 17969 4063
rect 17969 4029 18003 4063
rect 18003 4029 18012 4063
rect 17960 4020 18012 4029
rect 18696 4020 18748 4072
rect 19340 4088 19392 4140
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 2504 3952 2556 4004
rect 9220 3952 9272 4004
rect 15936 3952 15988 4004
rect 16948 3884 17000 3936
rect 17132 3927 17184 3936
rect 17132 3893 17141 3927
rect 17141 3893 17175 3927
rect 17175 3893 17184 3927
rect 17132 3884 17184 3893
rect 18420 3952 18472 4004
rect 20444 4020 20496 4072
rect 20904 4020 20956 4072
rect 20536 3952 20588 4004
rect 21456 4088 21508 4140
rect 18972 3884 19024 3936
rect 19524 3884 19576 3936
rect 19800 3927 19852 3936
rect 19800 3893 19809 3927
rect 19809 3893 19843 3927
rect 19843 3893 19852 3927
rect 19800 3884 19852 3893
rect 19892 3884 19944 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 3884 3680 3936 3732
rect 10968 3680 11020 3732
rect 16948 3680 17000 3732
rect 21180 3723 21232 3732
rect 21180 3689 21189 3723
rect 21189 3689 21223 3723
rect 21223 3689 21232 3723
rect 21180 3680 21232 3689
rect 4804 3612 4856 3664
rect 12348 3612 12400 3664
rect 18144 3612 18196 3664
rect 18604 3612 18656 3664
rect 8484 3544 8536 3596
rect 17040 3544 17092 3596
rect 18696 3587 18748 3596
rect 18696 3553 18705 3587
rect 18705 3553 18739 3587
rect 18739 3553 18748 3587
rect 18696 3544 18748 3553
rect 20260 3544 20312 3596
rect 2780 3476 2832 3528
rect 3424 3476 3476 3528
rect 9404 3476 9456 3528
rect 15568 3476 15620 3528
rect 16672 3519 16724 3528
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 17132 3476 17184 3528
rect 17316 3519 17368 3528
rect 17316 3485 17325 3519
rect 17325 3485 17359 3519
rect 17359 3485 17368 3519
rect 17316 3476 17368 3485
rect 17408 3476 17460 3528
rect 19340 3476 19392 3528
rect 19524 3519 19576 3528
rect 19524 3485 19533 3519
rect 19533 3485 19567 3519
rect 19567 3485 19576 3519
rect 19524 3476 19576 3485
rect 19616 3476 19668 3528
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 20168 3476 20220 3528
rect 22100 3476 22152 3528
rect 2044 3408 2096 3460
rect 7564 3408 7616 3460
rect 13544 3408 13596 3460
rect 16304 3408 16356 3460
rect 19800 3408 19852 3460
rect 9772 3340 9824 3392
rect 9864 3340 9916 3392
rect 15108 3340 15160 3392
rect 17224 3340 17276 3392
rect 17960 3340 18012 3392
rect 18328 3383 18380 3392
rect 18328 3349 18337 3383
rect 18337 3349 18371 3383
rect 18371 3349 18380 3383
rect 18328 3340 18380 3349
rect 19340 3340 19392 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 8024 3136 8076 3188
rect 13728 3136 13780 3188
rect 14280 3136 14332 3188
rect 17040 3136 17092 3188
rect 17408 3136 17460 3188
rect 18052 3179 18104 3188
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 18144 3136 18196 3188
rect 12164 3068 12216 3120
rect 19156 3068 19208 3120
rect 19432 3068 19484 3120
rect 12900 3043 12952 3052
rect 12900 3009 12909 3043
rect 12909 3009 12943 3043
rect 12943 3009 12952 3043
rect 12900 3000 12952 3009
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 16028 3043 16080 3052
rect 16028 3009 16037 3043
rect 16037 3009 16071 3043
rect 16071 3009 16080 3043
rect 16028 3000 16080 3009
rect 17776 3000 17828 3052
rect 19064 3000 19116 3052
rect 19340 3043 19392 3052
rect 19340 3009 19349 3043
rect 19349 3009 19383 3043
rect 19383 3009 19392 3043
rect 19340 3000 19392 3009
rect 19984 3068 20036 3120
rect 14464 2932 14516 2984
rect 16672 2932 16724 2984
rect 20352 3000 20404 3052
rect 20628 3000 20680 3052
rect 20260 2932 20312 2984
rect 11704 2864 11756 2916
rect 13544 2864 13596 2916
rect 17684 2864 17736 2916
rect 19984 2864 20036 2916
rect 12624 2796 12676 2848
rect 13084 2796 13136 2848
rect 15200 2796 15252 2848
rect 18788 2839 18840 2848
rect 18788 2805 18797 2839
rect 18797 2805 18831 2839
rect 18831 2805 18840 2839
rect 18788 2796 18840 2805
rect 19156 2839 19208 2848
rect 19156 2805 19165 2839
rect 19165 2805 19199 2839
rect 19199 2805 19208 2839
rect 19156 2796 19208 2805
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 15200 2592 15252 2644
rect 19708 2592 19760 2644
rect 19064 2524 19116 2576
rect 20260 2456 20312 2508
rect 19616 2388 19668 2440
rect 19800 2431 19852 2440
rect 19800 2397 19809 2431
rect 19809 2397 19843 2431
rect 19843 2397 19852 2431
rect 22376 2456 22428 2508
rect 19800 2388 19852 2397
rect 20996 2388 21048 2440
rect 21088 2431 21140 2440
rect 21088 2397 21097 2431
rect 21097 2397 21131 2431
rect 21131 2397 21140 2431
rect 21088 2388 21140 2397
rect 17960 2252 18012 2304
rect 18236 2252 18288 2304
rect 19340 2252 19392 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 5540 2048 5592 2100
rect 6184 2048 6236 2100
rect 17960 2048 18012 2100
rect 21088 2048 21140 2100
rect 18236 1980 18288 2032
rect 19800 1980 19852 2032
<< metal2 >>
rect 5722 22200 5778 23000
rect 16960 22222 17172 22250
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 5172 19984 5224 19990
rect 5170 19952 5172 19961
rect 5224 19952 5226 19961
rect 5170 19887 5226 19896
rect 4066 19816 4122 19825
rect 4066 19751 4122 19760
rect 4080 19718 4108 19751
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2044 3460 2096 3466
rect 2044 3402 2096 3408
rect 2056 800 2084 3402
rect 2516 800 2544 3946
rect 2792 3534 2820 9862
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2976 800 3004 10202
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3436 800 3464 3470
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3896 800 3924 3674
rect 4356 800 4384 9658
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4816 800 4844 3606
rect 5276 800 5304 8366
rect 5552 2106 5580 12650
rect 5736 7886 5764 22200
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 6550 20496 6606 20505
rect 6550 20431 6606 20440
rect 6564 20058 6592 20431
rect 16212 20392 16264 20398
rect 16212 20334 16264 20340
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 16224 20058 16252 20334
rect 6552 20052 6604 20058
rect 6552 19994 6604 20000
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 5908 19780 5960 19786
rect 5908 19722 5960 19728
rect 5920 19417 5948 19722
rect 9588 19712 9640 19718
rect 9640 19660 9720 19666
rect 9588 19654 9720 19660
rect 9600 19638 9720 19654
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 9692 19514 9720 19638
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 5906 19408 5962 19417
rect 5906 19343 5962 19352
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 9876 16250 9904 19790
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 10060 18834 10088 19314
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 10152 15162 10180 19450
rect 10508 19440 10560 19446
rect 10508 19382 10560 19388
rect 10520 17898 10548 19382
rect 10980 19378 11008 19926
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11256 19514 11284 19654
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10244 17870 10548 17898
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 10244 14618 10272 17870
rect 10612 16046 10640 18022
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11716 17338 11744 19790
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 14372 19440 14424 19446
rect 14372 19382 14424 19388
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 11900 18834 11928 19314
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 11900 16658 11928 17138
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10520 14482 10548 14962
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 7546 5672 7686
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5828 6914 5856 10678
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 5736 6886 5856 6914
rect 5540 2100 5592 2106
rect 5540 2042 5592 2048
rect 5736 800 5764 6886
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6184 2100 6236 2106
rect 6184 2042 6236 2048
rect 6196 800 6224 2042
rect 6656 800 6684 11018
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 800 7144 9318
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7576 800 7604 3402
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8036 800 8064 3130
rect 8496 800 8524 3538
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 9140 2530 9168 8298
rect 9232 4010 9260 14214
rect 11072 12986 11100 14214
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11624 11218 11652 11494
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11992 10198 12020 17070
rect 12360 16658 12388 17138
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12452 16590 12480 19178
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18748 12572 19110
rect 12624 18760 12676 18766
rect 12544 18720 12624 18748
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12256 15020 12308 15026
rect 12256 14962 12308 14968
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12176 11354 12204 12038
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12268 10810 12296 14962
rect 12452 14074 12480 14962
rect 12544 14958 12572 18720
rect 12624 18702 12676 18708
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12820 18086 12848 18634
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12728 14822 12756 16458
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12452 12918 12480 14010
rect 12440 12912 12492 12918
rect 12440 12854 12492 12860
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12544 11898 12572 12582
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12728 11694 12756 14758
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 12986 12848 13126
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12912 11354 12940 19314
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14188 18760 14240 18766
rect 14292 18748 14320 19246
rect 14240 18720 14320 18748
rect 14188 18702 14240 18708
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13832 18358 13860 18566
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 14200 18290 14228 18702
rect 14384 18578 14412 19382
rect 14292 18550 14412 18578
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13832 16574 13860 17138
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 13832 16546 13952 16574
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 16250 13860 16390
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 14006 13032 14350
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 13004 12850 13032 13942
rect 13280 12850 13308 14214
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12360 10742 12388 11018
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12348 10736 12400 10742
rect 12348 10678 12400 10684
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 12452 10062 12480 10610
rect 12728 10606 12756 10950
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 10266 12756 10542
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 12820 9450 12848 11086
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 8956 2502 9168 2530
rect 8956 800 8984 2502
rect 9416 800 9444 3470
rect 9784 3398 9812 6054
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9876 800 9904 3334
rect 10336 800 10364 4082
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10796 800 10824 4014
rect 10980 3738 11008 7142
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11256 800 11284 9114
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 13280 7954 13308 12786
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13372 9654 13400 9862
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 13372 9382 13400 9590
rect 13556 9518 13584 12786
rect 13740 12356 13768 16186
rect 13832 16114 13860 16186
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13924 15994 13952 16546
rect 13832 15966 13952 15994
rect 13832 14074 13860 15966
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13832 13530 13860 13738
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13648 12328 13768 12356
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13268 7948 13320 7954
rect 13268 7890 13320 7896
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 13372 6662 13400 9318
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13464 7002 13492 7482
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 12360 3670 12388 4422
rect 12348 3664 12400 3670
rect 12348 3606 12400 3612
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 11704 2916 11756 2922
rect 11704 2858 11756 2864
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11716 800 11744 2858
rect 12176 800 12204 3062
rect 12912 3058 12940 6190
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 13464 3058 13492 5578
rect 13556 3466 13584 7686
rect 13648 7546 13676 12328
rect 13832 12306 13860 13466
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13912 12368 13964 12374
rect 13912 12310 13964 12316
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13924 12186 13952 12310
rect 13832 12158 13952 12186
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13740 10266 13768 10610
rect 13728 10260 13780 10266
rect 13728 10202 13780 10208
rect 13740 9722 13768 10202
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13740 3194 13768 9386
rect 13832 8566 13860 12158
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 14292 10606 14320 18550
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14384 16590 14412 17138
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14384 16114 14412 16526
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14384 15026 14412 16050
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14384 12374 14412 14010
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14476 12186 14504 18294
rect 14568 17270 14596 19654
rect 14936 19446 14964 19654
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 15120 19378 15148 19722
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 14660 17338 14688 19314
rect 15200 18692 15252 18698
rect 15200 18634 15252 18640
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14568 16998 14596 17206
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14384 12158 14504 12186
rect 14280 10600 14332 10606
rect 14280 10542 14332 10548
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 14384 10010 14412 12158
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11898 14504 12038
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14462 11792 14518 11801
rect 14462 11727 14518 11736
rect 14292 9982 14412 10010
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 14292 7342 14320 9982
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14384 8090 14412 9862
rect 14476 8514 14504 11727
rect 14568 11218 14596 12922
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14568 8634 14596 8774
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14476 8486 14596 8514
rect 14568 8430 14596 8486
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14568 7478 14596 8366
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 14660 4690 14688 17274
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14844 13938 14872 14010
rect 14832 13932 14884 13938
rect 14832 13874 14884 13880
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14752 12986 14780 13466
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14844 12866 14872 13874
rect 14752 12838 14872 12866
rect 14752 11801 14780 12838
rect 14738 11792 14794 11801
rect 14738 11727 14794 11736
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14752 11150 14780 11630
rect 14844 11354 14872 11698
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14936 11218 14964 16186
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15120 15366 15148 16050
rect 15212 15994 15240 18634
rect 15304 18630 15332 19722
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 15304 16182 15332 18566
rect 15396 18222 15424 19110
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15396 16522 15424 16934
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15212 15966 15332 15994
rect 15304 15910 15332 15966
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15120 14618 15148 15302
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15212 13410 15240 14282
rect 15120 13382 15240 13410
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14740 11144 14792 11150
rect 14740 11086 14792 11092
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14752 5710 14780 10746
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14844 10266 14872 10610
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 15028 10130 15056 12582
rect 15120 11370 15148 13382
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15212 11558 15240 13194
rect 15304 11694 15332 15846
rect 15396 13818 15424 16458
rect 15568 16176 15620 16182
rect 15568 16118 15620 16124
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15488 14482 15516 14962
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15488 13938 15516 14418
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15396 13790 15516 13818
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15120 11342 15240 11370
rect 15396 11354 15424 11630
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 15212 9654 15240 11342
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15488 11286 15516 13790
rect 15580 12434 15608 16118
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 14346 15700 15846
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15672 13394 15700 13874
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15672 12918 15700 13330
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15580 12406 15700 12434
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15580 11898 15608 12038
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15488 9722 15516 10406
rect 15580 9994 15608 10950
rect 15672 10198 15700 12406
rect 15856 12306 15884 19450
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 16132 15434 16160 16390
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15568 9988 15620 9994
rect 15568 9930 15620 9936
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15488 9518 15516 9658
rect 15476 9512 15528 9518
rect 15476 9454 15528 9460
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15212 6322 15240 8774
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15304 7546 15332 7686
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15580 7342 15608 7686
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15290 6896 15346 6905
rect 15290 6831 15292 6840
rect 15344 6831 15346 6840
rect 15292 6802 15344 6808
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 12636 800 12664 2790
rect 13096 800 13124 2790
rect 13556 800 13584 2858
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14016 870 14136 898
rect 14016 800 14044 870
rect 2042 0 2098 800
rect 2502 0 2558 800
rect 2962 0 3018 800
rect 3422 0 3478 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5262 0 5318 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7562 0 7618 800
rect 8022 0 8078 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10782 0 10838 800
rect 11242 0 11298 800
rect 11702 0 11758 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14108 762 14136 870
rect 14292 762 14320 3130
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14476 800 14504 2926
rect 14936 800 14964 4694
rect 15106 4176 15162 4185
rect 15212 4146 15240 5510
rect 15106 4111 15162 4120
rect 15200 4140 15252 4146
rect 15120 3398 15148 4111
rect 15200 4082 15252 4088
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15212 2650 15240 2790
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15396 800 15424 4082
rect 15580 3534 15608 7278
rect 15672 6866 15700 7346
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15672 5681 15700 6598
rect 15658 5672 15714 5681
rect 15658 5607 15714 5616
rect 15672 5370 15700 5607
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15764 4826 15792 12038
rect 16132 11898 16160 12038
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 11082 15884 11494
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 10266 15976 10610
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16132 8974 16160 10202
rect 16224 9042 16252 19994
rect 16396 19780 16448 19786
rect 16396 19722 16448 19728
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16316 16250 16344 18158
rect 16408 17882 16436 19722
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16960 19378 16988 22222
rect 17144 22114 17172 22222
rect 17222 22200 17278 23000
rect 17236 22114 17264 22200
rect 17144 22086 17264 22114
rect 17958 21448 18014 21457
rect 17958 21383 18014 21392
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16592 18766 16620 19246
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16304 16244 16356 16250
rect 16304 16186 16356 16192
rect 16304 14544 16356 14550
rect 16302 14512 16304 14521
rect 16356 14512 16358 14521
rect 16302 14447 16358 14456
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16316 10130 16344 14350
rect 16408 10606 16436 17818
rect 16960 17610 16988 19314
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16960 14006 16988 16458
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16960 11286 16988 13942
rect 17052 11898 17080 20402
rect 17500 20392 17552 20398
rect 17500 20334 17552 20340
rect 17512 19854 17540 20334
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17972 18986 18000 21383
rect 18878 21040 18934 21049
rect 18878 20975 18934 20984
rect 18892 20534 18920 20975
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 18880 20528 18932 20534
rect 21192 20505 21220 20538
rect 18880 20470 18932 20476
rect 21178 20496 21234 20505
rect 18892 19854 18920 20470
rect 19708 20460 19760 20466
rect 21178 20431 21234 20440
rect 19708 20402 19760 20408
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18064 19446 18092 19790
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 18340 19514 18368 19722
rect 18144 19508 18196 19514
rect 18144 19450 18196 19456
rect 18328 19508 18380 19514
rect 18328 19450 18380 19456
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 18156 19281 18184 19450
rect 18142 19272 18198 19281
rect 18142 19207 18198 19216
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 17972 18958 18092 18986
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17144 14074 17172 18566
rect 17420 18290 17448 18702
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17420 17882 17448 18226
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17512 17678 17540 18566
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16960 10810 16988 10950
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17052 10742 17080 11018
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16592 10198 16620 10678
rect 17144 10674 17172 12038
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 16316 9654 16344 9862
rect 16304 9648 16356 9654
rect 16304 9590 16356 9596
rect 16408 9450 16436 9862
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16396 9444 16448 9450
rect 16396 9386 16448 9392
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 16040 7954 16068 8434
rect 16960 8362 16988 8842
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16776 7886 16804 8230
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15948 6118 15976 6394
rect 16040 6322 16068 7482
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15948 5574 15976 6054
rect 16040 5710 16068 6258
rect 16028 5704 16080 5710
rect 16028 5646 16080 5652
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15948 4690 15976 5510
rect 16028 5160 16080 5166
rect 16028 5102 16080 5108
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15948 4282 15976 4626
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15948 1986 15976 3946
rect 16040 3058 16068 5102
rect 16132 4622 16160 6598
rect 16316 6458 16344 6598
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16408 6390 16436 6802
rect 16684 6798 16712 7278
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16316 5370 16344 6190
rect 16960 5914 16988 7414
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 17052 5234 17080 9862
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17144 7546 17172 8570
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 17236 5778 17264 13194
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17328 8838 17356 13126
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17328 7274 17356 8434
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 17420 7206 17448 11222
rect 17512 11218 17540 17614
rect 17696 17338 17724 18634
rect 17774 17776 17830 17785
rect 17774 17711 17830 17720
rect 17960 17740 18012 17746
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17696 11694 17724 17274
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17604 10810 17632 11630
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 10130 17540 10406
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17512 9178 17540 9318
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17420 6866 17448 7142
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 6458 17448 6598
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17604 6338 17632 10134
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17696 8634 17724 9522
rect 17788 8634 17816 17711
rect 17960 17682 18012 17688
rect 17972 16794 18000 17682
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17972 16114 18000 16730
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17972 15570 18000 16050
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17880 14346 17908 14758
rect 17868 14340 17920 14346
rect 17868 14282 17920 14288
rect 17880 9738 17908 14282
rect 18064 11914 18092 18958
rect 18248 16794 18276 19110
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18420 17604 18472 17610
rect 18420 17546 18472 17552
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18248 16590 18276 16730
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 18156 14074 18184 14282
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18156 12434 18184 14010
rect 18156 12406 18276 12434
rect 18064 11886 18184 11914
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 17972 11218 18000 11698
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17972 10130 18000 10542
rect 18064 10538 18092 11698
rect 18156 11218 18184 11886
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18144 10736 18196 10742
rect 18144 10678 18196 10684
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17880 9710 18092 9738
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 17880 6934 17908 8774
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17868 6928 17920 6934
rect 17868 6870 17920 6876
rect 17880 6746 17908 6870
rect 17972 6866 18000 8366
rect 18064 6866 18092 9710
rect 18156 9382 18184 10678
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18156 8090 18184 8774
rect 18248 8430 18276 12406
rect 18340 10606 18368 17206
rect 18432 10606 18460 17546
rect 18708 16574 18736 18634
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18800 17270 18828 18022
rect 18984 17610 19012 20198
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 18972 17604 19024 17610
rect 18972 17546 19024 17552
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 19076 17202 19104 18702
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19536 17762 19564 20198
rect 19720 19514 19748 20402
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20732 19854 20760 20334
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20260 19780 20312 19786
rect 20260 19722 20312 19728
rect 19708 19508 19760 19514
rect 19708 19450 19760 19456
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19444 17734 19564 17762
rect 19444 17338 19472 17734
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19536 16590 19564 17614
rect 19064 16584 19116 16590
rect 18708 16546 19012 16574
rect 18708 16454 18736 16546
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18786 16144 18842 16153
rect 18786 16079 18842 16088
rect 18510 15600 18566 15609
rect 18510 15535 18566 15544
rect 18524 11898 18552 15535
rect 18694 15464 18750 15473
rect 18694 15399 18750 15408
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18616 13938 18644 14214
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18524 10674 18552 10950
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18340 9654 18368 9930
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18340 7886 18368 8434
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18156 7410 18184 7686
rect 18248 7546 18276 7754
rect 18432 7698 18460 10066
rect 18524 9926 18552 10610
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18340 7670 18460 7698
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18234 7304 18290 7313
rect 18234 7239 18290 7248
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18248 6798 18276 7239
rect 17420 6310 17632 6338
rect 17696 6718 17908 6746
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 17420 6254 17448 6310
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17132 5636 17184 5642
rect 17132 5578 17184 5584
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 17040 4480 17092 4486
rect 17144 4468 17172 5578
rect 17316 4548 17368 4554
rect 17316 4490 17368 4496
rect 17092 4440 17172 4468
rect 17040 4422 17092 4428
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16946 4312 17002 4321
rect 16946 4247 17002 4256
rect 16960 3942 16988 4247
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16672 3528 16724 3534
rect 16670 3496 16672 3505
rect 16724 3496 16726 3505
rect 16304 3460 16356 3466
rect 16670 3431 16726 3440
rect 16304 3402 16356 3408
rect 16028 3052 16080 3058
rect 16028 2994 16080 3000
rect 15856 1958 15976 1986
rect 15856 800 15884 1958
rect 16316 800 16344 3402
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 16670 3088 16726 3097
rect 16670 3023 16726 3032
rect 16684 2990 16712 3023
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16960 1714 16988 3674
rect 17052 3602 17080 4422
rect 17130 4040 17186 4049
rect 17130 3975 17186 3984
rect 17144 3942 17172 3975
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17130 3632 17186 3641
rect 17040 3596 17092 3602
rect 17130 3567 17186 3576
rect 17040 3538 17092 3544
rect 17144 3534 17172 3567
rect 17328 3534 17356 4490
rect 17420 4486 17448 6190
rect 17696 5370 17724 6718
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17880 6322 17908 6598
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17880 5914 17908 6258
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17682 5264 17738 5273
rect 17682 5199 17738 5208
rect 17696 5166 17724 5199
rect 17788 5166 17816 5510
rect 17972 5370 18000 6190
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17696 4690 17724 5102
rect 18064 4826 18092 6258
rect 18248 4826 18276 6734
rect 18340 6118 18368 7670
rect 18524 6730 18552 9862
rect 18616 8362 18644 13874
rect 18708 12442 18736 15399
rect 18696 12436 18748 12442
rect 18696 12378 18748 12384
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 11014 18736 11494
rect 18800 11354 18828 16079
rect 18878 12200 18934 12209
rect 18878 12135 18934 12144
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18892 11286 18920 12135
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18696 11008 18748 11014
rect 18696 10950 18748 10956
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18616 7954 18644 8298
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18708 7750 18736 8230
rect 18800 7818 18828 11154
rect 18892 11082 18920 11222
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18892 8362 18920 9454
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18604 7336 18656 7342
rect 18604 7278 18656 7284
rect 18512 6724 18564 6730
rect 18512 6666 18564 6672
rect 18616 6458 18644 7278
rect 18604 6452 18656 6458
rect 18604 6394 18656 6400
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 17684 4684 17736 4690
rect 17684 4626 17736 4632
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 17408 4480 17460 4486
rect 17408 4422 17460 4428
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17420 4078 17448 4150
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17038 3224 17094 3233
rect 17038 3159 17040 3168
rect 17092 3159 17094 3168
rect 17040 3130 17092 3136
rect 16776 1686 16988 1714
rect 16776 800 16804 1686
rect 17236 800 17264 3334
rect 17420 3194 17448 3470
rect 17972 3398 18000 4014
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 18064 3194 18092 4558
rect 18340 4554 18368 6054
rect 18708 5642 18736 7686
rect 18800 7041 18828 7754
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18786 7032 18842 7041
rect 18786 6967 18842 6976
rect 18800 6934 18828 6967
rect 18788 6928 18840 6934
rect 18788 6870 18840 6876
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18800 5794 18828 6054
rect 18892 5914 18920 7346
rect 18984 6254 19012 16546
rect 19064 16526 19116 16532
rect 19524 16584 19576 16590
rect 19628 16561 19656 18022
rect 19720 16574 19748 19450
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19904 16574 19932 17274
rect 19984 16584 20036 16590
rect 19524 16526 19576 16532
rect 19614 16552 19670 16561
rect 19076 16046 19104 16526
rect 19720 16546 19840 16574
rect 19614 16487 19670 16496
rect 19524 16176 19576 16182
rect 19524 16118 19576 16124
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 19076 15502 19104 15982
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19076 14414 19104 15438
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19076 14006 19104 14350
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19076 13394 19104 13942
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 19076 12850 19104 13330
rect 19536 12986 19564 16118
rect 19628 15502 19656 16487
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19062 11656 19118 11665
rect 19062 11591 19118 11600
rect 19076 8401 19104 11591
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19168 10538 19196 11018
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19260 9450 19288 9998
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19062 8392 19118 8401
rect 19062 8327 19118 8336
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19154 7984 19210 7993
rect 19536 7954 19564 12174
rect 19154 7919 19210 7928
rect 19524 7948 19576 7954
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19076 7546 19104 7822
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19168 7290 19196 7919
rect 19524 7890 19576 7896
rect 19522 7440 19578 7449
rect 19522 7375 19578 7384
rect 19536 7342 19564 7375
rect 19076 7262 19196 7290
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18800 5766 18920 5794
rect 18984 5778 19012 6190
rect 18892 5710 18920 5766
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 18432 4010 18460 5510
rect 18524 5370 18552 5510
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 18708 5098 18736 5578
rect 18892 5302 18920 5646
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 18696 5092 18748 5098
rect 18696 5034 18748 5040
rect 18708 4078 18736 5034
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 18142 3768 18198 3777
rect 18142 3703 18198 3712
rect 18156 3670 18184 3703
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18328 3392 18380 3398
rect 18326 3360 18328 3369
rect 18380 3360 18382 3369
rect 18326 3295 18382 3304
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17788 2961 17816 2994
rect 17774 2952 17830 2961
rect 17684 2916 17736 2922
rect 17774 2887 17830 2896
rect 17684 2858 17736 2864
rect 17696 800 17724 2858
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17972 2106 18000 2246
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 18156 800 18184 3130
rect 18236 2304 18288 2310
rect 18236 2246 18288 2252
rect 18248 2038 18276 2246
rect 18236 2032 18288 2038
rect 18236 1974 18288 1980
rect 18616 800 18644 3606
rect 18708 3602 18736 4014
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18788 2848 18840 2854
rect 18788 2790 18840 2796
rect 18800 2553 18828 2790
rect 18892 2774 18920 5238
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 18984 4486 19012 4966
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18984 3942 19012 4422
rect 19076 4214 19104 7262
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19628 6746 19656 15302
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19720 13258 19748 13670
rect 19708 13252 19760 13258
rect 19708 13194 19760 13200
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19720 10266 19748 10406
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19812 8430 19840 16546
rect 19904 16546 19984 16574
rect 19904 15366 19932 16546
rect 19984 16526 20036 16532
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19982 13288 20038 13297
rect 19982 13223 20038 13232
rect 20076 13252 20128 13258
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19904 9518 19932 12922
rect 19996 12442 20024 13223
rect 20076 13194 20128 13200
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19800 8424 19852 8430
rect 19706 8392 19762 8401
rect 19800 8366 19852 8372
rect 19706 8327 19762 8336
rect 19720 7426 19748 8327
rect 19720 7398 19840 7426
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 19444 6718 19656 6746
rect 19444 6390 19472 6718
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19444 6118 19472 6326
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19536 5914 19564 6598
rect 19628 6458 19656 6598
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19720 6186 19748 7210
rect 19708 6180 19760 6186
rect 19708 6122 19760 6128
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19628 5794 19656 6054
rect 19444 5766 19656 5794
rect 19444 5370 19472 5766
rect 19812 5658 19840 7398
rect 19904 5846 19932 9318
rect 20088 9110 20116 13194
rect 20166 11248 20222 11257
rect 20166 11183 20222 11192
rect 20180 10810 20208 11183
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20180 10266 20208 10746
rect 20272 10606 20300 19722
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 18737 20668 19654
rect 20732 19446 20760 19790
rect 20916 19553 20944 19790
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 20902 19544 20958 19553
rect 21742 19547 22050 19556
rect 20902 19479 20958 19488
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 20626 18728 20682 18737
rect 20626 18663 20682 18672
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20456 18290 20484 18566
rect 20732 18290 20760 19382
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20720 18284 20772 18290
rect 20720 18226 20772 18232
rect 20456 18193 20484 18226
rect 20442 18184 20498 18193
rect 20442 18119 20498 18128
rect 20732 17678 20760 18226
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20732 17270 20760 17614
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 21100 16998 21128 19314
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21364 17536 21416 17542
rect 21364 17478 21416 17484
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 20916 16574 20944 16934
rect 20534 16552 20590 16561
rect 20916 16546 21036 16574
rect 20534 16487 20590 16496
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20456 14074 20484 16050
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20456 12322 20484 14010
rect 20548 12442 20576 16487
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20626 12880 20682 12889
rect 20626 12815 20682 12824
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20456 12294 20576 12322
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20364 10742 20392 11018
rect 20352 10736 20404 10742
rect 20352 10678 20404 10684
rect 20260 10600 20312 10606
rect 20260 10542 20312 10548
rect 20364 10441 20392 10678
rect 20350 10432 20406 10441
rect 20350 10367 20406 10376
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20456 10130 20484 12174
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 20444 9580 20496 9586
rect 20444 9522 20496 9528
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 20350 8936 20406 8945
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19996 8090 20024 8366
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 20088 7546 20116 8910
rect 20350 8871 20406 8880
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 19982 6760 20038 6769
rect 19982 6695 20038 6704
rect 19892 5840 19944 5846
rect 19892 5782 19944 5788
rect 19536 5630 19840 5658
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19536 4706 19564 5630
rect 19616 5568 19668 5574
rect 19616 5510 19668 5516
rect 19352 4678 19564 4706
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 19076 3058 19104 4150
rect 19352 4146 19380 4678
rect 19628 4486 19656 5510
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19720 4826 19748 4966
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19628 4185 19656 4422
rect 19614 4176 19670 4185
rect 19340 4140 19392 4146
rect 19614 4111 19670 4120
rect 19340 4082 19392 4088
rect 19352 4049 19380 4082
rect 19338 4040 19394 4049
rect 19338 3975 19394 3984
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19536 3777 19564 3878
rect 19522 3768 19578 3777
rect 19522 3703 19578 3712
rect 19340 3528 19392 3534
rect 19524 3528 19576 3534
rect 19392 3476 19472 3482
rect 19340 3470 19472 3476
rect 19524 3470 19576 3476
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19352 3454 19472 3470
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19352 3233 19380 3334
rect 19338 3224 19394 3233
rect 19338 3159 19394 3168
rect 19444 3126 19472 3454
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 19432 3120 19484 3126
rect 19432 3062 19484 3068
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19168 2854 19196 3062
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19352 2961 19380 2994
rect 19338 2952 19394 2961
rect 19338 2887 19394 2896
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 18892 2746 19012 2774
rect 18786 2544 18842 2553
rect 18786 2479 18842 2488
rect 18984 2417 19012 2746
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19064 2576 19116 2582
rect 19536 2530 19564 3470
rect 19064 2518 19116 2524
rect 18970 2408 19026 2417
rect 18970 2343 19026 2352
rect 19076 800 19104 2518
rect 19444 2502 19564 2530
rect 19444 2394 19472 2502
rect 19628 2446 19656 3470
rect 19720 2774 19748 4762
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19812 3466 19840 3878
rect 19800 3460 19852 3466
rect 19800 3402 19852 3408
rect 19904 3097 19932 3878
rect 19996 3126 20024 6695
rect 20088 6118 20116 6938
rect 20180 6662 20208 8434
rect 20258 7440 20314 7449
rect 20258 7375 20314 7384
rect 20168 6656 20220 6662
rect 20168 6598 20220 6604
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 20074 5944 20130 5953
rect 20074 5879 20130 5888
rect 20088 3534 20116 5879
rect 20168 4480 20220 4486
rect 20168 4422 20220 4428
rect 20180 3913 20208 4422
rect 20166 3904 20222 3913
rect 20166 3839 20222 3848
rect 20272 3602 20300 7375
rect 20364 6474 20392 8871
rect 20456 8634 20484 9522
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20548 7478 20576 12294
rect 20640 11898 20668 12815
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20732 11778 20760 14962
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20824 14414 20852 14894
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20640 11750 20760 11778
rect 20812 11756 20864 11762
rect 20640 10198 20668 11750
rect 20812 11698 20864 11704
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20732 10674 20760 11630
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20628 10192 20680 10198
rect 20628 10134 20680 10140
rect 20626 9208 20682 9217
rect 20626 9143 20682 9152
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20364 6446 20484 6474
rect 20350 6352 20406 6361
rect 20350 6287 20406 6296
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20076 3528 20128 3534
rect 20168 3528 20220 3534
rect 20076 3470 20128 3476
rect 20166 3496 20168 3505
rect 20220 3496 20222 3505
rect 20166 3431 20222 3440
rect 19984 3120 20036 3126
rect 19890 3088 19946 3097
rect 19984 3062 20036 3068
rect 20364 3058 20392 6287
rect 20456 4468 20484 6446
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20548 5914 20576 6258
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 20640 4842 20668 9143
rect 20824 9042 20852 11698
rect 20916 9654 20944 13262
rect 21008 11234 21036 16546
rect 21192 15910 21220 17138
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21178 14512 21234 14521
rect 21178 14447 21234 14456
rect 21086 13696 21142 13705
rect 21086 13631 21142 13640
rect 21100 13530 21128 13631
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21100 12918 21128 13126
rect 21088 12912 21140 12918
rect 21088 12854 21140 12860
rect 21192 11354 21220 14447
rect 21284 13938 21312 15302
rect 21376 15026 21404 17478
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21638 17232 21694 17241
rect 21638 17167 21694 17176
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21454 14920 21510 14929
rect 21454 14855 21510 14864
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21284 12306 21312 13874
rect 21376 13870 21404 14350
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21376 12850 21404 13806
rect 21364 12844 21416 12850
rect 21364 12786 21416 12792
rect 21362 12472 21418 12481
rect 21468 12442 21496 14855
rect 21362 12407 21418 12416
rect 21456 12436 21508 12442
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21008 11206 21220 11234
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 20904 9648 20956 9654
rect 20904 9590 20956 9596
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 21008 8906 21036 11086
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20732 7002 20760 7686
rect 20824 7546 20852 7686
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20732 5778 20760 6802
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 20548 4814 20668 4842
rect 20548 4622 20576 4814
rect 20626 4720 20682 4729
rect 20626 4655 20682 4664
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20456 4440 20576 4468
rect 20548 4321 20576 4440
rect 20534 4312 20590 4321
rect 20534 4247 20590 4256
rect 20548 4146 20576 4247
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 19890 3023 19946 3032
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 19720 2746 19932 2774
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 19352 2366 19472 2394
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19352 2310 19380 2366
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19720 1170 19748 2586
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 19812 2038 19840 2382
rect 19800 2032 19852 2038
rect 19800 1974 19852 1980
rect 19904 1465 19932 2746
rect 19890 1456 19946 1465
rect 19890 1391 19946 1400
rect 19536 1142 19748 1170
rect 19536 800 19564 1142
rect 19996 800 20024 2858
rect 20272 2514 20300 2926
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 20456 800 20484 4014
rect 20536 4004 20588 4010
rect 20536 3946 20588 3952
rect 20548 3641 20576 3946
rect 20534 3632 20590 3641
rect 20534 3567 20590 3576
rect 20640 3058 20668 4655
rect 20732 4185 20760 5510
rect 20718 4176 20774 4185
rect 20718 4111 20774 4120
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20824 2774 20852 6054
rect 20916 4078 20944 8774
rect 21100 8498 21128 11018
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 21008 7410 21036 8230
rect 21192 7954 21220 11206
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21100 7546 21128 7754
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 21008 6322 21036 7346
rect 21100 6458 21128 7482
rect 21192 6934 21220 7890
rect 21180 6928 21232 6934
rect 21180 6870 21232 6876
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 20996 6316 21048 6322
rect 20996 6258 21048 6264
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 21192 5778 21220 6190
rect 21180 5772 21232 5778
rect 21180 5714 21232 5720
rect 20994 5672 21050 5681
rect 20994 5607 21050 5616
rect 21008 5574 21036 5607
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 20994 5400 21050 5409
rect 20994 5335 20996 5344
rect 21048 5335 21050 5344
rect 20996 5306 21048 5312
rect 20994 5264 21050 5273
rect 20994 5199 21050 5208
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 20824 2746 20944 2774
rect 20916 800 20944 2746
rect 21008 2446 21036 5199
rect 21086 5128 21142 5137
rect 21086 5063 21142 5072
rect 21100 2446 21128 5063
rect 21192 4826 21220 5714
rect 21284 5234 21312 12106
rect 21376 9654 21404 12407
rect 21456 12378 21508 12384
rect 21456 11620 21508 11626
rect 21456 11562 21508 11568
rect 21468 11082 21496 11562
rect 21456 11076 21508 11082
rect 21456 11018 21508 11024
rect 21364 9648 21416 9654
rect 21364 9590 21416 9596
rect 21454 9616 21510 9625
rect 21376 8974 21404 9590
rect 21454 9551 21510 9560
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21192 3738 21220 4762
rect 21376 4486 21404 6258
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21180 3732 21232 3738
rect 21180 3674 21232 3680
rect 21192 3369 21220 3674
rect 21178 3360 21234 3369
rect 21178 3295 21234 3304
rect 21376 2553 21404 4422
rect 21468 4146 21496 9551
rect 21560 7342 21588 15846
rect 21652 8634 21680 17167
rect 22006 16960 22062 16969
rect 22006 16895 22062 16904
rect 22020 16574 22048 16895
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22020 16546 22140 16574
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 22006 13968 22062 13977
rect 22006 13903 22062 13912
rect 22020 13870 22048 13903
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 22112 10810 22140 16546
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22006 10704 22062 10713
rect 22006 10639 22062 10648
rect 22020 10130 22048 10639
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22006 10024 22062 10033
rect 22062 9982 22140 10010
rect 22006 9959 22062 9968
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21640 8628 21692 8634
rect 21640 8570 21692 8576
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21560 6866 21588 7278
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21560 5574 21588 6598
rect 21652 5642 21680 6734
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21640 5636 21692 5642
rect 21640 5578 21692 5584
rect 21548 5568 21600 5574
rect 21548 5510 21600 5516
rect 21456 4140 21508 4146
rect 21456 4082 21508 4088
rect 21560 2689 21588 5510
rect 21652 3505 21680 5578
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 22112 3534 22140 9982
rect 22204 6730 22232 12242
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 22192 6724 22244 6730
rect 22192 6666 22244 6672
rect 22100 3528 22152 3534
rect 21638 3496 21694 3505
rect 22100 3470 22152 3476
rect 21638 3431 21694 3440
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 21546 2680 21602 2689
rect 21546 2615 21602 2624
rect 21362 2544 21418 2553
rect 22388 2514 22416 10066
rect 22480 6254 22508 16730
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22572 10266 22600 13806
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22468 6248 22520 6254
rect 22468 6190 22520 6196
rect 21362 2479 21418 2488
rect 22376 2508 22428 2514
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 21100 2106 21128 2382
rect 21088 2100 21140 2106
rect 21088 2042 21140 2048
rect 21376 1873 21404 2479
rect 22376 2450 22428 2456
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 21362 1864 21418 1873
rect 21362 1799 21418 1808
rect 14108 734 14320 762
rect 14462 0 14518 800
rect 14922 0 14978 800
rect 15382 0 15438 800
rect 15842 0 15898 800
rect 16302 0 16358 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20442 0 20498 800
rect 20902 0 20958 800
<< via2 >>
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 5170 19932 5172 19952
rect 5172 19932 5224 19952
rect 5224 19932 5226 19952
rect 5170 19896 5226 19932
rect 4066 19760 4122 19816
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 6550 20440 6606 20496
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 5906 19352 5962 19408
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 14462 11736 14518 11792
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 14738 11736 14794 11792
rect 15290 6860 15346 6896
rect 15290 6840 15292 6860
rect 15292 6840 15344 6860
rect 15344 6840 15346 6860
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 15106 4120 15162 4176
rect 15658 5616 15714 5672
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 17958 21392 18014 21448
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16302 14492 16304 14512
rect 16304 14492 16356 14512
rect 16356 14492 16358 14512
rect 16302 14456 16358 14492
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 18878 20984 18934 21040
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21178 20440 21234 20496
rect 18142 19216 18198 19272
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 17774 17720 17830 17776
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 18786 16088 18842 16144
rect 18510 15544 18566 15600
rect 18694 15408 18750 15464
rect 18234 7248 18290 7304
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16946 4256 17002 4312
rect 16670 3476 16672 3496
rect 16672 3476 16724 3496
rect 16724 3476 16726 3496
rect 16670 3440 16726 3476
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 16670 3032 16726 3088
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 17130 3984 17186 4040
rect 17130 3576 17186 3632
rect 17682 5208 17738 5264
rect 18878 12144 18934 12200
rect 17038 3188 17094 3224
rect 17038 3168 17040 3188
rect 17040 3168 17092 3188
rect 17092 3168 17094 3188
rect 18786 6976 18842 7032
rect 19614 16496 19670 16552
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19062 11600 19118 11656
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19062 8336 19118 8392
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19154 7928 19210 7984
rect 19522 7384 19578 7440
rect 18142 3712 18198 3768
rect 18326 3340 18328 3360
rect 18328 3340 18380 3360
rect 18380 3340 18382 3360
rect 18326 3304 18382 3340
rect 17774 2896 17830 2952
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19982 13232 20038 13288
rect 19706 8336 19762 8392
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 20166 11192 20222 11248
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 20902 19488 20958 19544
rect 20626 18672 20682 18728
rect 20442 18128 20498 18184
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 20534 16496 20590 16552
rect 20626 12824 20682 12880
rect 20350 10376 20406 10432
rect 20350 8880 20406 8936
rect 19982 6704 20038 6760
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19614 4120 19670 4176
rect 19338 3984 19394 4040
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19522 3712 19578 3768
rect 19338 3168 19394 3224
rect 19338 2896 19394 2952
rect 18786 2488 18842 2544
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 18970 2352 19026 2408
rect 20258 7384 20314 7440
rect 20074 5888 20130 5944
rect 20166 3848 20222 3904
rect 20626 9152 20682 9208
rect 20350 6296 20406 6352
rect 20166 3476 20168 3496
rect 20168 3476 20220 3496
rect 20220 3476 20222 3496
rect 20166 3440 20222 3476
rect 19890 3032 19946 3088
rect 21178 14456 21234 14512
rect 21086 13640 21142 13696
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21638 17176 21694 17232
rect 21454 14864 21510 14920
rect 21362 12416 21418 12472
rect 20626 4664 20682 4720
rect 20534 4256 20590 4312
rect 19890 1400 19946 1456
rect 20534 3576 20590 3632
rect 20718 4120 20774 4176
rect 20994 5616 21050 5672
rect 20994 5364 21050 5400
rect 20994 5344 20996 5364
rect 20996 5344 21048 5364
rect 21048 5344 21050 5364
rect 20994 5208 21050 5264
rect 21086 5072 21142 5128
rect 21454 9560 21510 9616
rect 21178 3304 21234 3360
rect 22006 16904 22062 16960
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 22006 13912 22062 13968
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 22006 10648 22062 10704
rect 22006 9968 22062 10024
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21638 3440 21694 3496
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21546 2624 21602 2680
rect 21362 2488 21418 2544
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
rect 21362 1808 21418 1864
<< metal3 >>
rect 17953 21450 18019 21453
rect 22200 21450 23000 21480
rect 17953 21448 23000 21450
rect 17953 21392 17958 21448
rect 18014 21392 23000 21448
rect 17953 21390 23000 21392
rect 17953 21387 18019 21390
rect 22200 21360 23000 21390
rect 18873 21042 18939 21045
rect 22200 21042 23000 21072
rect 18873 21040 23000 21042
rect 18873 20984 18878 21040
rect 18934 20984 23000 21040
rect 18873 20982 23000 20984
rect 18873 20979 18939 20982
rect 22200 20952 23000 20982
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 22200 20634 23000 20664
rect 22142 20544 23000 20634
rect 6545 20498 6611 20501
rect 21173 20498 21239 20501
rect 22142 20498 22202 20544
rect 6545 20496 19626 20498
rect 6545 20440 6550 20496
rect 6606 20440 19626 20496
rect 6545 20438 19626 20440
rect 6545 20435 6611 20438
rect 19566 20226 19626 20438
rect 21173 20496 22202 20498
rect 21173 20440 21178 20496
rect 21234 20440 22202 20496
rect 21173 20438 22202 20440
rect 21173 20435 21239 20438
rect 22200 20226 23000 20256
rect 19566 20166 23000 20226
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 22200 20136 23000 20166
rect 19139 20095 19455 20096
rect 5165 19954 5231 19957
rect 5165 19952 19442 19954
rect 5165 19896 5170 19952
rect 5226 19896 19442 19952
rect 5165 19894 19442 19896
rect 5165 19891 5231 19894
rect 4061 19818 4127 19821
rect 19382 19818 19442 19894
rect 22200 19818 23000 19848
rect 4061 19816 19258 19818
rect 4061 19760 4066 19816
rect 4122 19760 19258 19816
rect 4061 19758 19258 19760
rect 19382 19758 23000 19818
rect 4061 19755 4127 19758
rect 19198 19682 19258 19758
rect 22200 19728 23000 19758
rect 19198 19622 21098 19682
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 20897 19546 20963 19549
rect 18646 19544 20963 19546
rect 18646 19488 20902 19544
rect 20958 19488 20963 19544
rect 18646 19486 20963 19488
rect 5901 19410 5967 19413
rect 18646 19410 18706 19486
rect 20897 19483 20963 19486
rect 5901 19408 18706 19410
rect 5901 19352 5906 19408
rect 5962 19352 18706 19408
rect 5901 19350 18706 19352
rect 21038 19410 21098 19622
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 22200 19410 23000 19440
rect 21038 19350 23000 19410
rect 5901 19347 5967 19350
rect 22200 19320 23000 19350
rect 18137 19274 18203 19277
rect 18137 19272 19626 19274
rect 18137 19216 18142 19272
rect 18198 19216 19626 19272
rect 18137 19214 19626 19216
rect 18137 19211 18203 19214
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 19566 19002 19626 19214
rect 22200 19002 23000 19032
rect 19566 18942 23000 19002
rect 22200 18912 23000 18942
rect 20621 18730 20687 18733
rect 20621 18728 22202 18730
rect 20621 18672 20626 18728
rect 20682 18672 22202 18728
rect 20621 18670 22202 18672
rect 20621 18667 20687 18670
rect 22142 18624 22202 18670
rect 22142 18534 23000 18624
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 22200 18504 23000 18534
rect 21738 18463 22054 18464
rect 19558 18124 19564 18188
rect 19628 18186 19634 18188
rect 20437 18186 20503 18189
rect 19628 18184 20503 18186
rect 19628 18128 20442 18184
rect 20498 18128 20503 18184
rect 19628 18126 20503 18128
rect 19628 18124 19634 18126
rect 20437 18123 20503 18126
rect 20662 18124 20668 18188
rect 20732 18186 20738 18188
rect 22200 18186 23000 18216
rect 20732 18126 23000 18186
rect 20732 18124 20738 18126
rect 22200 18096 23000 18126
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 17769 17778 17835 17781
rect 22200 17778 23000 17808
rect 17769 17776 23000 17778
rect 17769 17720 17774 17776
rect 17830 17720 23000 17776
rect 17769 17718 23000 17720
rect 17769 17715 17835 17718
rect 22200 17688 23000 17718
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 22200 17370 23000 17400
rect 22142 17280 23000 17370
rect 21633 17234 21699 17237
rect 22142 17234 22202 17280
rect 21633 17232 22202 17234
rect 21633 17176 21638 17232
rect 21694 17176 22202 17232
rect 21633 17174 22202 17176
rect 21633 17171 21699 17174
rect 22001 16962 22067 16965
rect 22200 16962 23000 16992
rect 22001 16960 23000 16962
rect 22001 16904 22006 16960
rect 22062 16904 23000 16960
rect 22001 16902 23000 16904
rect 22001 16899 22067 16902
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 22200 16872 23000 16902
rect 19139 16831 19455 16832
rect 17718 16492 17724 16556
rect 17788 16554 17794 16556
rect 19609 16554 19675 16557
rect 17788 16552 19675 16554
rect 17788 16496 19614 16552
rect 19670 16496 19675 16552
rect 17788 16494 19675 16496
rect 17788 16492 17794 16494
rect 19609 16491 19675 16494
rect 20529 16554 20595 16557
rect 22200 16554 23000 16584
rect 20529 16552 23000 16554
rect 20529 16496 20534 16552
rect 20590 16496 23000 16552
rect 20529 16494 23000 16496
rect 20529 16491 20595 16494
rect 22200 16464 23000 16494
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 18781 16146 18847 16149
rect 22200 16146 23000 16176
rect 18781 16144 23000 16146
rect 18781 16088 18786 16144
rect 18842 16088 23000 16144
rect 18781 16086 23000 16088
rect 18781 16083 18847 16086
rect 22200 16056 23000 16086
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 22200 15738 23000 15768
rect 19566 15678 23000 15738
rect 18505 15602 18571 15605
rect 19566 15602 19626 15678
rect 22200 15648 23000 15678
rect 18505 15600 19626 15602
rect 18505 15544 18510 15600
rect 18566 15544 19626 15600
rect 18505 15542 19626 15544
rect 18505 15539 18571 15542
rect 18689 15466 18755 15469
rect 18689 15464 22202 15466
rect 18689 15408 18694 15464
rect 18750 15408 22202 15464
rect 18689 15406 22202 15408
rect 18689 15403 18755 15406
rect 22142 15360 22202 15406
rect 22142 15270 23000 15360
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 22200 15240 23000 15270
rect 21738 15199 22054 15200
rect 21449 14922 21515 14925
rect 22200 14922 23000 14952
rect 21449 14920 23000 14922
rect 21449 14864 21454 14920
rect 21510 14864 23000 14920
rect 21449 14862 23000 14864
rect 21449 14859 21515 14862
rect 22200 14832 23000 14862
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 16297 14516 16363 14517
rect 16246 14514 16252 14516
rect 16206 14454 16252 14514
rect 16316 14512 16363 14516
rect 16358 14456 16363 14512
rect 16246 14452 16252 14454
rect 16316 14452 16363 14456
rect 16297 14451 16363 14452
rect 21173 14514 21239 14517
rect 22200 14514 23000 14544
rect 21173 14512 23000 14514
rect 21173 14456 21178 14512
rect 21234 14456 23000 14512
rect 21173 14454 23000 14456
rect 21173 14451 21239 14454
rect 22200 14424 23000 14454
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 22200 14106 23000 14136
rect 22142 14016 23000 14106
rect 22001 13970 22067 13973
rect 22142 13970 22202 14016
rect 22001 13968 22202 13970
rect 22001 13912 22006 13968
rect 22062 13912 22202 13968
rect 22001 13910 22202 13912
rect 22001 13907 22067 13910
rect 21081 13698 21147 13701
rect 22200 13698 23000 13728
rect 21081 13696 23000 13698
rect 21081 13640 21086 13696
rect 21142 13640 23000 13696
rect 21081 13638 23000 13640
rect 21081 13635 21147 13638
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 22200 13608 23000 13638
rect 19139 13567 19455 13568
rect 19977 13290 20043 13293
rect 22200 13290 23000 13320
rect 19977 13288 23000 13290
rect 19977 13232 19982 13288
rect 20038 13232 23000 13288
rect 19977 13230 23000 13232
rect 19977 13227 20043 13230
rect 22200 13200 23000 13230
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 20621 12882 20687 12885
rect 22200 12882 23000 12912
rect 20621 12880 23000 12882
rect 20621 12824 20626 12880
rect 20682 12824 23000 12880
rect 20621 12822 23000 12824
rect 20621 12819 20687 12822
rect 22200 12792 23000 12822
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 21357 12474 21423 12477
rect 22200 12474 23000 12504
rect 21357 12472 23000 12474
rect 21357 12416 21362 12472
rect 21418 12416 23000 12472
rect 21357 12414 23000 12416
rect 21357 12411 21423 12414
rect 22200 12384 23000 12414
rect 18873 12202 18939 12205
rect 18873 12200 22202 12202
rect 18873 12144 18878 12200
rect 18934 12144 22202 12200
rect 18873 12142 22202 12144
rect 18873 12139 18939 12142
rect 22142 12096 22202 12142
rect 22142 12006 23000 12096
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 22200 11976 23000 12006
rect 21738 11935 22054 11936
rect 14457 11794 14523 11797
rect 14733 11794 14799 11797
rect 14457 11792 14799 11794
rect 14457 11736 14462 11792
rect 14518 11736 14738 11792
rect 14794 11736 14799 11792
rect 14457 11734 14799 11736
rect 14457 11731 14523 11734
rect 14733 11731 14799 11734
rect 19057 11658 19123 11661
rect 22200 11658 23000 11688
rect 19057 11656 23000 11658
rect 19057 11600 19062 11656
rect 19118 11600 23000 11656
rect 19057 11598 23000 11600
rect 19057 11595 19123 11598
rect 22200 11568 23000 11598
rect 0 11522 800 11552
rect 0 11462 3434 11522
rect 0 11432 800 11462
rect 3374 11250 3434 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 15326 11250 15332 11252
rect 3374 11190 15332 11250
rect 15326 11188 15332 11190
rect 15396 11250 15402 11252
rect 16246 11250 16252 11252
rect 15396 11190 16252 11250
rect 15396 11188 15402 11190
rect 16246 11188 16252 11190
rect 16316 11188 16322 11252
rect 20161 11250 20227 11253
rect 22200 11250 23000 11280
rect 20161 11248 23000 11250
rect 20161 11192 20166 11248
rect 20222 11192 23000 11248
rect 20161 11190 23000 11192
rect 20161 11187 20227 11190
rect 22200 11160 23000 11190
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 22200 10842 23000 10872
rect 22142 10752 23000 10842
rect 22001 10706 22067 10709
rect 22142 10706 22202 10752
rect 22001 10704 22202 10706
rect 22001 10648 22006 10704
rect 22062 10648 22202 10704
rect 22001 10646 22202 10648
rect 22001 10643 22067 10646
rect 20345 10434 20411 10437
rect 22200 10434 23000 10464
rect 20345 10432 23000 10434
rect 20345 10376 20350 10432
rect 20406 10376 23000 10432
rect 20345 10374 23000 10376
rect 20345 10371 20411 10374
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 22200 10344 23000 10374
rect 19139 10303 19455 10304
rect 22001 10026 22067 10029
rect 22200 10026 23000 10056
rect 22001 10024 23000 10026
rect 22001 9968 22006 10024
rect 22062 9968 23000 10024
rect 22001 9966 23000 9968
rect 22001 9963 22067 9966
rect 22200 9936 23000 9966
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 21449 9618 21515 9621
rect 22200 9618 23000 9648
rect 21449 9616 23000 9618
rect 21449 9560 21454 9616
rect 21510 9560 23000 9616
rect 21449 9558 23000 9560
rect 21449 9555 21515 9558
rect 22200 9528 23000 9558
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 20621 9210 20687 9213
rect 22200 9210 23000 9240
rect 20621 9208 23000 9210
rect 20621 9152 20626 9208
rect 20682 9152 23000 9208
rect 20621 9150 23000 9152
rect 20621 9147 20687 9150
rect 22200 9120 23000 9150
rect 20345 8938 20411 8941
rect 20345 8936 22202 8938
rect 20345 8880 20350 8936
rect 20406 8880 22202 8936
rect 20345 8878 22202 8880
rect 20345 8875 20411 8878
rect 22142 8832 22202 8878
rect 22142 8742 23000 8832
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 22200 8712 23000 8742
rect 21738 8671 22054 8672
rect 19057 8396 19123 8397
rect 19006 8394 19012 8396
rect 18966 8334 19012 8394
rect 19076 8392 19123 8396
rect 19118 8336 19123 8392
rect 19006 8332 19012 8334
rect 19076 8332 19123 8336
rect 19057 8331 19123 8332
rect 19701 8394 19767 8397
rect 22200 8394 23000 8424
rect 19701 8392 23000 8394
rect 19701 8336 19706 8392
rect 19762 8336 23000 8392
rect 19701 8334 23000 8336
rect 19701 8331 19767 8334
rect 22200 8304 23000 8334
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 19149 7986 19215 7989
rect 22200 7986 23000 8016
rect 19149 7984 23000 7986
rect 19149 7928 19154 7984
rect 19210 7928 23000 7984
rect 19149 7926 23000 7928
rect 19149 7923 19215 7926
rect 22200 7896 23000 7926
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 22200 7578 23000 7608
rect 22142 7488 23000 7578
rect 19517 7444 19583 7445
rect 19517 7442 19564 7444
rect 19472 7440 19564 7442
rect 19472 7384 19522 7440
rect 19472 7382 19564 7384
rect 19517 7380 19564 7382
rect 19628 7380 19634 7444
rect 20253 7442 20319 7445
rect 22142 7442 22202 7488
rect 20253 7440 22202 7442
rect 20253 7384 20258 7440
rect 20314 7384 22202 7440
rect 20253 7382 22202 7384
rect 19517 7379 19583 7380
rect 20253 7379 20319 7382
rect 18229 7306 18295 7309
rect 18229 7304 19626 7306
rect 18229 7248 18234 7304
rect 18290 7248 19626 7304
rect 18229 7246 19626 7248
rect 18229 7243 18295 7246
rect 19566 7170 19626 7246
rect 22200 7170 23000 7200
rect 19566 7110 23000 7170
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 22200 7080 23000 7110
rect 19139 7039 19455 7040
rect 18270 6972 18276 7036
rect 18340 7034 18346 7036
rect 18781 7034 18847 7037
rect 18340 7032 18847 7034
rect 18340 6976 18786 7032
rect 18842 6976 18847 7032
rect 18340 6974 18847 6976
rect 18340 6972 18346 6974
rect 18781 6971 18847 6974
rect 15285 6900 15351 6901
rect 15285 6898 15332 6900
rect 15240 6896 15332 6898
rect 15240 6840 15290 6896
rect 15240 6838 15332 6840
rect 15285 6836 15332 6838
rect 15396 6836 15402 6900
rect 15285 6835 15351 6836
rect 19977 6762 20043 6765
rect 22200 6762 23000 6792
rect 19977 6760 23000 6762
rect 19977 6704 19982 6760
rect 20038 6704 23000 6760
rect 19977 6702 23000 6704
rect 19977 6699 20043 6702
rect 22200 6672 23000 6702
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 20345 6354 20411 6357
rect 22200 6354 23000 6384
rect 20345 6352 23000 6354
rect 20345 6296 20350 6352
rect 20406 6296 23000 6352
rect 20345 6294 23000 6296
rect 20345 6291 20411 6294
rect 22200 6264 23000 6294
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 20069 5946 20135 5949
rect 22200 5946 23000 5976
rect 20069 5944 23000 5946
rect 20069 5888 20074 5944
rect 20130 5888 23000 5944
rect 20069 5886 23000 5888
rect 20069 5883 20135 5886
rect 22200 5856 23000 5886
rect 15653 5674 15719 5677
rect 20989 5674 21055 5677
rect 15653 5672 21055 5674
rect 15653 5616 15658 5672
rect 15714 5616 20994 5672
rect 21050 5616 21055 5672
rect 15653 5614 21055 5616
rect 15653 5611 15719 5614
rect 20989 5611 21055 5614
rect 21176 5614 22202 5674
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 20662 5340 20668 5404
rect 20732 5402 20738 5404
rect 20989 5402 21055 5405
rect 20732 5400 21055 5402
rect 20732 5344 20994 5400
rect 21050 5344 21055 5400
rect 20732 5342 21055 5344
rect 20732 5340 20738 5342
rect 20989 5339 21055 5342
rect 17677 5268 17743 5269
rect 17677 5266 17724 5268
rect 17632 5264 17724 5266
rect 17632 5208 17682 5264
rect 17632 5206 17724 5208
rect 17677 5204 17724 5206
rect 17788 5204 17794 5268
rect 20989 5266 21055 5269
rect 21176 5266 21236 5614
rect 22142 5568 22202 5614
rect 22142 5478 23000 5568
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 22200 5448 23000 5478
rect 21738 5407 22054 5408
rect 20989 5264 21236 5266
rect 20989 5208 20994 5264
rect 21050 5208 21236 5264
rect 20989 5206 21236 5208
rect 17677 5203 17743 5204
rect 20989 5203 21055 5206
rect 21081 5130 21147 5133
rect 22200 5130 23000 5160
rect 21081 5128 23000 5130
rect 21081 5072 21086 5128
rect 21142 5072 23000 5128
rect 21081 5070 23000 5072
rect 21081 5067 21147 5070
rect 22200 5040 23000 5070
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 20621 4722 20687 4725
rect 22200 4722 23000 4752
rect 20621 4720 23000 4722
rect 20621 4664 20626 4720
rect 20682 4664 23000 4720
rect 20621 4662 23000 4664
rect 20621 4659 20687 4662
rect 22200 4632 23000 4662
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 16941 4314 17007 4317
rect 20529 4314 20595 4317
rect 22200 4314 23000 4344
rect 16941 4312 20595 4314
rect 16941 4256 16946 4312
rect 17002 4256 20534 4312
rect 20590 4256 20595 4312
rect 16941 4254 20595 4256
rect 16941 4251 17007 4254
rect 20529 4251 20595 4254
rect 22142 4224 23000 4314
rect 15101 4178 15167 4181
rect 19609 4178 19675 4181
rect 15101 4176 19675 4178
rect 15101 4120 15106 4176
rect 15162 4120 19614 4176
rect 19670 4120 19675 4176
rect 15101 4118 19675 4120
rect 15101 4115 15167 4118
rect 19609 4115 19675 4118
rect 20713 4178 20779 4181
rect 22142 4178 22202 4224
rect 20713 4176 22202 4178
rect 20713 4120 20718 4176
rect 20774 4120 22202 4176
rect 20713 4118 22202 4120
rect 20713 4115 20779 4118
rect 17125 4042 17191 4045
rect 19333 4042 19399 4045
rect 17125 4040 19399 4042
rect 17125 3984 17130 4040
rect 17186 3984 19338 4040
rect 19394 3984 19399 4040
rect 17125 3982 19399 3984
rect 17125 3979 17191 3982
rect 19333 3979 19399 3982
rect 20161 3906 20227 3909
rect 22200 3906 23000 3936
rect 20161 3904 23000 3906
rect 20161 3848 20166 3904
rect 20222 3848 23000 3904
rect 20161 3846 23000 3848
rect 20161 3843 20227 3846
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 22200 3816 23000 3846
rect 19139 3775 19455 3776
rect 18137 3770 18203 3773
rect 18270 3770 18276 3772
rect 18137 3768 18276 3770
rect 18137 3712 18142 3768
rect 18198 3712 18276 3768
rect 18137 3710 18276 3712
rect 18137 3707 18203 3710
rect 18270 3708 18276 3710
rect 18340 3708 18346 3772
rect 19517 3770 19583 3773
rect 19517 3768 21420 3770
rect 19517 3712 19522 3768
rect 19578 3712 21420 3768
rect 19517 3710 21420 3712
rect 19517 3707 19583 3710
rect 17125 3634 17191 3637
rect 20529 3634 20595 3637
rect 17125 3632 20595 3634
rect 17125 3576 17130 3632
rect 17186 3576 20534 3632
rect 20590 3576 20595 3632
rect 17125 3574 20595 3576
rect 17125 3571 17191 3574
rect 20529 3571 20595 3574
rect 16665 3498 16731 3501
rect 20161 3498 20227 3501
rect 16665 3496 20227 3498
rect 16665 3440 16670 3496
rect 16726 3440 20166 3496
rect 20222 3440 20227 3496
rect 16665 3438 20227 3440
rect 16665 3435 16731 3438
rect 20161 3435 20227 3438
rect 18321 3362 18387 3365
rect 21173 3362 21239 3365
rect 18321 3360 21239 3362
rect 18321 3304 18326 3360
rect 18382 3304 21178 3360
rect 21234 3304 21239 3360
rect 18321 3302 21239 3304
rect 18321 3299 18387 3302
rect 21173 3299 21239 3302
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 17033 3226 17099 3229
rect 19333 3226 19399 3229
rect 17033 3224 19399 3226
rect 17033 3168 17038 3224
rect 17094 3168 19338 3224
rect 19394 3168 19399 3224
rect 17033 3166 19399 3168
rect 17033 3163 17099 3166
rect 19333 3163 19399 3166
rect 16665 3090 16731 3093
rect 19885 3090 19951 3093
rect 16665 3088 19951 3090
rect 16665 3032 16670 3088
rect 16726 3032 19890 3088
rect 19946 3032 19951 3088
rect 16665 3030 19951 3032
rect 21360 3090 21420 3710
rect 21633 3498 21699 3501
rect 22200 3498 23000 3528
rect 21633 3496 23000 3498
rect 21633 3440 21638 3496
rect 21694 3440 23000 3496
rect 21633 3438 23000 3440
rect 21633 3435 21699 3438
rect 22200 3408 23000 3438
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 22200 3090 23000 3120
rect 21360 3030 23000 3090
rect 16665 3027 16731 3030
rect 19885 3027 19951 3030
rect 22200 3000 23000 3030
rect 17769 2954 17835 2957
rect 19006 2954 19012 2956
rect 17769 2952 19012 2954
rect 17769 2896 17774 2952
rect 17830 2896 19012 2952
rect 17769 2894 19012 2896
rect 17769 2891 17835 2894
rect 19006 2892 19012 2894
rect 19076 2954 19082 2956
rect 19333 2954 19399 2957
rect 19076 2952 19399 2954
rect 19076 2896 19338 2952
rect 19394 2896 19399 2952
rect 19076 2894 19399 2896
rect 19076 2892 19082 2894
rect 19333 2891 19399 2894
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 21541 2682 21607 2685
rect 22200 2682 23000 2712
rect 21541 2680 23000 2682
rect 21541 2624 21546 2680
rect 21602 2624 23000 2680
rect 21541 2622 23000 2624
rect 21541 2619 21607 2622
rect 22200 2592 23000 2622
rect 18781 2546 18847 2549
rect 21357 2546 21423 2549
rect 18781 2544 21423 2546
rect 18781 2488 18786 2544
rect 18842 2488 21362 2544
rect 21418 2488 21423 2544
rect 18781 2486 21423 2488
rect 18781 2483 18847 2486
rect 21357 2483 21423 2486
rect 18965 2410 19031 2413
rect 18965 2408 22202 2410
rect 18965 2352 18970 2408
rect 19026 2352 22202 2408
rect 18965 2350 22202 2352
rect 18965 2347 19031 2350
rect 22142 2304 22202 2350
rect 22142 2214 23000 2304
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 22200 2184 23000 2214
rect 21738 2143 22054 2144
rect 21357 1866 21423 1869
rect 22200 1866 23000 1896
rect 21357 1864 23000 1866
rect 21357 1808 21362 1864
rect 21418 1808 23000 1864
rect 21357 1806 23000 1808
rect 21357 1803 21423 1806
rect 22200 1776 23000 1806
rect 19885 1458 19951 1461
rect 22200 1458 23000 1488
rect 19885 1456 23000 1458
rect 19885 1400 19890 1456
rect 19946 1400 23000 1456
rect 19885 1398 23000 1400
rect 19885 1395 19951 1398
rect 22200 1368 23000 1398
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 19564 18124 19628 18188
rect 20668 18124 20732 18188
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 17724 16492 17788 16556
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 16252 14512 16316 14516
rect 16252 14456 16302 14512
rect 16302 14456 16316 14512
rect 16252 14452 16316 14456
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 15332 11188 15396 11252
rect 16252 11188 16316 11252
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 19012 8392 19076 8396
rect 19012 8336 19062 8392
rect 19062 8336 19076 8392
rect 19012 8332 19076 8336
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 19564 7440 19628 7444
rect 19564 7384 19578 7440
rect 19578 7384 19628 7440
rect 19564 7380 19628 7384
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 18276 6972 18340 7036
rect 15332 6896 15396 6900
rect 15332 6840 15346 6896
rect 15346 6840 15396 6896
rect 15332 6836 15396 6840
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 20668 5340 20732 5404
rect 17724 5264 17788 5268
rect 17724 5208 17738 5264
rect 17738 5208 17788 5264
rect 17724 5204 17788 5208
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 18276 3708 18340 3772
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 19012 2892 19076 2956
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 19563 18188 19629 18189
rect 19563 18124 19564 18188
rect 19628 18124 19629 18188
rect 19563 18123 19629 18124
rect 20667 18188 20733 18189
rect 20667 18124 20668 18188
rect 20732 18124 20733 18188
rect 20667 18123 20733 18124
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 17723 16556 17789 16557
rect 17723 16492 17724 16556
rect 17788 16492 17789 16556
rect 17723 16491 17789 16492
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16251 14516 16317 14517
rect 16251 14452 16252 14516
rect 16316 14452 16317 14516
rect 16251 14451 16317 14452
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 16254 11253 16314 14451
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 15331 11252 15397 11253
rect 15331 11188 15332 11252
rect 15396 11188 15397 11252
rect 15331 11187 15397 11188
rect 16251 11252 16317 11253
rect 16251 11188 16252 11252
rect 16316 11188 16317 11252
rect 16251 11187 16317 11188
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 15334 6901 15394 11187
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 15331 6900 15397 6901
rect 15331 6836 15332 6900
rect 15396 6836 15397 6900
rect 15331 6835 15397 6836
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 17726 5269 17786 16491
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19011 8396 19077 8397
rect 19011 8332 19012 8396
rect 19076 8332 19077 8396
rect 19011 8331 19077 8332
rect 18275 7036 18341 7037
rect 18275 6972 18276 7036
rect 18340 6972 18341 7036
rect 18275 6971 18341 6972
rect 17723 5268 17789 5269
rect 17723 5204 17724 5268
rect 17788 5204 17789 5268
rect 17723 5203 17789 5204
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 18278 3773 18338 6971
rect 18275 3772 18341 3773
rect 18275 3708 18276 3772
rect 18340 3708 18341 3772
rect 18275 3707 18341 3708
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 19014 2957 19074 8331
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19566 7445 19626 18123
rect 19563 7444 19629 7445
rect 19563 7380 19564 7444
rect 19628 7380 19629 7444
rect 19563 7379 19629 7380
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 20670 5405 20730 18123
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 20667 5404 20733 5405
rect 20667 5340 20668 5404
rect 20732 5340 20733 5404
rect 20667 5339 20733 5340
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19011 2956 19077 2957
rect 19011 2892 19012 2956
rect 19076 2892 19077 2956
rect 19011 2891 19077 2892
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 17756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform -1 0 18216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform -1 0 16744 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1649977179
transform -1 0 17112 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1649977179
transform -1 0 18124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1649977179
transform -1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1649977179
transform -1 0 17204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1649977179
transform -1 0 18492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1649977179
transform -1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1649977179
transform -1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1649977179
transform -1 0 17020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1649977179
transform -1 0 18584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1649977179
transform -1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1649977179
transform -1 0 17112 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__87__A
timestamp 1649977179
transform -1 0 17480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__88__A
timestamp 1649977179
transform 1 0 21252 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 19504 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 19964 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 20608 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 20332 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 15088 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 18032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 20884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 15088 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 21344 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 18768 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 19872 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 19964 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 18768 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 15272 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 17480 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14536 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 19596 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18676 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 18400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 19688 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18676 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 19964 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 15272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 15272 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 11224 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12236 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14628 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 12236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13248 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13248 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9292 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17480 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 19780 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 17296 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_174 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17112 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1649977179
transform 1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_186
timestamp 1649977179
transform 1 0 18216 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_190
timestamp 1649977179
transform 1 0 18584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1649977179
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_212
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1649977179
transform 1 0 21160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1649977179
transform 1 0 21528 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_135
timestamp 1649977179
transform 1 0 13524 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_147
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_185
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_189
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_211
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_218
timestamp 1649977179
transform 1 0 21160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_222
timestamp 1649977179
transform 1 0 21528 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_170
timestamp 1649977179
transform 1 0 16744 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_174
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_180
timestamp 1649977179
transform 1 0 17664 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_184
timestamp 1649977179
transform 1 0 18032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1649977179
transform 1 0 19596 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_211
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_216
timestamp 1649977179
transform 1 0 20976 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_220
timestamp 1649977179
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_149 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_157
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_162
timestamp 1649977179
transform 1 0 16008 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_171
timestamp 1649977179
transform 1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_175
timestamp 1649977179
transform 1 0 17204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_179
timestamp 1649977179
transform 1 0 17572 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_190
timestamp 1649977179
transform 1 0 18584 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_194
timestamp 1649977179
transform 1 0 18952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1649977179
transform 1 0 19504 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_206
timestamp 1649977179
transform 1 0 20056 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_212
timestamp 1649977179
transform 1 0 20608 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_218
timestamp 1649977179
transform 1 0 21160 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_222
timestamp 1649977179
transform 1 0 21528 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1649977179
transform 1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_160
timestamp 1649977179
transform 1 0 15824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_169
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_173
timestamp 1649977179
transform 1 0 17020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_186
timestamp 1649977179
transform 1 0 18216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1649977179
transform 1 0 18584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1649977179
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_199
timestamp 1649977179
transform 1 0 19412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_203
timestamp 1649977179
transform 1 0 19780 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_207
timestamp 1649977179
transform 1 0 20148 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_213
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_217
timestamp 1649977179
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_154
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_158
timestamp 1649977179
transform 1 0 15640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_162
timestamp 1649977179
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_175
timestamp 1649977179
transform 1 0 17204 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_187
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_194
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_198
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_202
timestamp 1649977179
transform 1 0 19688 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_206
timestamp 1649977179
transform 1 0 20056 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_210
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1649977179
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_147
timestamp 1649977179
transform 1 0 14628 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_151
timestamp 1649977179
transform 1 0 14996 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1649977179
transform 1 0 15272 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_170
timestamp 1649977179
transform 1 0 16744 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_182
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_178
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_198
timestamp 1649977179
transform 1 0 19320 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_209
timestamp 1649977179
transform 1 0 20332 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_220
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_145
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_148
timestamp 1649977179
transform 1 0 14720 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_152
timestamp 1649977179
transform 1 0 15088 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_157
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_168
timestamp 1649977179
transform 1 0 16560 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_179
timestamp 1649977179
transform 1 0 17572 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1649977179
transform 1 0 18584 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_206
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_210
timestamp 1649977179
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_131
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_134
timestamp 1649977179
transform 1 0 13432 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp 1649977179
transform 1 0 14444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_153
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1649977179
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_172
timestamp 1649977179
transform 1 0 16928 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_185
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_196
timestamp 1649977179
transform 1 0 19136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_207
timestamp 1649977179
transform 1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_47
timestamp 1649977179
transform 1 0 5428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1649977179
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_56
timestamp 1649977179
transform 1 0 6256 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_68
timestamp 1649977179
transform 1 0 7360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_150
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1649977179
transform 1 0 15272 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_158
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_163
timestamp 1649977179
transform 1 0 16100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_168
timestamp 1649977179
transform 1 0 16560 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_176
timestamp 1649977179
transform 1 0 17296 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1649977179
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_203
timestamp 1649977179
transform 1 0 19780 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_207
timestamp 1649977179
transform 1 0 20148 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_218
timestamp 1649977179
transform 1 0 21160 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_222
timestamp 1649977179
transform 1 0 21528 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_140
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_151
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1649977179
transform 1 0 15364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_178
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_189
timestamp 1649977179
transform 1 0 18492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1649977179
transform 1 0 19504 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_211
timestamp 1649977179
transform 1 0 20516 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_218
timestamp 1649977179
transform 1 0 21160 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_222
timestamp 1649977179
transform 1 0 21528 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_147
timestamp 1649977179
transform 1 0 14628 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_159
timestamp 1649977179
transform 1 0 15732 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_169
timestamp 1649977179
transform 1 0 16652 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_174
timestamp 1649977179
transform 1 0 17112 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_180
timestamp 1649977179
transform 1 0 17664 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1649977179
transform 1 0 19780 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1649977179
transform 1 0 20516 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1649977179
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1649977179
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_117
timestamp 1649977179
transform 1 0 11868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_128
timestamp 1649977179
transform 1 0 12880 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_134
timestamp 1649977179
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_138
timestamp 1649977179
transform 1 0 13800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_150
timestamp 1649977179
transform 1 0 14904 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_154
timestamp 1649977179
transform 1 0 15272 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_172
timestamp 1649977179
transform 1 0 16928 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1649977179
transform 1 0 17664 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 1649977179
transform 1 0 19136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_207
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_132
timestamp 1649977179
transform 1 0 13248 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_150
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_155
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_159
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_170
timestamp 1649977179
transform 1 0 16744 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_182
timestamp 1649977179
transform 1 0 17848 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_187
timestamp 1649977179
transform 1 0 18308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1649977179
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_203
timestamp 1649977179
transform 1 0 19780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_207
timestamp 1649977179
transform 1 0 20148 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1649977179
transform 1 0 20608 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1649977179
transform 1 0 21160 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_222
timestamp 1649977179
transform 1 0 21528 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1649977179
transform 1 0 12420 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_127
timestamp 1649977179
transform 1 0 12788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_131
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_134
timestamp 1649977179
transform 1 0 13432 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_146
timestamp 1649977179
transform 1 0 14536 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_154
timestamp 1649977179
transform 1 0 15272 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1649977179
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_178
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_189
timestamp 1649977179
transform 1 0 18492 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1649977179
transform 1 0 19504 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_211
timestamp 1649977179
transform 1 0 20516 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_218
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_222
timestamp 1649977179
transform 1 0 21528 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_105
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_110
timestamp 1649977179
transform 1 0 11224 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_132
timestamp 1649977179
transform 1 0 13248 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_150
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 1649977179
transform 1 0 15272 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_164
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_169
timestamp 1649977179
transform 1 0 16652 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_181
timestamp 1649977179
transform 1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_186
timestamp 1649977179
transform 1 0 18216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_190
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1649977179
transform 1 0 19596 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_205
timestamp 1649977179
transform 1 0 19964 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1649977179
transform 1 0 20700 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1649977179
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_222
timestamp 1649977179
transform 1 0 21528 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_121
timestamp 1649977179
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_133
timestamp 1649977179
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_138
timestamp 1649977179
transform 1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1649977179
transform 1 0 14260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1649977179
transform 1 0 14996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1649977179
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1649977179
transform 1 0 16928 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_183
timestamp 1649977179
transform 1 0 17940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_191
timestamp 1649977179
transform 1 0 18676 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_207
timestamp 1649977179
transform 1 0 20148 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_213
timestamp 1649977179
transform 1 0 20700 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_218
timestamp 1649977179
transform 1 0 21160 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_222
timestamp 1649977179
transform 1 0 21528 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_150
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_168
timestamp 1649977179
transform 1 0 16560 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_172
timestamp 1649977179
transform 1 0 16928 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_179
timestamp 1649977179
transform 1 0 17572 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1649977179
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1649977179
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_207
timestamp 1649977179
transform 1 0 20148 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_213
timestamp 1649977179
transform 1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1649977179
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_145
timestamp 1649977179
transform 1 0 14444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_191
timestamp 1649977179
transform 1 0 18676 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1649977179
transform 1 0 19780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_159
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_167
timestamp 1649977179
transform 1 0 16468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_186
timestamp 1649977179
transform 1 0 18216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_213
timestamp 1649977179
transform 1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_121
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1649977179
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_185
timestamp 1649977179
transform 1 0 18124 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_203
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_89
timestamp 1649977179
transform 1 0 9292 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_100
timestamp 1649977179
transform 1 0 10304 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_105
timestamp 1649977179
transform 1 0 10764 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_181
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1649977179
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_213
timestamp 1649977179
transform 1 0 20700 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_97
timestamp 1649977179
transform 1 0 10028 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1649977179
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_145
timestamp 1649977179
transform 1 0 14444 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1649977179
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_149
timestamp 1649977179
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_168
timestamp 1649977179
transform 1 0 16560 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_180
timestamp 1649977179
transform 1 0 17664 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_216
timestamp 1649977179
transform 1 0 20976 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_222
timestamp 1649977179
transform 1 0 21528 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1649977179
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1649977179
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_142
timestamp 1649977179
transform 1 0 14168 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_160
timestamp 1649977179
transform 1 0 15824 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_185
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_197
timestamp 1649977179
transform 1 0 19228 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_219
timestamp 1649977179
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_118
timestamp 1649977179
transform 1 0 11960 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_149
timestamp 1649977179
transform 1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_168
timestamp 1649977179
transform 1 0 16560 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_174
timestamp 1649977179
transform 1 0 17112 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_191
timestamp 1649977179
transform 1 0 18676 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_199
timestamp 1649977179
transform 1 0 19412 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1649977179
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_220
timestamp 1649977179
transform 1 0 21344 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_122
timestamp 1649977179
transform 1 0 12328 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_159
timestamp 1649977179
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_177
timestamp 1649977179
transform 1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_196
timestamp 1649977179
transform 1 0 19136 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_202
timestamp 1649977179
transform 1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_182
timestamp 1649977179
transform 1 0 17848 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1649977179
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_203
timestamp 1649977179
transform 1 0 19780 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_220
timestamp 1649977179
transform 1 0 21344 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_143
timestamp 1649977179
transform 1 0 14260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_155
timestamp 1649977179
transform 1 0 15364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_197
timestamp 1649977179
transform 1 0 19228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_214
timestamp 1649977179
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_222
timestamp 1649977179
transform 1 0 21528 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_100
timestamp 1649977179
transform 1 0 10304 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_111
timestamp 1649977179
transform 1 0 11316 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_119
timestamp 1649977179
transform 1 0 12052 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_157
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_175
timestamp 1649977179
transform 1 0 17204 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1649977179
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_213
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_102
timestamp 1649977179
transform 1 0 10488 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1649977179
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1649977179
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_142
timestamp 1649977179
transform 1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_160
timestamp 1649977179
transform 1 0 15824 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1649977179
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_185
timestamp 1649977179
transform 1 0 18124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1649977179
transform 1 0 19780 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_35
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_47
timestamp 1649977179
transform 1 0 5428 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_56
timestamp 1649977179
transform 1 0 6256 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_62
timestamp 1649977179
transform 1 0 6808 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_74
timestamp 1649977179
transform 1 0 7912 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1649977179
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_101
timestamp 1649977179
transform 1 0 10396 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_116
timestamp 1649977179
transform 1 0 11776 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_128
timestamp 1649977179
transform 1 0 12880 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_157
timestamp 1649977179
transform 1 0 15548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_161
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_178
timestamp 1649977179
transform 1 0 17480 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_213
timestamp 1649977179
transform 1 0 20700 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_219
timestamp 1649977179
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_157
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1649977179
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_176
timestamp 1649977179
transform 1 0 17296 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_214
timestamp 1649977179
transform 1 0 20792 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_220
timestamp 1649977179
transform 1 0 21344 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _24_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1649977179
transform -1 0 14628 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1649977179
transform -1 0 11960 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1649977179
transform -1 0 11316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1649977179
transform 1 0 17940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1649977179
transform -1 0 19320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1649977179
transform -1 0 15548 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1649977179
transform 1 0 15824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1649977179
transform -1 0 16652 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1649977179
transform 1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1649977179
transform 1 0 18032 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1649977179
transform 1 0 18676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1649977179
transform -1 0 19136 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1649977179
transform 1 0 15088 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1649977179
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1649977179
transform -1 0 14260 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1649977179
transform 1 0 16468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _48_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1649977179
transform 1 0 20792 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1649977179
transform 1 0 20792 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1649977179
transform 1 0 20884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1649977179
transform 1 0 20792 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1649977179
transform 1 0 20792 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1649977179
transform 1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1649977179
transform 1 0 20792 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1649977179
transform 1 0 20884 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1649977179
transform 1 0 16008 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1649977179
transform -1 0 4324 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1649977179
transform -1 0 5428 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1649977179
transform -1 0 6808 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1649977179
transform 1 0 20976 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1649977179
transform -1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1649977179
transform -1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1649977179
transform -1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1649977179
transform -1 0 19872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1649977179
transform -1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1649977179
transform -1 0 20976 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1649977179
transform -1 0 21160 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1649977179
transform -1 0 20700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1649977179
transform -1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1649977179
transform -1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1649977179
transform -1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1649977179
transform -1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1649977179
transform 1 0 17296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1649977179
transform -1 0 19964 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1649977179
transform -1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1649977179
transform -1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1649977179
transform -1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1649977179
transform -1 0 21160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1649977179
transform -1 0 21160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1649977179
transform -1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18860 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17848 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16008 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20700 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17480 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19872 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20884 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17756 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20792 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19504 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19780 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21344 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20792 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19872 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18308 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18676 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16192 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18216 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15732 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13892 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14444 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12696 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15732 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14352 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19780 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14168 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12328 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14260 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14260 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15088 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16560 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14352 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17388 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19136 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16928 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19688 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15824 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14812 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18676 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17020 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17756 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15732 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20516 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20516 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 18584 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19504 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 18952 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20148 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19964 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18216 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18492 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 16284 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 19136 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20608 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20608 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 19504 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 20056 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20516 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20516 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16376 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17572 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 16100 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 17664 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17940 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18492 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 16376 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18676 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17848 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19320 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14720 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12880 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12236 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17020 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12420 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13340 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19596 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15364 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17296 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 14996 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15824 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16560 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17756 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10120 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6256 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13616 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9844 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12420 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11776 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12420 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10488 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10672 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10304 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9660 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17664 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17112 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16192 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18952 0 1 19584
box -38 -48 1142 592
<< labels >>
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 SC_IN_TOP
port 0 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 1 nsew signal tristate
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_1_
port 4 nsew signal input
flabel metal2 s 17222 22200 17278 23000 0 FreeSans 224 90 0 0 ccff_head
port 5 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 ccff_tail
port 6 nsew signal tristate
flabel metal3 s 22200 4632 23000 4752 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 7 nsew signal input
flabel metal3 s 22200 8712 23000 8832 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 8 nsew signal input
flabel metal3 s 22200 9120 23000 9240 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 9 nsew signal input
flabel metal3 s 22200 9528 23000 9648 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 10 nsew signal input
flabel metal3 s 22200 9936 23000 10056 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 11 nsew signal input
flabel metal3 s 22200 10344 23000 10464 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 12 nsew signal input
flabel metal3 s 22200 10752 23000 10872 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 13 nsew signal input
flabel metal3 s 22200 11160 23000 11280 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 14 nsew signal input
flabel metal3 s 22200 11568 23000 11688 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 15 nsew signal input
flabel metal3 s 22200 11976 23000 12096 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 16 nsew signal input
flabel metal3 s 22200 12384 23000 12504 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 17 nsew signal input
flabel metal3 s 22200 5040 23000 5160 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 18 nsew signal input
flabel metal3 s 22200 5448 23000 5568 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 19 nsew signal input
flabel metal3 s 22200 5856 23000 5976 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 20 nsew signal input
flabel metal3 s 22200 6264 23000 6384 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 21 nsew signal input
flabel metal3 s 22200 6672 23000 6792 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 22 nsew signal input
flabel metal3 s 22200 7080 23000 7200 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 23 nsew signal input
flabel metal3 s 22200 7488 23000 7608 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 24 nsew signal input
flabel metal3 s 22200 7896 23000 8016 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 25 nsew signal input
flabel metal3 s 22200 8304 23000 8424 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 26 nsew signal input
flabel metal3 s 22200 12792 23000 12912 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 27 nsew signal tristate
flabel metal3 s 22200 16872 23000 16992 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 28 nsew signal tristate
flabel metal3 s 22200 17280 23000 17400 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 29 nsew signal tristate
flabel metal3 s 22200 17688 23000 17808 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 30 nsew signal tristate
flabel metal3 s 22200 18096 23000 18216 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 31 nsew signal tristate
flabel metal3 s 22200 18504 23000 18624 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 32 nsew signal tristate
flabel metal3 s 22200 18912 23000 19032 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 33 nsew signal tristate
flabel metal3 s 22200 19320 23000 19440 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 34 nsew signal tristate
flabel metal3 s 22200 19728 23000 19848 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 35 nsew signal tristate
flabel metal3 s 22200 20136 23000 20256 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 36 nsew signal tristate
flabel metal3 s 22200 20544 23000 20664 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 37 nsew signal tristate
flabel metal3 s 22200 13200 23000 13320 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 38 nsew signal tristate
flabel metal3 s 22200 13608 23000 13728 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 39 nsew signal tristate
flabel metal3 s 22200 14016 23000 14136 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 40 nsew signal tristate
flabel metal3 s 22200 14424 23000 14544 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 41 nsew signal tristate
flabel metal3 s 22200 14832 23000 14952 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 42 nsew signal tristate
flabel metal3 s 22200 15240 23000 15360 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 43 nsew signal tristate
flabel metal3 s 22200 15648 23000 15768 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 44 nsew signal tristate
flabel metal3 s 22200 16056 23000 16176 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 45 nsew signal tristate
flabel metal3 s 22200 16464 23000 16584 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 46 nsew signal tristate
flabel metal2 s 2502 0 2558 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 47 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 48 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 49 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 50 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 51 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 52 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 53 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 54 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 55 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 56 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 57 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 58 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 59 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 60 nsew signal input
flabel metal2 s 4342 0 4398 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 61 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 62 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 63 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 64 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 65 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 66 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 67 nsew signal tristate
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 68 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 69 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 70 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 71 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 72 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 73 nsew signal tristate
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 74 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 75 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 76 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 77 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 78 nsew signal tristate
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 79 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 80 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 81 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 82 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 83 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 84 nsew signal tristate
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 85 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 86 nsew signal tristate
flabel metal3 s 22200 20952 23000 21072 0 FreeSans 480 0 0 0 prog_clk_0_E_in
port 87 nsew signal input
flabel metal3 s 22200 1368 23000 1488 0 FreeSans 480 0 0 0 right_bottom_grid_pin_34_
port 88 nsew signal input
flabel metal3 s 22200 1776 23000 1896 0 FreeSans 480 0 0 0 right_bottom_grid_pin_35_
port 89 nsew signal input
flabel metal3 s 22200 2184 23000 2304 0 FreeSans 480 0 0 0 right_bottom_grid_pin_36_
port 90 nsew signal input
flabel metal3 s 22200 2592 23000 2712 0 FreeSans 480 0 0 0 right_bottom_grid_pin_37_
port 91 nsew signal input
flabel metal3 s 22200 3000 23000 3120 0 FreeSans 480 0 0 0 right_bottom_grid_pin_38_
port 92 nsew signal input
flabel metal3 s 22200 3408 23000 3528 0 FreeSans 480 0 0 0 right_bottom_grid_pin_39_
port 93 nsew signal input
flabel metal3 s 22200 3816 23000 3936 0 FreeSans 480 0 0 0 right_bottom_grid_pin_40_
port 94 nsew signal input
flabel metal3 s 22200 4224 23000 4344 0 FreeSans 480 0 0 0 right_bottom_grid_pin_41_
port 95 nsew signal input
flabel metal3 s 22200 21360 23000 21480 0 FreeSans 480 0 0 0 right_top_grid_pin_1_
port 96 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
