magic
tech sky130A
magscale 1 2
timestamp 1680087882
<< viali >>
rect 6561 24361 6595 24395
rect 15025 24361 15059 24395
rect 16957 24361 16991 24395
rect 21925 24361 21959 24395
rect 24409 24361 24443 24395
rect 9137 24293 9171 24327
rect 11713 24293 11747 24327
rect 15577 24293 15611 24327
rect 18153 24293 18187 24327
rect 3249 24225 3283 24259
rect 8217 24225 8251 24259
rect 10977 24225 11011 24259
rect 12817 24225 12851 24259
rect 16037 24225 16071 24259
rect 16221 24225 16255 24259
rect 17601 24225 17635 24259
rect 18797 24225 18831 24259
rect 25145 24225 25179 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 6745 24157 6779 24191
rect 7205 24157 7239 24191
rect 9321 24157 9355 24191
rect 9781 24157 9815 24191
rect 11897 24157 11931 24191
rect 12449 24157 12483 24191
rect 15945 24157 15979 24191
rect 20269 24157 20303 24191
rect 21005 24157 21039 24191
rect 22293 24157 22327 24191
rect 24961 24157 24995 24191
rect 5825 24089 5859 24123
rect 14933 24089 14967 24123
rect 19441 24089 19475 24123
rect 22569 24089 22603 24123
rect 3985 24021 4019 24055
rect 17325 24021 17359 24055
rect 17417 24021 17451 24055
rect 18521 24021 18555 24055
rect 18613 24021 18647 24055
rect 24041 24021 24075 24055
rect 24593 24021 24627 24055
rect 25053 24021 25087 24055
rect 25421 24021 25455 24055
rect 14105 23817 14139 23851
rect 14473 23817 14507 23851
rect 24317 23817 24351 23851
rect 3985 23749 4019 23783
rect 5825 23749 5859 23783
rect 9137 23749 9171 23783
rect 10885 23749 10919 23783
rect 16037 23749 16071 23783
rect 17233 23749 17267 23783
rect 20085 23749 20119 23783
rect 20269 23749 20303 23783
rect 21833 23749 21867 23783
rect 24777 23749 24811 23783
rect 25145 23749 25179 23783
rect 1685 23681 1719 23715
rect 2145 23681 2179 23715
rect 2973 23681 3007 23715
rect 4813 23681 4847 23715
rect 7941 23681 7975 23715
rect 9781 23681 9815 23715
rect 12081 23681 12115 23715
rect 15853 23681 15887 23715
rect 18061 23681 18095 23715
rect 20637 23681 20671 23715
rect 1869 23613 1903 23647
rect 6561 23613 6595 23647
rect 6837 23613 6871 23647
rect 12541 23613 12575 23647
rect 14565 23613 14599 23647
rect 14749 23613 14783 23647
rect 17325 23613 17359 23647
rect 17509 23613 17543 23647
rect 18337 23613 18371 23647
rect 20913 23613 20947 23647
rect 22293 23613 22327 23647
rect 22569 23613 22603 23647
rect 24041 23613 24075 23647
rect 11621 23545 11655 23579
rect 25329 23545 25363 23579
rect 2513 23477 2547 23511
rect 16405 23477 16439 23511
rect 16865 23477 16899 23511
rect 19809 23477 19843 23511
rect 24593 23477 24627 23511
rect 4261 23205 4295 23239
rect 21189 23205 21223 23239
rect 24593 23205 24627 23239
rect 10517 23137 10551 23171
rect 12173 23137 12207 23171
rect 15301 23137 15335 23171
rect 17693 23137 17727 23171
rect 17877 23137 17911 23171
rect 21649 23137 21683 23171
rect 25145 23137 25179 23171
rect 2237 23069 2271 23103
rect 4077 23069 4111 23103
rect 5457 23069 5491 23103
rect 7205 23069 7239 23103
rect 8217 23069 8251 23103
rect 9413 23069 9447 23103
rect 9873 23069 9907 23103
rect 11713 23069 11747 23103
rect 13737 23069 13771 23103
rect 15025 23069 15059 23103
rect 17601 23069 17635 23103
rect 19441 23069 19475 23103
rect 3249 23001 3283 23035
rect 6377 23001 6411 23035
rect 14381 23001 14415 23035
rect 18521 23001 18555 23035
rect 18705 23001 18739 23035
rect 19717 23001 19751 23035
rect 21925 23001 21959 23035
rect 24501 23001 24535 23035
rect 4721 22933 4755 22967
rect 9229 22933 9263 22967
rect 13553 22933 13587 22967
rect 14473 22933 14507 22967
rect 16773 22933 16807 22967
rect 17233 22933 17267 22967
rect 23397 22933 23431 22967
rect 23857 22933 23891 22967
rect 24961 22933 24995 22967
rect 25053 22933 25087 22967
rect 2513 22729 2547 22763
rect 12081 22729 12115 22763
rect 13093 22729 13127 22763
rect 15393 22729 15427 22763
rect 16405 22729 16439 22763
rect 18613 22729 18647 22763
rect 19073 22729 19107 22763
rect 20269 22729 20303 22763
rect 21281 22729 21315 22763
rect 3985 22661 4019 22695
rect 5733 22661 5767 22695
rect 7297 22661 7331 22695
rect 8769 22661 8803 22695
rect 13921 22661 13955 22695
rect 23581 22661 23615 22695
rect 25329 22661 25363 22695
rect 1685 22593 1719 22627
rect 2145 22593 2179 22627
rect 2973 22593 3007 22627
rect 4813 22593 4847 22627
rect 6653 22593 6687 22627
rect 7573 22593 7607 22627
rect 12173 22593 12207 22627
rect 13001 22593 13035 22627
rect 13645 22593 13679 22627
rect 15945 22593 15979 22627
rect 16129 22593 16163 22627
rect 16865 22593 16899 22627
rect 19441 22593 19475 22627
rect 20637 22593 20671 22627
rect 21649 22593 21683 22627
rect 22017 22593 22051 22627
rect 23305 22593 23339 22627
rect 9413 22525 9447 22559
rect 9689 22525 9723 22559
rect 12265 22525 12299 22559
rect 17141 22525 17175 22559
rect 19533 22525 19567 22559
rect 19625 22525 19659 22559
rect 20729 22525 20763 22559
rect 20821 22525 20855 22559
rect 22293 22525 22327 22559
rect 1869 22457 1903 22491
rect 6745 22389 6779 22423
rect 11161 22389 11195 22423
rect 11713 22389 11747 22423
rect 25053 22389 25087 22423
rect 14552 22185 14586 22219
rect 2881 22049 2915 22083
rect 6101 22049 6135 22083
rect 8309 22049 8343 22083
rect 10701 22049 10735 22083
rect 12449 22049 12483 22083
rect 17049 22049 17083 22083
rect 18245 22049 18279 22083
rect 20637 22049 20671 22083
rect 23489 22049 23523 22083
rect 25053 22049 25087 22083
rect 25145 22049 25179 22083
rect 2237 21981 2271 22015
rect 3985 21981 4019 22015
rect 4261 21981 4295 22015
rect 5549 21981 5583 22015
rect 7389 21981 7423 22015
rect 8953 21981 8987 22015
rect 9505 21981 9539 22015
rect 13737 21981 13771 22015
rect 14289 21981 14323 22015
rect 16957 21981 16991 22015
rect 20361 21981 20395 22015
rect 22753 21981 22787 22015
rect 23213 21981 23247 22015
rect 10977 21913 11011 21947
rect 13553 21913 13587 21947
rect 18061 21913 18095 21947
rect 18705 21913 18739 21947
rect 19533 21913 19567 21947
rect 9321 21845 9355 21879
rect 10057 21845 10091 21879
rect 12725 21845 12759 21879
rect 16037 21845 16071 21879
rect 16497 21845 16531 21879
rect 16865 21845 16899 21879
rect 17693 21845 17727 21879
rect 18153 21845 18187 21879
rect 18889 21845 18923 21879
rect 19625 21845 19659 21879
rect 22109 21845 22143 21879
rect 22569 21845 22603 21879
rect 24593 21845 24627 21879
rect 24961 21845 24995 21879
rect 12633 21641 12667 21675
rect 14289 21641 14323 21675
rect 1685 21573 1719 21607
rect 2145 21573 2179 21607
rect 12725 21573 12759 21607
rect 23121 21573 23155 21607
rect 25421 21573 25455 21607
rect 2973 21505 3007 21539
rect 4813 21505 4847 21539
rect 6745 21505 6779 21539
rect 7389 21505 7423 21539
rect 9045 21505 9079 21539
rect 11069 21505 11103 21539
rect 11253 21505 11287 21539
rect 14197 21505 14231 21539
rect 15393 21505 15427 21539
rect 16405 21505 16439 21539
rect 17417 21505 17451 21539
rect 18245 21505 18279 21539
rect 20821 21505 20855 21539
rect 22385 21505 22419 21539
rect 23397 21505 23431 21539
rect 3525 21437 3559 21471
rect 5089 21437 5123 21471
rect 7665 21437 7699 21471
rect 9321 21437 9355 21471
rect 12909 21437 12943 21471
rect 14381 21437 14415 21471
rect 15485 21437 15519 21471
rect 15669 21437 15703 21471
rect 17509 21437 17543 21471
rect 17601 21437 17635 21471
rect 20913 21437 20947 21471
rect 21097 21437 21131 21471
rect 21557 21437 21591 21471
rect 22477 21437 22511 21471
rect 22661 21437 22695 21471
rect 23673 21437 23707 21471
rect 1869 21369 1903 21403
rect 15025 21369 15059 21403
rect 22017 21369 22051 21403
rect 6561 21301 6595 21335
rect 10793 21301 10827 21335
rect 12265 21301 12299 21335
rect 13829 21301 13863 21335
rect 16129 21301 16163 21335
rect 17049 21301 17083 21335
rect 19533 21301 19567 21335
rect 20453 21301 20487 21335
rect 25145 21301 25179 21335
rect 6377 21097 6411 21131
rect 12909 21097 12943 21131
rect 14473 21097 14507 21131
rect 18889 21097 18923 21131
rect 21189 21097 21223 21131
rect 24041 21097 24075 21131
rect 9965 21029 9999 21063
rect 15485 21029 15519 21063
rect 16681 21029 16715 21063
rect 17877 21029 17911 21063
rect 2789 20961 2823 20995
rect 4445 20961 4479 20995
rect 7389 20961 7423 20995
rect 10609 20961 10643 20995
rect 11161 20961 11195 20995
rect 11437 20961 11471 20995
rect 13737 20961 13771 20995
rect 15945 20961 15979 20995
rect 16037 20961 16071 20995
rect 17233 20961 17267 20995
rect 18337 20961 18371 20995
rect 18521 20961 18555 20995
rect 19717 20961 19751 20995
rect 22201 20961 22235 20995
rect 23397 20961 23431 20995
rect 25145 20961 25179 20995
rect 2237 20893 2271 20927
rect 4169 20893 4203 20927
rect 6009 20893 6043 20927
rect 6929 20893 6963 20927
rect 13553 20893 13587 20927
rect 19441 20893 19475 20927
rect 22017 20893 22051 20927
rect 24961 20893 24995 20927
rect 14381 20825 14415 20859
rect 15853 20825 15887 20859
rect 17049 20825 17083 20859
rect 18245 20825 18279 20859
rect 22109 20825 22143 20859
rect 22661 20825 22695 20859
rect 23213 20825 23247 20859
rect 23305 20825 23339 20859
rect 23949 20825 23983 20859
rect 5825 20757 5859 20791
rect 9321 20757 9355 20791
rect 10333 20757 10367 20791
rect 10425 20757 10459 20791
rect 17141 20757 17175 20791
rect 21649 20757 21683 20791
rect 22845 20757 22879 20791
rect 24593 20757 24627 20791
rect 25053 20757 25087 20791
rect 2237 20553 2271 20587
rect 5089 20553 5123 20587
rect 5181 20553 5215 20587
rect 7757 20553 7791 20587
rect 12081 20553 12115 20587
rect 12449 20553 12483 20587
rect 12541 20553 12575 20587
rect 18705 20553 18739 20587
rect 21005 20553 21039 20587
rect 22109 20553 22143 20587
rect 4905 20485 4939 20519
rect 11161 20485 11195 20519
rect 13093 20485 13127 20519
rect 22477 20485 22511 20519
rect 23765 20485 23799 20519
rect 1777 20417 1811 20451
rect 2421 20417 2455 20451
rect 3065 20417 3099 20451
rect 6009 20417 6043 20451
rect 7297 20417 7331 20451
rect 8585 20417 8619 20451
rect 9045 20417 9079 20451
rect 15853 20417 15887 20451
rect 16957 20417 16991 20451
rect 23489 20417 23523 20451
rect 3341 20349 3375 20383
rect 9321 20349 9355 20383
rect 12633 20349 12667 20383
rect 13553 20349 13587 20383
rect 13829 20349 13863 20383
rect 17233 20349 17267 20383
rect 19257 20349 19291 20383
rect 19533 20349 19567 20383
rect 22569 20349 22603 20383
rect 22661 20349 22695 20383
rect 23213 20349 23247 20383
rect 1593 20213 1627 20247
rect 5825 20213 5859 20247
rect 7113 20213 7147 20247
rect 8401 20213 8435 20247
rect 10793 20213 10827 20247
rect 15301 20213 15335 20247
rect 15945 20213 15979 20247
rect 16313 20213 16347 20247
rect 21281 20213 21315 20247
rect 21465 20213 21499 20247
rect 25237 20213 25271 20247
rect 10425 20009 10459 20043
rect 14933 20009 14967 20043
rect 17325 20009 17359 20043
rect 17693 20009 17727 20043
rect 18889 20009 18923 20043
rect 20729 20009 20763 20043
rect 22845 20009 22879 20043
rect 24593 20009 24627 20043
rect 13369 19941 13403 19975
rect 13645 19941 13679 19975
rect 13829 19941 13863 19975
rect 16865 19941 16899 19975
rect 18797 19941 18831 19975
rect 2513 19873 2547 19907
rect 10885 19873 10919 19907
rect 10977 19873 11011 19907
rect 15485 19873 15519 19907
rect 18245 19873 18279 19907
rect 19993 19873 20027 19907
rect 21097 19873 21131 19907
rect 23949 19873 23983 19907
rect 25145 19873 25179 19907
rect 2237 19805 2271 19839
rect 4721 19805 4755 19839
rect 5181 19805 5215 19839
rect 5457 19805 5491 19839
rect 6653 19805 6687 19839
rect 7113 19805 7147 19839
rect 7389 19805 7423 19839
rect 11621 19805 11655 19839
rect 14289 19805 14323 19839
rect 17049 19805 17083 19839
rect 18153 19805 18187 19839
rect 25053 19805 25087 19839
rect 8401 19737 8435 19771
rect 10793 19737 10827 19771
rect 11897 19737 11931 19771
rect 15393 19737 15427 19771
rect 16221 19737 16255 19771
rect 19809 19737 19843 19771
rect 21373 19737 21407 19771
rect 23765 19737 23799 19771
rect 24961 19737 24995 19771
rect 4537 19669 4571 19703
rect 6469 19669 6503 19703
rect 9137 19669 9171 19703
rect 9781 19669 9815 19703
rect 15301 19669 15335 19703
rect 16313 19669 16347 19703
rect 18061 19669 18095 19703
rect 19441 19669 19475 19703
rect 19901 19669 19935 19703
rect 23121 19669 23155 19703
rect 23305 19669 23339 19703
rect 23673 19669 23707 19703
rect 3893 19465 3927 19499
rect 5825 19465 5859 19499
rect 7113 19465 7147 19499
rect 11069 19465 11103 19499
rect 11621 19465 11655 19499
rect 11713 19465 11747 19499
rect 14473 19465 14507 19499
rect 14933 19465 14967 19499
rect 15301 19465 15335 19499
rect 18797 19465 18831 19499
rect 19625 19465 19659 19499
rect 20453 19465 20487 19499
rect 20821 19465 20855 19499
rect 22017 19465 22051 19499
rect 22385 19465 22419 19499
rect 22477 19465 22511 19499
rect 25053 19465 25087 19499
rect 9321 19397 9355 19431
rect 15393 19397 15427 19431
rect 20913 19397 20947 19431
rect 1961 19329 1995 19363
rect 4077 19329 4111 19363
rect 4813 19329 4847 19363
rect 6009 19329 6043 19363
rect 7297 19329 7331 19363
rect 7941 19329 7975 19363
rect 8585 19329 8619 19363
rect 9045 19329 9079 19363
rect 12725 19329 12759 19363
rect 16313 19329 16347 19363
rect 17049 19329 17083 19363
rect 19717 19329 19751 19363
rect 23305 19329 23339 19363
rect 2237 19261 2271 19295
rect 4537 19261 4571 19295
rect 6469 19261 6503 19295
rect 6653 19261 6687 19295
rect 6837 19261 6871 19295
rect 12081 19261 12115 19295
rect 13001 19261 13035 19295
rect 15577 19261 15611 19295
rect 16773 19261 16807 19295
rect 17325 19261 17359 19295
rect 19901 19261 19935 19295
rect 21005 19261 21039 19295
rect 22569 19261 22603 19295
rect 23581 19261 23615 19295
rect 25329 19261 25363 19295
rect 7757 19193 7791 19227
rect 8401 19193 8435 19227
rect 10793 19125 10827 19159
rect 11253 19125 11287 19159
rect 16129 19125 16163 19159
rect 19257 19125 19291 19159
rect 21557 19125 21591 19159
rect 1961 18921 1995 18955
rect 3801 18921 3835 18955
rect 4261 18921 4295 18955
rect 5825 18921 5859 18955
rect 8401 18921 8435 18955
rect 9229 18921 9263 18955
rect 13001 18921 13035 18955
rect 14289 18921 14323 18955
rect 17693 18921 17727 18955
rect 2605 18853 2639 18887
rect 18061 18853 18095 18887
rect 7389 18785 7423 18819
rect 9781 18785 9815 18819
rect 13645 18785 13679 18819
rect 14749 18785 14783 18819
rect 14933 18785 14967 18819
rect 15485 18785 15519 18819
rect 17233 18785 17267 18819
rect 18521 18785 18555 18819
rect 18613 18785 18647 18819
rect 19441 18785 19475 18819
rect 20637 18785 20671 18819
rect 23121 18785 23155 18819
rect 23765 18785 23799 18819
rect 25237 18785 25271 18819
rect 1685 18717 1719 18751
rect 2145 18717 2179 18751
rect 2789 18717 2823 18751
rect 3433 18717 3467 18751
rect 4721 18717 4755 18751
rect 5365 18717 5399 18751
rect 6009 18717 6043 18751
rect 6653 18717 6687 18751
rect 7113 18717 7147 18751
rect 8585 18717 8619 18751
rect 9597 18717 9631 18751
rect 13461 18717 13495 18751
rect 20361 18717 20395 18751
rect 25053 18717 25087 18751
rect 10425 18649 10459 18683
rect 13369 18649 13403 18683
rect 14657 18649 14691 18683
rect 15761 18649 15795 18683
rect 22937 18649 22971 18683
rect 23029 18649 23063 18683
rect 3249 18581 3283 18615
rect 4537 18581 4571 18615
rect 5181 18581 5215 18615
rect 6469 18581 6503 18615
rect 9689 18581 9723 18615
rect 11897 18581 11931 18615
rect 17509 18581 17543 18615
rect 18429 18581 18463 18615
rect 22109 18581 22143 18615
rect 22569 18581 22603 18615
rect 24593 18581 24627 18615
rect 24961 18581 24995 18615
rect 1593 18377 1627 18411
rect 2145 18377 2179 18411
rect 2237 18377 2271 18411
rect 4537 18377 4571 18411
rect 5181 18377 5215 18411
rect 5825 18377 5859 18411
rect 8309 18377 8343 18411
rect 11805 18377 11839 18411
rect 12173 18377 12207 18411
rect 15577 18377 15611 18411
rect 15669 18377 15703 18411
rect 18521 18377 18555 18411
rect 23305 18377 23339 18411
rect 25053 18377 25087 18411
rect 6745 18309 6779 18343
rect 11069 18309 11103 18343
rect 11345 18309 11379 18343
rect 14749 18309 14783 18343
rect 20821 18309 20855 18343
rect 20913 18309 20947 18343
rect 1777 18241 1811 18275
rect 2789 18241 2823 18275
rect 2973 18241 3007 18275
rect 3433 18241 3467 18275
rect 4721 18241 4755 18275
rect 5365 18241 5399 18275
rect 6009 18241 6043 18275
rect 7205 18241 7239 18275
rect 7849 18241 7883 18275
rect 8493 18241 8527 18275
rect 8953 18241 8987 18275
rect 12265 18241 12299 18275
rect 13001 18241 13035 18275
rect 17233 18241 17267 18275
rect 17325 18241 17359 18275
rect 18429 18241 18463 18275
rect 19625 18241 19659 18275
rect 22017 18241 22051 18275
rect 24961 18241 24995 18275
rect 3801 18173 3835 18207
rect 3893 18173 3927 18207
rect 6561 18173 6595 18207
rect 9229 18173 9263 18207
rect 12449 18173 12483 18207
rect 15761 18173 15795 18207
rect 17509 18173 17543 18207
rect 18705 18173 18739 18207
rect 19717 18173 19751 18207
rect 19809 18173 19843 18207
rect 21005 18173 21039 18207
rect 21465 18173 21499 18207
rect 24409 18173 24443 18207
rect 25237 18173 25271 18207
rect 7021 18105 7055 18139
rect 15209 18105 15243 18139
rect 16865 18105 16899 18139
rect 3249 18037 3283 18071
rect 7665 18037 7699 18071
rect 10701 18037 10735 18071
rect 16221 18037 16255 18071
rect 18061 18037 18095 18071
rect 19257 18037 19291 18071
rect 20453 18037 20487 18071
rect 24593 18037 24627 18071
rect 3249 17833 3283 17867
rect 6469 17833 6503 17867
rect 7757 17833 7791 17867
rect 11529 17833 11563 17867
rect 13737 17833 13771 17867
rect 17141 17833 17175 17867
rect 20992 17833 21026 17867
rect 22477 17833 22511 17867
rect 16681 17765 16715 17799
rect 5181 17697 5215 17731
rect 5457 17697 5491 17731
rect 9781 17697 9815 17731
rect 11989 17697 12023 17731
rect 12265 17697 12299 17731
rect 14289 17697 14323 17731
rect 14933 17697 14967 17731
rect 15209 17697 15243 17731
rect 17693 17697 17727 17731
rect 19901 17697 19935 17731
rect 20085 17697 20119 17731
rect 20729 17697 20763 17731
rect 23857 17697 23891 17731
rect 3433 17629 3467 17663
rect 4261 17629 4295 17663
rect 4721 17629 4755 17663
rect 6653 17629 6687 17663
rect 7297 17629 7331 17663
rect 7941 17629 7975 17663
rect 8585 17629 8619 17663
rect 9321 17629 9355 17663
rect 17601 17629 17635 17663
rect 18797 17629 18831 17663
rect 23673 17629 23707 17663
rect 23765 17629 23799 17663
rect 10057 17561 10091 17595
rect 22845 17561 22879 17595
rect 24501 17561 24535 17595
rect 24777 17561 24811 17595
rect 24961 17561 24995 17595
rect 4537 17493 4571 17527
rect 7113 17493 7147 17527
rect 8401 17493 8435 17527
rect 9137 17493 9171 17527
rect 17509 17493 17543 17527
rect 18153 17493 18187 17527
rect 18613 17493 18647 17527
rect 19441 17493 19475 17527
rect 19809 17493 19843 17527
rect 22937 17493 22971 17527
rect 23305 17493 23339 17527
rect 3893 17289 3927 17323
rect 6561 17289 6595 17323
rect 7205 17289 7239 17323
rect 7849 17289 7883 17323
rect 15853 17289 15887 17323
rect 20545 17289 20579 17323
rect 24317 17289 24351 17323
rect 9505 17221 9539 17255
rect 11989 17221 12023 17255
rect 3801 17153 3835 17187
rect 4077 17153 4111 17187
rect 6745 17153 6779 17187
rect 7389 17153 7423 17187
rect 8033 17153 8067 17187
rect 8769 17153 8803 17187
rect 9229 17153 9263 17187
rect 11713 17153 11747 17187
rect 14473 17153 14507 17187
rect 15025 17153 15059 17187
rect 17233 17153 17267 17187
rect 18337 17153 18371 17187
rect 21373 17153 21407 17187
rect 22569 17153 22603 17187
rect 24869 17153 24903 17187
rect 4537 17085 4571 17119
rect 4813 17085 4847 17119
rect 10977 17085 11011 17119
rect 13921 17085 13955 17119
rect 15945 17085 15979 17119
rect 16037 17085 16071 17119
rect 17325 17085 17359 17119
rect 17417 17085 17451 17119
rect 18613 17085 18647 17119
rect 20085 17085 20119 17119
rect 21833 17085 21867 17119
rect 22017 17085 22051 17119
rect 22293 17085 22327 17119
rect 22845 17085 22879 17119
rect 8585 17017 8619 17051
rect 13461 17017 13495 17051
rect 14841 17017 14875 17051
rect 17969 17017 18003 17051
rect 25053 17017 25087 17051
rect 11253 16949 11287 16983
rect 15485 16949 15519 16983
rect 16865 16949 16899 16983
rect 21189 16949 21223 16983
rect 6837 16745 6871 16779
rect 7297 16745 7331 16779
rect 16037 16745 16071 16779
rect 16497 16745 16531 16779
rect 7757 16677 7791 16711
rect 9505 16677 9539 16711
rect 5273 16609 5307 16643
rect 7481 16609 7515 16643
rect 9045 16609 9079 16643
rect 11437 16609 11471 16643
rect 12265 16609 12299 16643
rect 14289 16609 14323 16643
rect 17417 16609 17451 16643
rect 19441 16609 19475 16643
rect 22293 16609 22327 16643
rect 22569 16609 22603 16643
rect 24869 16609 24903 16643
rect 4905 16541 4939 16575
rect 7941 16541 7975 16575
rect 8585 16537 8619 16571
rect 9689 16541 9723 16575
rect 11161 16541 11195 16575
rect 11253 16541 11287 16575
rect 11989 16541 12023 16575
rect 16681 16541 16715 16575
rect 17141 16541 17175 16575
rect 9229 16473 9263 16507
rect 14565 16473 14599 16507
rect 19717 16473 19751 16507
rect 24685 16473 24719 16507
rect 4721 16405 4755 16439
rect 8401 16405 8435 16439
rect 10149 16405 10183 16439
rect 10793 16405 10827 16439
rect 13737 16405 13771 16439
rect 18889 16405 18923 16439
rect 21189 16405 21223 16439
rect 21649 16405 21683 16439
rect 24041 16405 24075 16439
rect 8125 16201 8159 16235
rect 10793 16201 10827 16235
rect 10885 16201 10919 16235
rect 14381 16201 14415 16235
rect 19349 16201 19383 16235
rect 21005 16201 21039 16235
rect 23857 16201 23891 16235
rect 11989 16133 12023 16167
rect 15945 16133 15979 16167
rect 19809 16133 19843 16167
rect 20913 16133 20947 16167
rect 22385 16133 22419 16167
rect 24685 16133 24719 16167
rect 8401 16065 8435 16099
rect 8677 16065 8711 16099
rect 9321 16065 9355 16099
rect 9965 16065 9999 16099
rect 14289 16065 14323 16099
rect 15853 16065 15887 16099
rect 17141 16065 17175 16099
rect 19717 16065 19751 16099
rect 21557 16065 21591 16099
rect 23765 16065 23799 16099
rect 11069 15997 11103 16031
rect 11713 15997 11747 16031
rect 13461 15997 13495 16031
rect 14565 15997 14599 16031
rect 16037 15997 16071 16031
rect 19901 15997 19935 16031
rect 21097 15997 21131 16031
rect 22477 15997 22511 16031
rect 22569 15997 22603 16031
rect 23949 15997 23983 16031
rect 9137 15929 9171 15963
rect 9781 15929 9815 15963
rect 10425 15929 10459 15963
rect 15485 15929 15519 15963
rect 23029 15929 23063 15963
rect 24869 15929 24903 15963
rect 8493 15861 8527 15895
rect 13921 15861 13955 15895
rect 15025 15861 15059 15895
rect 16681 15861 16715 15895
rect 18429 15861 18463 15895
rect 20545 15861 20579 15895
rect 22017 15861 22051 15895
rect 23397 15861 23431 15895
rect 8769 15657 8803 15691
rect 9873 15657 9907 15691
rect 18705 15657 18739 15691
rect 16037 15589 16071 15623
rect 16313 15589 16347 15623
rect 10793 15521 10827 15555
rect 13185 15521 13219 15555
rect 13369 15521 13403 15555
rect 14289 15521 14323 15555
rect 16957 15521 16991 15555
rect 17233 15521 17267 15555
rect 20085 15521 20119 15555
rect 21189 15521 21223 15555
rect 21281 15521 21315 15555
rect 22201 15521 22235 15555
rect 9413 15453 9447 15487
rect 10057 15453 10091 15487
rect 10517 15453 10551 15487
rect 13093 15453 13127 15487
rect 19993 15453 20027 15487
rect 21097 15453 21131 15487
rect 22017 15453 22051 15487
rect 23397 15453 23431 15487
rect 24777 15453 24811 15487
rect 14565 15385 14599 15419
rect 16681 15385 16715 15419
rect 19901 15385 19935 15419
rect 22753 15385 22787 15419
rect 9229 15317 9263 15351
rect 12265 15317 12299 15351
rect 12725 15317 12759 15351
rect 13829 15317 13863 15351
rect 18981 15317 19015 15351
rect 19533 15317 19567 15351
rect 20729 15317 20763 15351
rect 22845 15317 22879 15351
rect 24593 15317 24627 15351
rect 9505 15113 9539 15147
rect 9689 15113 9723 15147
rect 10333 15113 10367 15147
rect 24593 15113 24627 15147
rect 9873 15045 9907 15079
rect 13921 15045 13955 15079
rect 15485 15045 15519 15079
rect 16129 15045 16163 15079
rect 17141 15045 17175 15079
rect 21465 15045 21499 15079
rect 22109 15045 22143 15079
rect 23121 15045 23155 15079
rect 10517 14977 10551 15011
rect 11161 14977 11195 15011
rect 14565 14977 14599 15011
rect 15025 14977 15059 15011
rect 10057 14909 10091 14943
rect 11713 14909 11747 14943
rect 11989 14909 12023 14943
rect 13461 14909 13495 14943
rect 16865 14909 16899 14943
rect 19349 14909 19383 14943
rect 19625 14909 19659 14943
rect 21097 14909 21131 14943
rect 22845 14909 22879 14943
rect 25053 14909 25087 14943
rect 10977 14773 11011 14807
rect 14841 14773 14875 14807
rect 18613 14773 18647 14807
rect 19073 14773 19107 14807
rect 22201 14773 22235 14807
rect 10425 14569 10459 14603
rect 12909 14569 12943 14603
rect 20545 14569 20579 14603
rect 22293 14569 22327 14603
rect 25421 14569 25455 14603
rect 18245 14501 18279 14535
rect 19441 14501 19475 14535
rect 22845 14501 22879 14535
rect 25237 14501 25271 14535
rect 10977 14433 11011 14467
rect 12449 14433 12483 14467
rect 13553 14433 13587 14467
rect 14289 14433 14323 14467
rect 14565 14433 14599 14467
rect 16497 14433 16531 14467
rect 16773 14433 16807 14467
rect 19993 14433 20027 14467
rect 23765 14433 23799 14467
rect 23949 14433 23983 14467
rect 10701 14365 10735 14399
rect 13093 14365 13127 14399
rect 20821 14365 20855 14399
rect 23673 14365 23707 14399
rect 19809 14297 19843 14331
rect 19901 14297 19935 14331
rect 24685 14297 24719 14331
rect 16037 14229 16071 14263
rect 18705 14229 18739 14263
rect 23305 14229 23339 14263
rect 24777 14229 24811 14263
rect 11345 14025 11379 14059
rect 15485 14025 15519 14059
rect 16129 14025 16163 14059
rect 17049 14025 17083 14059
rect 17509 14025 17543 14059
rect 19533 14025 19567 14059
rect 20361 14025 20395 14059
rect 21097 14025 21131 14059
rect 11161 13957 11195 13991
rect 18245 13957 18279 13991
rect 23121 13957 23155 13991
rect 25145 13957 25179 13991
rect 11989 13889 12023 13923
rect 12633 13889 12667 13923
rect 13277 13889 13311 13923
rect 13737 13889 13771 13923
rect 15761 13889 15795 13923
rect 16313 13889 16347 13923
rect 17417 13889 17451 13923
rect 22109 13889 22143 13923
rect 22845 13889 22879 13923
rect 16681 13821 16715 13855
rect 17693 13821 17727 13855
rect 21189 13821 21223 13855
rect 21281 13821 21315 13855
rect 24593 13821 24627 13855
rect 25329 13821 25363 13855
rect 11805 13753 11839 13787
rect 12449 13753 12483 13787
rect 13093 13753 13127 13787
rect 22293 13753 22327 13787
rect 14000 13685 14034 13719
rect 20729 13685 20763 13719
rect 13829 13481 13863 13515
rect 16037 13481 16071 13515
rect 18705 13481 18739 13515
rect 21465 13481 21499 13515
rect 24593 13481 24627 13515
rect 13553 13413 13587 13447
rect 19349 13413 19383 13447
rect 23949 13413 23983 13447
rect 24133 13413 24167 13447
rect 14289 13345 14323 13379
rect 16497 13345 16531 13379
rect 16773 13345 16807 13379
rect 19717 13345 19751 13379
rect 21925 13345 21959 13379
rect 25145 13345 25179 13379
rect 9597 13277 9631 13311
rect 11805 13277 11839 13311
rect 18889 13277 18923 13311
rect 25053 13277 25087 13311
rect 12081 13209 12115 13243
rect 14565 13209 14599 13243
rect 19993 13209 20027 13243
rect 22201 13209 22235 13243
rect 24961 13209 24995 13243
rect 10885 13141 10919 13175
rect 18245 13141 18279 13175
rect 23673 13141 23707 13175
rect 12541 12937 12575 12971
rect 14289 12937 14323 12971
rect 15439 12937 15473 12971
rect 23765 12937 23799 12971
rect 24869 12937 24903 12971
rect 13001 12869 13035 12903
rect 16313 12869 16347 12903
rect 21557 12869 21591 12903
rect 15209 12801 15243 12835
rect 19441 12801 19475 12835
rect 20637 12801 20671 12835
rect 22017 12801 22051 12835
rect 24409 12801 24443 12835
rect 16865 12733 16899 12767
rect 17141 12733 17175 12767
rect 19533 12733 19567 12767
rect 19625 12733 19659 12767
rect 20729 12733 20763 12767
rect 20821 12733 20855 12767
rect 21281 12733 21315 12767
rect 22293 12733 22327 12767
rect 18613 12665 18647 12699
rect 24225 12665 24259 12699
rect 19073 12597 19107 12631
rect 20269 12597 20303 12631
rect 25329 12597 25363 12631
rect 13737 12393 13771 12427
rect 13921 12393 13955 12427
rect 15393 12393 15427 12427
rect 17509 12393 17543 12427
rect 24041 12393 24075 12427
rect 25329 12393 25363 12427
rect 14289 12257 14323 12291
rect 15761 12257 15795 12291
rect 17969 12257 18003 12291
rect 18889 12257 18923 12291
rect 19717 12257 19751 12291
rect 22293 12257 22327 12291
rect 22569 12257 22603 12291
rect 24593 12257 24627 12291
rect 14565 12189 14599 12223
rect 19441 12189 19475 12223
rect 21649 12189 21683 12223
rect 16037 12121 16071 12155
rect 18705 12121 18739 12155
rect 21189 12053 21223 12087
rect 25053 12053 25087 12087
rect 14565 11849 14599 11883
rect 15117 11849 15151 11883
rect 15669 11849 15703 11883
rect 19717 11781 19751 11815
rect 23305 11781 23339 11815
rect 12817 11713 12851 11747
rect 15301 11713 15335 11747
rect 16313 11713 16347 11747
rect 17141 11713 17175 11747
rect 19441 11713 19475 11747
rect 21465 11713 21499 11747
rect 22109 11713 22143 11747
rect 23949 11713 23983 11747
rect 13093 11645 13127 11679
rect 17417 11645 17451 11679
rect 24777 11645 24811 11679
rect 16129 11577 16163 11611
rect 21189 11577 21223 11611
rect 16773 11509 16807 11543
rect 18889 11509 18923 11543
rect 14749 11305 14783 11339
rect 15485 11305 15519 11339
rect 16773 11305 16807 11339
rect 17417 11305 17451 11339
rect 18705 11305 18739 11339
rect 22017 11305 22051 11339
rect 16129 11237 16163 11271
rect 19349 11237 19383 11271
rect 19441 11237 19475 11271
rect 20913 11237 20947 11271
rect 21189 11237 21223 11271
rect 18061 11169 18095 11203
rect 23857 11169 23891 11203
rect 15669 11101 15703 11135
rect 16313 11101 16347 11135
rect 16957 11101 16991 11135
rect 17601 11101 17635 11135
rect 18889 11101 18923 11135
rect 20453 11101 20487 11135
rect 21373 11101 21407 11135
rect 21649 11101 21683 11135
rect 22201 11101 22235 11135
rect 22661 11101 22695 11135
rect 24777 11101 24811 11135
rect 19717 11033 19751 11067
rect 19993 11033 20027 11067
rect 20177 11033 20211 11067
rect 20729 11033 20763 11067
rect 24593 10965 24627 10999
rect 15761 10761 15795 10795
rect 16405 10761 16439 10795
rect 17049 10761 17083 10795
rect 18705 10761 18739 10795
rect 17417 10693 17451 10727
rect 23305 10693 23339 10727
rect 18245 10625 18279 10659
rect 18889 10625 18923 10659
rect 19533 10625 19567 10659
rect 20177 10625 20211 10659
rect 20821 10625 20855 10659
rect 21465 10625 21499 10659
rect 22109 10625 22143 10659
rect 23949 10625 23983 10659
rect 24685 10557 24719 10591
rect 18061 10489 18095 10523
rect 19349 10489 19383 10523
rect 19993 10489 20027 10523
rect 20637 10421 20671 10455
rect 21281 10421 21315 10455
rect 17785 10217 17819 10251
rect 19441 10217 19475 10251
rect 20729 10217 20763 10251
rect 21636 10217 21670 10251
rect 24593 10217 24627 10251
rect 23121 10149 23155 10183
rect 18061 10081 18095 10115
rect 21373 10081 21407 10115
rect 25145 10081 25179 10115
rect 18337 10013 18371 10047
rect 19625 10013 19659 10047
rect 20913 10013 20947 10047
rect 24041 10013 24075 10047
rect 25053 10013 25087 10047
rect 24961 9945 24995 9979
rect 20085 9877 20119 9911
rect 23857 9877 23891 9911
rect 21649 9673 21683 9707
rect 23305 9605 23339 9639
rect 18245 9537 18279 9571
rect 18889 9537 18923 9571
rect 19533 9537 19567 9571
rect 20177 9537 20211 9571
rect 20913 9537 20947 9571
rect 21281 9537 21315 9571
rect 22109 9537 22143 9571
rect 23949 9537 23983 9571
rect 21373 9469 21407 9503
rect 24777 9469 24811 9503
rect 18705 9401 18739 9435
rect 19349 9401 19383 9435
rect 20729 9401 20763 9435
rect 18061 9333 18095 9367
rect 19993 9333 20027 9367
rect 11805 9129 11839 9163
rect 24777 9129 24811 9163
rect 19073 9061 19107 9095
rect 21281 9061 21315 9095
rect 10057 8993 10091 9027
rect 19441 8993 19475 9027
rect 23857 8993 23891 9027
rect 19717 8925 19751 8959
rect 21465 8925 21499 8959
rect 22109 8925 22143 8959
rect 22661 8925 22695 8959
rect 10333 8857 10367 8891
rect 12081 8857 12115 8891
rect 24685 8857 24719 8891
rect 21925 8789 21959 8823
rect 19441 8585 19475 8619
rect 21649 8585 21683 8619
rect 19625 8449 19659 8483
rect 20269 8449 20303 8483
rect 20913 8449 20947 8483
rect 21281 8449 21315 8483
rect 22293 8449 22327 8483
rect 23949 8449 23983 8483
rect 23305 8381 23339 8415
rect 24777 8381 24811 8415
rect 20085 8313 20119 8347
rect 20729 8313 20763 8347
rect 21373 8041 21407 8075
rect 22017 7973 22051 8007
rect 23857 7905 23891 7939
rect 20913 7837 20947 7871
rect 21557 7837 21591 7871
rect 22201 7837 22235 7871
rect 22845 7837 22879 7871
rect 24869 7837 24903 7871
rect 20729 7701 20763 7735
rect 24685 7701 24719 7735
rect 21281 7497 21315 7531
rect 23305 7429 23339 7463
rect 25145 7429 25179 7463
rect 20821 7361 20855 7395
rect 21465 7361 21499 7395
rect 22293 7361 22327 7395
rect 23949 7361 23983 7395
rect 20637 7225 20671 7259
rect 23857 6817 23891 6851
rect 21557 6749 21591 6783
rect 22661 6749 22695 6783
rect 24685 6749 24719 6783
rect 24869 6681 24903 6715
rect 21373 6613 21407 6647
rect 22017 6613 22051 6647
rect 23305 6341 23339 6375
rect 22293 6273 22327 6307
rect 24133 6273 24167 6307
rect 24777 6205 24811 6239
rect 22017 5865 22051 5899
rect 21373 5797 21407 5831
rect 21557 5661 21591 5695
rect 22201 5661 22235 5695
rect 22845 5661 22879 5695
rect 24869 5661 24903 5695
rect 23857 5593 23891 5627
rect 24685 5525 24719 5559
rect 22293 5185 22327 5219
rect 23949 5185 23983 5219
rect 23305 5117 23339 5151
rect 24685 5117 24719 5151
rect 22385 4777 22419 4811
rect 22661 4573 22695 4607
rect 24869 4573 24903 4607
rect 23857 4505 23891 4539
rect 24685 4437 24719 4471
rect 20269 4097 20303 4131
rect 22293 4097 22327 4131
rect 23949 4097 23983 4131
rect 21281 4029 21315 4063
rect 23305 4029 23339 4063
rect 24777 4029 24811 4063
rect 20821 3485 20855 3519
rect 22845 3485 22879 3519
rect 24777 3485 24811 3519
rect 22017 3417 22051 3451
rect 23857 3417 23891 3451
rect 24593 3349 24627 3383
rect 23305 3077 23339 3111
rect 25145 3077 25179 3111
rect 18429 3009 18463 3043
rect 20085 3009 20119 3043
rect 22293 3009 22327 3043
rect 24133 3009 24167 3043
rect 19441 2941 19475 2975
rect 21281 2941 21315 2975
rect 6837 2601 6871 2635
rect 7021 2397 7055 2431
rect 7297 2397 7331 2431
rect 20269 2397 20303 2431
rect 22845 2397 22879 2431
rect 21281 2329 21315 2363
rect 23857 2329 23891 2363
<< metal1 >>
rect 3050 26392 3056 26444
rect 3108 26432 3114 26444
rect 3326 26432 3332 26444
rect 3108 26404 3332 26432
rect 3108 26392 3114 26404
rect 3326 26392 3332 26404
rect 3384 26392 3390 26444
rect 5442 26324 5448 26376
rect 5500 26364 5506 26376
rect 21266 26364 21272 26376
rect 5500 26336 21272 26364
rect 5500 26324 5506 26336
rect 21266 26324 21272 26336
rect 21324 26324 21330 26376
rect 4890 26256 4896 26308
rect 4948 26296 4954 26308
rect 20162 26296 20168 26308
rect 4948 26268 20168 26296
rect 4948 26256 4954 26268
rect 20162 26256 20168 26268
rect 20220 26256 20226 26308
rect 5994 25032 6000 25084
rect 6052 25072 6058 25084
rect 13722 25072 13728 25084
rect 6052 25044 13728 25072
rect 6052 25032 6058 25044
rect 13722 25032 13728 25044
rect 13780 25032 13786 25084
rect 9122 24964 9128 25016
rect 9180 25004 9186 25016
rect 20346 25004 20352 25016
rect 9180 24976 20352 25004
rect 9180 24964 9186 24976
rect 20346 24964 20352 24976
rect 20404 24964 20410 25016
rect 1946 24896 1952 24948
rect 2004 24936 2010 24948
rect 16022 24936 16028 24948
rect 2004 24908 16028 24936
rect 2004 24896 2010 24908
rect 16022 24896 16028 24908
rect 16080 24896 16086 24948
rect 6730 24828 6736 24880
rect 6788 24868 6794 24880
rect 26142 24868 26148 24880
rect 6788 24840 26148 24868
rect 6788 24828 6794 24840
rect 26142 24828 26148 24840
rect 26200 24828 26206 24880
rect 14090 24692 14096 24744
rect 14148 24732 14154 24744
rect 23382 24732 23388 24744
rect 14148 24704 23388 24732
rect 14148 24692 14154 24704
rect 23382 24692 23388 24704
rect 23440 24692 23446 24744
rect 16850 24624 16856 24676
rect 16908 24664 16914 24676
rect 24854 24664 24860 24676
rect 16908 24636 24860 24664
rect 16908 24624 16914 24636
rect 24854 24624 24860 24636
rect 24912 24624 24918 24676
rect 4798 24556 4804 24608
rect 4856 24596 4862 24608
rect 12618 24596 12624 24608
rect 4856 24568 12624 24596
rect 4856 24556 4862 24568
rect 12618 24556 12624 24568
rect 12676 24556 12682 24608
rect 16942 24556 16948 24608
rect 17000 24596 17006 24608
rect 24946 24596 24952 24608
rect 17000 24568 24952 24596
rect 17000 24556 17006 24568
rect 24946 24556 24952 24568
rect 25004 24556 25010 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 6546 24352 6552 24404
rect 6604 24352 6610 24404
rect 6638 24352 6644 24404
rect 6696 24392 6702 24404
rect 15013 24395 15071 24401
rect 15013 24392 15025 24395
rect 6696 24364 15025 24392
rect 6696 24352 6702 24364
rect 15013 24361 15025 24364
rect 15059 24361 15071 24395
rect 15013 24355 15071 24361
rect 16942 24352 16948 24404
rect 17000 24352 17006 24404
rect 19150 24392 19156 24404
rect 17512 24364 19156 24392
rect 4982 24284 4988 24336
rect 5040 24324 5046 24336
rect 5040 24296 7236 24324
rect 5040 24284 5046 24296
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 6178 24256 6184 24268
rect 3283 24228 6184 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 6178 24216 6184 24228
rect 6236 24216 6242 24268
rect 2225 24191 2283 24197
rect 2225 24157 2237 24191
rect 2271 24188 2283 24191
rect 3878 24188 3884 24200
rect 2271 24160 3884 24188
rect 2271 24157 2283 24160
rect 2225 24151 2283 24157
rect 3878 24148 3884 24160
rect 3936 24148 3942 24200
rect 4154 24148 4160 24200
rect 4212 24148 4218 24200
rect 4801 24191 4859 24197
rect 4801 24157 4813 24191
rect 4847 24188 4859 24191
rect 6638 24188 6644 24200
rect 4847 24160 6644 24188
rect 4847 24157 4859 24160
rect 4801 24151 4859 24157
rect 6638 24148 6644 24160
rect 6696 24148 6702 24200
rect 6733 24191 6791 24197
rect 6733 24157 6745 24191
rect 6779 24188 6791 24191
rect 7006 24188 7012 24200
rect 6779 24160 7012 24188
rect 6779 24157 6791 24160
rect 6733 24151 6791 24157
rect 7006 24148 7012 24160
rect 7064 24148 7070 24200
rect 7208 24197 7236 24296
rect 9122 24284 9128 24336
rect 9180 24284 9186 24336
rect 11698 24284 11704 24336
rect 11756 24284 11762 24336
rect 12342 24284 12348 24336
rect 12400 24324 12406 24336
rect 15565 24327 15623 24333
rect 12400 24296 12848 24324
rect 12400 24284 12406 24296
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9674 24256 9680 24268
rect 8251 24228 9680 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 10965 24259 11023 24265
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 11238 24256 11244 24268
rect 11011 24228 11244 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 11238 24216 11244 24228
rect 11296 24216 11302 24268
rect 12820 24265 12848 24296
rect 15565 24293 15577 24327
rect 15611 24324 15623 24327
rect 16390 24324 16396 24336
rect 15611 24296 16396 24324
rect 15611 24293 15623 24296
rect 15565 24287 15623 24293
rect 16390 24284 16396 24296
rect 16448 24284 16454 24336
rect 12805 24259 12863 24265
rect 11900 24228 12756 24256
rect 7193 24191 7251 24197
rect 7193 24157 7205 24191
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24157 9367 24191
rect 9309 24151 9367 24157
rect 5813 24123 5871 24129
rect 5813 24089 5825 24123
rect 5859 24120 5871 24123
rect 8662 24120 8668 24132
rect 5859 24092 8668 24120
rect 5859 24089 5871 24092
rect 5813 24083 5871 24089
rect 8662 24080 8668 24092
rect 8720 24080 8726 24132
rect 9324 24120 9352 24151
rect 9490 24148 9496 24200
rect 9548 24188 9554 24200
rect 11900 24197 11928 24228
rect 9769 24191 9827 24197
rect 9769 24188 9781 24191
rect 9548 24160 9781 24188
rect 9548 24148 9554 24160
rect 9769 24157 9781 24160
rect 9815 24157 9827 24191
rect 9769 24151 9827 24157
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24157 11943 24191
rect 11885 24151 11943 24157
rect 12434 24148 12440 24200
rect 12492 24148 12498 24200
rect 12728 24188 12756 24228
rect 12805 24225 12817 24259
rect 12851 24225 12863 24259
rect 12805 24219 12863 24225
rect 16022 24216 16028 24268
rect 16080 24216 16086 24268
rect 16209 24259 16267 24265
rect 16209 24225 16221 24259
rect 16255 24256 16267 24259
rect 17512 24256 17540 24364
rect 19150 24352 19156 24364
rect 19208 24352 19214 24404
rect 21913 24395 21971 24401
rect 21913 24361 21925 24395
rect 21959 24392 21971 24395
rect 22002 24392 22008 24404
rect 21959 24364 22008 24392
rect 21959 24361 21971 24364
rect 21913 24355 21971 24361
rect 22002 24352 22008 24364
rect 22060 24352 22066 24404
rect 24302 24392 24308 24404
rect 22388 24364 24308 24392
rect 18046 24324 18052 24336
rect 17604 24296 18052 24324
rect 17604 24265 17632 24296
rect 18046 24284 18052 24296
rect 18104 24284 18110 24336
rect 18141 24327 18199 24333
rect 18141 24293 18153 24327
rect 18187 24293 18199 24327
rect 18141 24287 18199 24293
rect 16255 24228 17540 24256
rect 17589 24259 17647 24265
rect 16255 24225 16267 24228
rect 16209 24219 16267 24225
rect 17589 24225 17601 24259
rect 17635 24225 17647 24259
rect 17589 24219 17647 24225
rect 17954 24216 17960 24268
rect 18012 24256 18018 24268
rect 18156 24256 18184 24287
rect 18230 24284 18236 24336
rect 18288 24324 18294 24336
rect 21726 24324 21732 24336
rect 18288 24296 21732 24324
rect 18288 24284 18294 24296
rect 21726 24284 21732 24296
rect 21784 24284 21790 24336
rect 18012 24228 18184 24256
rect 18012 24216 18018 24228
rect 18782 24216 18788 24268
rect 18840 24216 18846 24268
rect 22388 24256 22416 24364
rect 24302 24352 24308 24364
rect 24360 24352 24366 24404
rect 24394 24352 24400 24404
rect 24452 24352 24458 24404
rect 20272 24228 22416 24256
rect 15102 24188 15108 24200
rect 12728 24160 15108 24188
rect 15102 24148 15108 24160
rect 15160 24148 15166 24200
rect 20272 24197 20300 24228
rect 23198 24216 23204 24268
rect 23256 24256 23262 24268
rect 25133 24259 25191 24265
rect 25133 24256 25145 24259
rect 23256 24228 25145 24256
rect 23256 24216 23262 24228
rect 25133 24225 25145 24228
rect 25179 24225 25191 24259
rect 25133 24219 25191 24225
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24188 15991 24191
rect 20257 24191 20315 24197
rect 15979 24160 20208 24188
rect 15979 24157 15991 24160
rect 15933 24151 15991 24157
rect 12802 24120 12808 24132
rect 9324 24092 12808 24120
rect 12802 24080 12808 24092
rect 12860 24120 12866 24132
rect 14550 24120 14556 24132
rect 12860 24092 14556 24120
rect 12860 24080 12866 24092
rect 14550 24080 14556 24092
rect 14608 24080 14614 24132
rect 14921 24123 14979 24129
rect 14921 24089 14933 24123
rect 14967 24089 14979 24123
rect 14921 24083 14979 24089
rect 3973 24055 4031 24061
rect 3973 24021 3985 24055
rect 4019 24052 4031 24055
rect 6454 24052 6460 24064
rect 4019 24024 6460 24052
rect 4019 24021 4031 24024
rect 3973 24015 4031 24021
rect 6454 24012 6460 24024
rect 6512 24012 6518 24064
rect 10226 24012 10232 24064
rect 10284 24052 10290 24064
rect 14936 24052 14964 24083
rect 15010 24080 15016 24132
rect 15068 24120 15074 24132
rect 19429 24123 19487 24129
rect 19429 24120 19441 24123
rect 15068 24092 19441 24120
rect 15068 24080 15074 24092
rect 19429 24089 19441 24092
rect 19475 24089 19487 24123
rect 20180 24120 20208 24160
rect 20257 24157 20269 24191
rect 20303 24157 20315 24191
rect 20257 24151 20315 24157
rect 20806 24148 20812 24200
rect 20864 24188 20870 24200
rect 20993 24191 21051 24197
rect 20993 24188 21005 24191
rect 20864 24160 21005 24188
rect 20864 24148 20870 24160
rect 20993 24157 21005 24160
rect 21039 24157 21051 24191
rect 20993 24151 21051 24157
rect 22278 24148 22284 24200
rect 22336 24148 22342 24200
rect 24394 24148 24400 24200
rect 24452 24188 24458 24200
rect 24949 24191 25007 24197
rect 24949 24188 24961 24191
rect 24452 24160 24961 24188
rect 24452 24148 24458 24160
rect 24949 24157 24961 24160
rect 24995 24157 25007 24191
rect 24949 24151 25007 24157
rect 20898 24120 20904 24132
rect 20180 24092 20904 24120
rect 19429 24083 19487 24089
rect 20898 24080 20904 24092
rect 20956 24080 20962 24132
rect 22557 24123 22615 24129
rect 22557 24089 22569 24123
rect 22603 24120 22615 24123
rect 22646 24120 22652 24132
rect 22603 24092 22652 24120
rect 22603 24089 22615 24092
rect 22557 24083 22615 24089
rect 22646 24080 22652 24092
rect 22704 24080 22710 24132
rect 23934 24120 23940 24132
rect 23782 24092 23940 24120
rect 23934 24080 23940 24092
rect 23992 24080 23998 24132
rect 10284 24024 14964 24052
rect 10284 24012 10290 24024
rect 16942 24012 16948 24064
rect 17000 24052 17006 24064
rect 17313 24055 17371 24061
rect 17313 24052 17325 24055
rect 17000 24024 17325 24052
rect 17000 24012 17006 24024
rect 17313 24021 17325 24024
rect 17359 24021 17371 24055
rect 17313 24015 17371 24021
rect 17402 24012 17408 24064
rect 17460 24012 17466 24064
rect 17678 24012 17684 24064
rect 17736 24052 17742 24064
rect 18509 24055 18567 24061
rect 18509 24052 18521 24055
rect 17736 24024 18521 24052
rect 17736 24012 17742 24024
rect 18509 24021 18521 24024
rect 18555 24021 18567 24055
rect 18509 24015 18567 24021
rect 18601 24055 18659 24061
rect 18601 24021 18613 24055
rect 18647 24052 18659 24055
rect 19242 24052 19248 24064
rect 18647 24024 19248 24052
rect 18647 24021 18659 24024
rect 18601 24015 18659 24021
rect 19242 24012 19248 24024
rect 19300 24012 19306 24064
rect 19794 24012 19800 24064
rect 19852 24052 19858 24064
rect 23198 24052 23204 24064
rect 19852 24024 23204 24052
rect 19852 24012 19858 24024
rect 23198 24012 23204 24024
rect 23256 24012 23262 24064
rect 23566 24012 23572 24064
rect 23624 24052 23630 24064
rect 24029 24055 24087 24061
rect 24029 24052 24041 24055
rect 23624 24024 24041 24052
rect 23624 24012 23630 24024
rect 24029 24021 24041 24024
rect 24075 24021 24087 24055
rect 24029 24015 24087 24021
rect 24486 24012 24492 24064
rect 24544 24052 24550 24064
rect 24581 24055 24639 24061
rect 24581 24052 24593 24055
rect 24544 24024 24593 24052
rect 24544 24012 24550 24024
rect 24581 24021 24593 24024
rect 24627 24021 24639 24055
rect 24581 24015 24639 24021
rect 25041 24055 25099 24061
rect 25041 24021 25053 24055
rect 25087 24052 25099 24055
rect 25406 24052 25412 24064
rect 25087 24024 25412 24052
rect 25087 24021 25099 24024
rect 25041 24015 25099 24021
rect 25406 24012 25412 24024
rect 25464 24012 25470 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 2976 23820 12434 23848
rect 1302 23672 1308 23724
rect 1360 23712 1366 23724
rect 2976 23721 3004 23820
rect 3973 23783 4031 23789
rect 3973 23749 3985 23783
rect 4019 23780 4031 23783
rect 5166 23780 5172 23792
rect 4019 23752 5172 23780
rect 4019 23749 4031 23752
rect 3973 23743 4031 23749
rect 5166 23740 5172 23752
rect 5224 23740 5230 23792
rect 5813 23783 5871 23789
rect 5813 23749 5825 23783
rect 5859 23780 5871 23783
rect 7558 23780 7564 23792
rect 5859 23752 7564 23780
rect 5859 23749 5871 23752
rect 5813 23743 5871 23749
rect 7558 23740 7564 23752
rect 7616 23740 7622 23792
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 10134 23780 10140 23792
rect 9171 23752 10140 23780
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 10134 23740 10140 23752
rect 10192 23740 10198 23792
rect 10870 23740 10876 23792
rect 10928 23740 10934 23792
rect 12406 23780 12434 23820
rect 13722 23808 13728 23860
rect 13780 23848 13786 23860
rect 14093 23851 14151 23857
rect 14093 23848 14105 23851
rect 13780 23820 14105 23848
rect 13780 23808 13786 23820
rect 14093 23817 14105 23820
rect 14139 23817 14151 23851
rect 14093 23811 14151 23817
rect 14461 23851 14519 23857
rect 14461 23817 14473 23851
rect 14507 23848 14519 23851
rect 15010 23848 15016 23860
rect 14507 23820 15016 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 15010 23808 15016 23820
rect 15068 23808 15074 23860
rect 15378 23808 15384 23860
rect 15436 23848 15442 23860
rect 17678 23848 17684 23860
rect 15436 23820 17684 23848
rect 15436 23808 15442 23820
rect 17678 23808 17684 23820
rect 17736 23808 17742 23860
rect 23566 23848 23572 23860
rect 17972 23820 21956 23848
rect 16025 23783 16083 23789
rect 16025 23780 16037 23783
rect 12406 23752 16037 23780
rect 16025 23749 16037 23752
rect 16071 23749 16083 23783
rect 16025 23743 16083 23749
rect 17221 23783 17279 23789
rect 17221 23749 17233 23783
rect 17267 23780 17279 23783
rect 17310 23780 17316 23792
rect 17267 23752 17316 23780
rect 17267 23749 17279 23752
rect 17221 23743 17279 23749
rect 17310 23740 17316 23752
rect 17368 23740 17374 23792
rect 1673 23715 1731 23721
rect 1673 23712 1685 23715
rect 1360 23684 1685 23712
rect 1360 23672 1366 23684
rect 1673 23681 1685 23684
rect 1719 23712 1731 23715
rect 2133 23715 2191 23721
rect 2133 23712 2145 23715
rect 1719 23684 2145 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 2133 23681 2145 23684
rect 2179 23681 2191 23715
rect 2133 23675 2191 23681
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23681 3019 23715
rect 2961 23675 3019 23681
rect 4798 23672 4804 23724
rect 4856 23672 4862 23724
rect 5442 23672 5448 23724
rect 5500 23712 5506 23724
rect 7929 23715 7987 23721
rect 7929 23712 7941 23715
rect 5500 23684 7941 23712
rect 5500 23672 5506 23684
rect 7929 23681 7941 23684
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 9769 23715 9827 23721
rect 9769 23681 9781 23715
rect 9815 23681 9827 23715
rect 12069 23715 12127 23721
rect 12069 23712 12081 23715
rect 9769 23675 9827 23681
rect 9876 23684 12081 23712
rect 1857 23647 1915 23653
rect 1857 23613 1869 23647
rect 1903 23644 1915 23647
rect 6549 23647 6607 23653
rect 1903 23616 6316 23644
rect 1903 23613 1915 23616
rect 1857 23607 1915 23613
rect 6288 23576 6316 23616
rect 6549 23613 6561 23647
rect 6595 23644 6607 23647
rect 6638 23644 6644 23656
rect 6595 23616 6644 23644
rect 6595 23613 6607 23616
rect 6549 23607 6607 23613
rect 6638 23604 6644 23616
rect 6696 23604 6702 23656
rect 6730 23604 6736 23656
rect 6788 23644 6794 23656
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 6788 23616 6837 23644
rect 6788 23604 6794 23616
rect 6825 23613 6837 23616
rect 6871 23613 6883 23647
rect 6825 23607 6883 23613
rect 6914 23604 6920 23656
rect 6972 23644 6978 23656
rect 6972 23616 7696 23644
rect 6972 23604 6978 23616
rect 7098 23576 7104 23588
rect 6288 23548 7104 23576
rect 7098 23536 7104 23548
rect 7156 23536 7162 23588
rect 7668 23576 7696 23616
rect 7834 23604 7840 23656
rect 7892 23644 7898 23656
rect 9784 23644 9812 23675
rect 7892 23616 9812 23644
rect 7892 23604 7898 23616
rect 9876 23576 9904 23684
rect 12069 23681 12081 23684
rect 12115 23681 12127 23715
rect 12069 23675 12127 23681
rect 15841 23715 15899 23721
rect 15841 23681 15853 23715
rect 15887 23712 15899 23715
rect 16114 23712 16120 23724
rect 15887 23684 16120 23712
rect 15887 23681 15899 23684
rect 15841 23675 15899 23681
rect 16114 23672 16120 23684
rect 16172 23672 16178 23724
rect 17126 23672 17132 23724
rect 17184 23712 17190 23724
rect 17862 23712 17868 23724
rect 17184 23684 17868 23712
rect 17184 23672 17190 23684
rect 17862 23672 17868 23684
rect 17920 23672 17926 23724
rect 11974 23604 11980 23656
rect 12032 23644 12038 23656
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 12032 23616 12541 23644
rect 12032 23604 12038 23616
rect 12529 23613 12541 23616
rect 12575 23613 12587 23647
rect 12529 23607 12587 23613
rect 14553 23647 14611 23653
rect 14553 23613 14565 23647
rect 14599 23613 14611 23647
rect 14553 23607 14611 23613
rect 7668 23548 9904 23576
rect 11609 23579 11667 23585
rect 11609 23545 11621 23579
rect 11655 23576 11667 23579
rect 12802 23576 12808 23588
rect 11655 23548 12808 23576
rect 11655 23545 11667 23548
rect 11609 23539 11667 23545
rect 12802 23536 12808 23548
rect 12860 23536 12866 23588
rect 14568 23576 14596 23607
rect 14734 23604 14740 23656
rect 14792 23604 14798 23656
rect 14918 23604 14924 23656
rect 14976 23644 14982 23656
rect 17313 23647 17371 23653
rect 17313 23644 17325 23647
rect 14976 23616 17325 23644
rect 14976 23604 14982 23616
rect 17313 23613 17325 23616
rect 17359 23613 17371 23647
rect 17313 23607 17371 23613
rect 17497 23647 17555 23653
rect 17497 23613 17509 23647
rect 17543 23644 17555 23647
rect 17972 23644 18000 23820
rect 20073 23783 20131 23789
rect 20073 23780 20085 23783
rect 19550 23752 20085 23780
rect 20073 23749 20085 23752
rect 20119 23780 20131 23783
rect 20257 23783 20315 23789
rect 20257 23780 20269 23783
rect 20119 23752 20269 23780
rect 20119 23749 20131 23752
rect 20073 23743 20131 23749
rect 20257 23749 20269 23752
rect 20303 23780 20315 23783
rect 20806 23780 20812 23792
rect 20303 23752 20812 23780
rect 20303 23749 20315 23752
rect 20257 23743 20315 23749
rect 20806 23740 20812 23752
rect 20864 23780 20870 23792
rect 21821 23783 21879 23789
rect 21821 23780 21833 23783
rect 20864 23752 21833 23780
rect 20864 23740 20870 23752
rect 21821 23749 21833 23752
rect 21867 23749 21879 23783
rect 21928 23780 21956 23820
rect 22066 23820 23572 23848
rect 22066 23780 22094 23820
rect 23566 23808 23572 23820
rect 23624 23808 23630 23860
rect 24302 23808 24308 23860
rect 24360 23808 24366 23860
rect 23934 23780 23940 23792
rect 21928 23752 22094 23780
rect 23782 23752 23940 23780
rect 21821 23743 21879 23749
rect 23934 23740 23940 23752
rect 23992 23780 23998 23792
rect 24578 23780 24584 23792
rect 23992 23752 24584 23780
rect 23992 23740 23998 23752
rect 24578 23740 24584 23752
rect 24636 23740 24642 23792
rect 24762 23740 24768 23792
rect 24820 23780 24826 23792
rect 25133 23783 25191 23789
rect 25133 23780 25145 23783
rect 24820 23752 25145 23780
rect 24820 23740 24826 23752
rect 25133 23749 25145 23752
rect 25179 23749 25191 23783
rect 25133 23743 25191 23749
rect 18046 23672 18052 23724
rect 18104 23672 18110 23724
rect 20625 23715 20683 23721
rect 20625 23681 20637 23715
rect 20671 23712 20683 23715
rect 22002 23712 22008 23724
rect 20671 23684 22008 23712
rect 20671 23681 20683 23684
rect 20625 23675 20683 23681
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 17543 23616 18000 23644
rect 18325 23647 18383 23653
rect 17543 23613 17555 23616
rect 17497 23607 17555 23613
rect 18325 23613 18337 23647
rect 18371 23644 18383 23647
rect 18782 23644 18788 23656
rect 18371 23616 18788 23644
rect 18371 23613 18383 23616
rect 18325 23607 18383 23613
rect 18782 23604 18788 23616
rect 18840 23644 18846 23656
rect 20714 23644 20720 23656
rect 18840 23616 20720 23644
rect 18840 23604 18846 23616
rect 20714 23604 20720 23616
rect 20772 23604 20778 23656
rect 20898 23604 20904 23656
rect 20956 23604 20962 23656
rect 22278 23604 22284 23656
rect 22336 23604 22342 23656
rect 22554 23644 22560 23656
rect 22388 23616 22560 23644
rect 17770 23576 17776 23588
rect 14568 23548 17776 23576
rect 17770 23536 17776 23548
rect 17828 23536 17834 23588
rect 20254 23576 20260 23588
rect 19720 23548 20260 23576
rect 2501 23511 2559 23517
rect 2501 23477 2513 23511
rect 2547 23508 2559 23511
rect 7006 23508 7012 23520
rect 2547 23480 7012 23508
rect 2547 23477 2559 23480
rect 2501 23471 2559 23477
rect 7006 23468 7012 23480
rect 7064 23508 7070 23520
rect 13630 23508 13636 23520
rect 7064 23480 13636 23508
rect 7064 23468 7070 23480
rect 13630 23468 13636 23480
rect 13688 23468 13694 23520
rect 15838 23468 15844 23520
rect 15896 23508 15902 23520
rect 16393 23511 16451 23517
rect 16393 23508 16405 23511
rect 15896 23480 16405 23508
rect 15896 23468 15902 23480
rect 16393 23477 16405 23480
rect 16439 23477 16451 23511
rect 16393 23471 16451 23477
rect 16850 23468 16856 23520
rect 16908 23468 16914 23520
rect 16942 23468 16948 23520
rect 17000 23508 17006 23520
rect 19720 23508 19748 23548
rect 20254 23536 20260 23548
rect 20312 23536 20318 23588
rect 21726 23536 21732 23588
rect 21784 23576 21790 23588
rect 22388 23576 22416 23616
rect 22554 23604 22560 23616
rect 22612 23604 22618 23656
rect 22646 23604 22652 23656
rect 22704 23644 22710 23656
rect 24029 23647 24087 23653
rect 24029 23644 24041 23647
rect 22704 23616 24041 23644
rect 22704 23604 22710 23616
rect 24029 23613 24041 23616
rect 24075 23644 24087 23647
rect 25498 23644 25504 23656
rect 24075 23616 25504 23644
rect 24075 23613 24087 23616
rect 24029 23607 24087 23613
rect 25498 23604 25504 23616
rect 25556 23604 25562 23656
rect 25317 23579 25375 23585
rect 25317 23576 25329 23579
rect 21784 23548 22416 23576
rect 23676 23548 25329 23576
rect 21784 23536 21790 23548
rect 17000 23480 19748 23508
rect 17000 23468 17006 23480
rect 19794 23468 19800 23520
rect 19852 23468 19858 23520
rect 21634 23468 21640 23520
rect 21692 23508 21698 23520
rect 23676 23508 23704 23548
rect 25317 23545 25329 23548
rect 25363 23545 25375 23579
rect 25317 23539 25375 23545
rect 21692 23480 23704 23508
rect 21692 23468 21698 23480
rect 24578 23468 24584 23520
rect 24636 23468 24642 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 6638 23264 6644 23316
rect 6696 23304 6702 23316
rect 7374 23304 7380 23316
rect 6696 23276 7380 23304
rect 6696 23264 6702 23276
rect 7374 23264 7380 23276
rect 7432 23304 7438 23316
rect 11790 23304 11796 23316
rect 7432 23276 11796 23304
rect 7432 23264 7438 23276
rect 11790 23264 11796 23276
rect 11848 23264 11854 23316
rect 11900 23276 13584 23304
rect 4249 23239 4307 23245
rect 4249 23205 4261 23239
rect 4295 23236 4307 23239
rect 7282 23236 7288 23248
rect 4295 23208 7288 23236
rect 4295 23205 4307 23208
rect 4249 23199 4307 23205
rect 7282 23196 7288 23208
rect 7340 23196 7346 23248
rect 7466 23196 7472 23248
rect 7524 23236 7530 23248
rect 11900 23236 11928 23276
rect 7524 23208 9904 23236
rect 7524 23196 7530 23208
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 8386 23168 8392 23180
rect 2832 23140 4016 23168
rect 2832 23128 2838 23140
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23100 2283 23103
rect 2271 23072 2774 23100
rect 2271 23069 2283 23072
rect 2225 23063 2283 23069
rect 2746 22964 2774 23072
rect 3988 23096 4016 23140
rect 5460 23140 8392 23168
rect 5460 23109 5488 23140
rect 8386 23128 8392 23140
rect 8444 23128 8450 23180
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 9272 23140 9536 23168
rect 9272 23128 9278 23140
rect 4065 23103 4123 23109
rect 4065 23096 4077 23103
rect 3988 23069 4077 23096
rect 4111 23069 4123 23103
rect 3988 23068 4123 23069
rect 4065 23063 4123 23068
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23069 5503 23103
rect 5445 23063 5503 23069
rect 5902 23060 5908 23112
rect 5960 23100 5966 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 5960 23072 7205 23100
rect 5960 23060 5966 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 8205 23103 8263 23109
rect 8205 23069 8217 23103
rect 8251 23100 8263 23103
rect 9306 23100 9312 23112
rect 8251 23072 9312 23100
rect 8251 23069 8263 23072
rect 8205 23063 8263 23069
rect 9306 23060 9312 23072
rect 9364 23060 9370 23112
rect 9401 23103 9459 23109
rect 9401 23069 9413 23103
rect 9447 23069 9459 23103
rect 9401 23063 9459 23069
rect 3237 23035 3295 23041
rect 3237 23001 3249 23035
rect 3283 23032 3295 23035
rect 4338 23032 4344 23044
rect 3283 23004 4344 23032
rect 3283 23001 3295 23004
rect 3237 22995 3295 23001
rect 4338 22992 4344 23004
rect 4396 22992 4402 23044
rect 6270 23032 6276 23044
rect 4632 23004 6276 23032
rect 4632 22964 4660 23004
rect 6270 22992 6276 23004
rect 6328 22992 6334 23044
rect 6365 23035 6423 23041
rect 6365 23001 6377 23035
rect 6411 23001 6423 23035
rect 6365 22995 6423 23001
rect 2746 22936 4660 22964
rect 4706 22924 4712 22976
rect 4764 22924 4770 22976
rect 6380 22964 6408 22995
rect 6454 22992 6460 23044
rect 6512 23032 6518 23044
rect 9416 23032 9444 23063
rect 6512 23004 9444 23032
rect 9508 23032 9536 23140
rect 9876 23109 9904 23208
rect 9968 23208 11928 23236
rect 9861 23103 9919 23109
rect 9861 23069 9873 23103
rect 9907 23069 9919 23103
rect 9861 23063 9919 23069
rect 9968 23032 9996 23208
rect 12526 23196 12532 23248
rect 12584 23236 12590 23248
rect 13446 23236 13452 23248
rect 12584 23208 13452 23236
rect 12584 23196 12590 23208
rect 13446 23196 13452 23208
rect 13504 23196 13510 23248
rect 13556 23236 13584 23276
rect 13630 23264 13636 23316
rect 13688 23304 13694 23316
rect 14826 23304 14832 23316
rect 13688 23276 14832 23304
rect 13688 23264 13694 23276
rect 14826 23264 14832 23276
rect 14884 23264 14890 23316
rect 16298 23304 16304 23316
rect 14936 23276 16304 23304
rect 14936 23236 14964 23276
rect 16298 23264 16304 23276
rect 16356 23264 16362 23316
rect 17954 23264 17960 23316
rect 18012 23304 18018 23316
rect 24486 23304 24492 23316
rect 18012 23276 24492 23304
rect 18012 23264 18018 23276
rect 24486 23264 24492 23276
rect 24544 23264 24550 23316
rect 13556 23208 14964 23236
rect 16942 23196 16948 23248
rect 17000 23236 17006 23248
rect 19334 23236 19340 23248
rect 17000 23208 19340 23236
rect 17000 23196 17006 23208
rect 19334 23196 19340 23208
rect 19392 23196 19398 23248
rect 20714 23196 20720 23248
rect 20772 23236 20778 23248
rect 21177 23239 21235 23245
rect 21177 23236 21189 23239
rect 20772 23208 21189 23236
rect 20772 23196 20778 23208
rect 21177 23205 21189 23208
rect 21223 23205 21235 23239
rect 21177 23199 21235 23205
rect 23382 23196 23388 23248
rect 23440 23236 23446 23248
rect 24581 23239 24639 23245
rect 24581 23236 24593 23239
rect 23440 23208 24593 23236
rect 23440 23196 23446 23208
rect 24581 23205 24593 23208
rect 24627 23205 24639 23239
rect 24581 23199 24639 23205
rect 10502 23128 10508 23180
rect 10560 23128 10566 23180
rect 11606 23128 11612 23180
rect 11664 23168 11670 23180
rect 12161 23171 12219 23177
rect 12161 23168 12173 23171
rect 11664 23140 12173 23168
rect 11664 23128 11670 23140
rect 12161 23137 12173 23140
rect 12207 23137 12219 23171
rect 13906 23168 13912 23180
rect 12161 23131 12219 23137
rect 13280 23140 13912 23168
rect 11701 23103 11759 23109
rect 11701 23069 11713 23103
rect 11747 23069 11759 23103
rect 11701 23063 11759 23069
rect 9508 23004 9996 23032
rect 6512 22992 6518 23004
rect 7650 22964 7656 22976
rect 6380 22936 7656 22964
rect 7650 22924 7656 22936
rect 7708 22924 7714 22976
rect 9217 22967 9275 22973
rect 9217 22933 9229 22967
rect 9263 22964 9275 22967
rect 11716 22964 11744 23063
rect 11790 23060 11796 23112
rect 11848 23100 11854 23112
rect 13280 23100 13308 23140
rect 13906 23128 13912 23140
rect 13964 23128 13970 23180
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 17126 23168 17132 23180
rect 15335 23140 17132 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 17126 23128 17132 23140
rect 17184 23128 17190 23180
rect 17402 23128 17408 23180
rect 17460 23168 17466 23180
rect 17681 23171 17739 23177
rect 17681 23168 17693 23171
rect 17460 23140 17693 23168
rect 17460 23128 17466 23140
rect 17681 23137 17693 23140
rect 17727 23137 17739 23171
rect 17681 23131 17739 23137
rect 17862 23128 17868 23180
rect 17920 23168 17926 23180
rect 18414 23168 18420 23180
rect 17920 23140 18420 23168
rect 17920 23128 17926 23140
rect 18414 23128 18420 23140
rect 18472 23128 18478 23180
rect 18690 23128 18696 23180
rect 18748 23168 18754 23180
rect 20990 23168 20996 23180
rect 18748 23140 20996 23168
rect 18748 23128 18754 23140
rect 20990 23128 20996 23140
rect 21048 23128 21054 23180
rect 21637 23171 21695 23177
rect 21637 23137 21649 23171
rect 21683 23168 21695 23171
rect 22278 23168 22284 23180
rect 21683 23140 22284 23168
rect 21683 23137 21695 23140
rect 21637 23131 21695 23137
rect 22278 23128 22284 23140
rect 22336 23168 22342 23180
rect 23290 23168 23296 23180
rect 22336 23140 23296 23168
rect 22336 23128 22342 23140
rect 23290 23128 23296 23140
rect 23348 23128 23354 23180
rect 25133 23171 25191 23177
rect 25133 23137 25145 23171
rect 25179 23137 25191 23171
rect 25133 23131 25191 23137
rect 11848 23072 13308 23100
rect 11848 23060 11854 23072
rect 13722 23060 13728 23112
rect 13780 23060 13786 23112
rect 14274 23060 14280 23112
rect 14332 23100 14338 23112
rect 15013 23103 15071 23109
rect 15013 23100 15025 23103
rect 14332 23072 15025 23100
rect 14332 23060 14338 23072
rect 15013 23069 15025 23072
rect 15059 23069 15071 23103
rect 15013 23063 15071 23069
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23096 17647 23103
rect 17954 23100 17960 23112
rect 17696 23096 17960 23100
rect 17635 23072 17960 23096
rect 17635 23069 17724 23072
rect 17589 23068 17724 23069
rect 17589 23063 17647 23068
rect 17954 23060 17960 23072
rect 18012 23060 18018 23112
rect 18046 23060 18052 23112
rect 18104 23100 18110 23112
rect 19334 23100 19340 23112
rect 18104 23072 19340 23100
rect 18104 23060 18110 23072
rect 19334 23060 19340 23072
rect 19392 23100 19398 23112
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 19392 23072 19441 23100
rect 19392 23060 19398 23072
rect 19429 23069 19441 23072
rect 19475 23069 19487 23103
rect 19429 23063 19487 23069
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 21266 23100 21272 23112
rect 20864 23072 21272 23100
rect 20864 23060 20870 23072
rect 21266 23060 21272 23072
rect 21324 23060 21330 23112
rect 23198 23060 23204 23112
rect 23256 23100 23262 23112
rect 25148 23100 25176 23131
rect 23256 23072 25176 23100
rect 23256 23060 23262 23072
rect 13446 22992 13452 23044
rect 13504 23032 13510 23044
rect 13504 23004 13952 23032
rect 13504 22992 13510 23004
rect 9263 22936 11744 22964
rect 9263 22933 9275 22936
rect 9217 22927 9275 22933
rect 13538 22924 13544 22976
rect 13596 22924 13602 22976
rect 13924 22964 13952 23004
rect 14366 22992 14372 23044
rect 14424 22992 14430 23044
rect 15838 22992 15844 23044
rect 15896 22992 15902 23044
rect 17126 22992 17132 23044
rect 17184 23032 17190 23044
rect 17402 23032 17408 23044
rect 17184 23004 17408 23032
rect 17184 22992 17190 23004
rect 17402 22992 17408 23004
rect 17460 22992 17466 23044
rect 18506 22992 18512 23044
rect 18564 22992 18570 23044
rect 18598 22992 18604 23044
rect 18656 23032 18662 23044
rect 18693 23035 18751 23041
rect 18693 23032 18705 23035
rect 18656 23004 18705 23032
rect 18656 22992 18662 23004
rect 18693 23001 18705 23004
rect 18739 23001 18751 23035
rect 18693 22995 18751 23001
rect 19702 22992 19708 23044
rect 19760 22992 19766 23044
rect 21913 23035 21971 23041
rect 21913 23001 21925 23035
rect 21959 23032 21971 23035
rect 22002 23032 22008 23044
rect 21959 23004 22008 23032
rect 21959 23001 21971 23004
rect 21913 22995 21971 23001
rect 22002 22992 22008 23004
rect 22060 22992 22066 23044
rect 23658 23032 23664 23044
rect 23138 23004 23664 23032
rect 23658 22992 23664 23004
rect 23716 22992 23722 23044
rect 24489 23035 24547 23041
rect 24489 23001 24501 23035
rect 24535 23032 24547 23035
rect 24535 23004 25084 23032
rect 24535 23001 24547 23004
rect 24489 22995 24547 23001
rect 14461 22967 14519 22973
rect 14461 22964 14473 22967
rect 13924 22936 14473 22964
rect 14461 22933 14473 22936
rect 14507 22933 14519 22967
rect 14461 22927 14519 22933
rect 14642 22924 14648 22976
rect 14700 22964 14706 22976
rect 16666 22964 16672 22976
rect 14700 22936 16672 22964
rect 14700 22924 14706 22936
rect 16666 22924 16672 22936
rect 16724 22964 16730 22976
rect 16761 22967 16819 22973
rect 16761 22964 16773 22967
rect 16724 22936 16773 22964
rect 16724 22924 16730 22936
rect 16761 22933 16773 22936
rect 16807 22933 16819 22967
rect 16761 22927 16819 22933
rect 16850 22924 16856 22976
rect 16908 22964 16914 22976
rect 17221 22967 17279 22973
rect 17221 22964 17233 22967
rect 16908 22936 17233 22964
rect 16908 22924 16914 22936
rect 17221 22933 17233 22936
rect 17267 22933 17279 22967
rect 17221 22927 17279 22933
rect 17862 22924 17868 22976
rect 17920 22964 17926 22976
rect 19794 22964 19800 22976
rect 17920 22936 19800 22964
rect 17920 22924 17926 22936
rect 19794 22924 19800 22936
rect 19852 22924 19858 22976
rect 22554 22924 22560 22976
rect 22612 22964 22618 22976
rect 23385 22967 23443 22973
rect 23385 22964 23397 22967
rect 22612 22936 23397 22964
rect 22612 22924 22618 22936
rect 23385 22933 23397 22936
rect 23431 22933 23443 22967
rect 23385 22927 23443 22933
rect 23845 22967 23903 22973
rect 23845 22933 23857 22967
rect 23891 22964 23903 22967
rect 24026 22964 24032 22976
rect 23891 22936 24032 22964
rect 23891 22933 23903 22936
rect 23845 22927 23903 22933
rect 24026 22924 24032 22936
rect 24084 22924 24090 22976
rect 24762 22924 24768 22976
rect 24820 22964 24826 22976
rect 25056 22973 25084 23004
rect 24949 22967 25007 22973
rect 24949 22964 24961 22967
rect 24820 22936 24961 22964
rect 24820 22924 24826 22936
rect 24949 22933 24961 22936
rect 24995 22933 25007 22967
rect 24949 22927 25007 22933
rect 25041 22967 25099 22973
rect 25041 22933 25053 22967
rect 25087 22964 25099 22967
rect 25958 22964 25964 22976
rect 25087 22936 25964 22964
rect 25087 22933 25099 22936
rect 25041 22927 25099 22933
rect 25958 22924 25964 22936
rect 26016 22924 26022 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 2501 22763 2559 22769
rect 2501 22729 2513 22763
rect 2547 22760 2559 22763
rect 2774 22760 2780 22772
rect 2547 22732 2780 22760
rect 2547 22729 2559 22732
rect 2501 22723 2559 22729
rect 2774 22720 2780 22732
rect 2832 22720 2838 22772
rect 4706 22720 4712 22772
rect 4764 22760 4770 22772
rect 12069 22763 12127 22769
rect 12069 22760 12081 22763
rect 4764 22732 12081 22760
rect 4764 22720 4770 22732
rect 12069 22729 12081 22732
rect 12115 22729 12127 22763
rect 12069 22723 12127 22729
rect 12618 22720 12624 22772
rect 12676 22760 12682 22772
rect 13081 22763 13139 22769
rect 13081 22760 13093 22763
rect 12676 22732 13093 22760
rect 12676 22720 12682 22732
rect 13081 22729 13093 22732
rect 13127 22729 13139 22763
rect 14642 22760 14648 22772
rect 13081 22723 13139 22729
rect 13924 22732 14648 22760
rect 3973 22695 4031 22701
rect 3973 22661 3985 22695
rect 4019 22692 4031 22695
rect 4246 22692 4252 22704
rect 4019 22664 4252 22692
rect 4019 22661 4031 22664
rect 3973 22655 4031 22661
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 5718 22652 5724 22704
rect 5776 22652 5782 22704
rect 7285 22695 7343 22701
rect 7285 22661 7297 22695
rect 7331 22692 7343 22695
rect 7374 22692 7380 22704
rect 7331 22664 7380 22692
rect 7331 22661 7343 22664
rect 7285 22655 7343 22661
rect 7374 22652 7380 22664
rect 7432 22652 7438 22704
rect 8754 22652 8760 22704
rect 8812 22652 8818 22704
rect 10410 22652 10416 22704
rect 10468 22652 10474 22704
rect 11606 22652 11612 22704
rect 11664 22692 11670 22704
rect 13538 22692 13544 22704
rect 11664 22664 13544 22692
rect 11664 22652 11670 22664
rect 13538 22652 13544 22664
rect 13596 22652 13602 22704
rect 13924 22701 13952 22732
rect 14642 22720 14648 22732
rect 14700 22720 14706 22772
rect 14734 22720 14740 22772
rect 14792 22760 14798 22772
rect 15381 22763 15439 22769
rect 15381 22760 15393 22763
rect 14792 22732 15393 22760
rect 14792 22720 14798 22732
rect 15381 22729 15393 22732
rect 15427 22729 15439 22763
rect 15381 22723 15439 22729
rect 15838 22720 15844 22772
rect 15896 22760 15902 22772
rect 16393 22763 16451 22769
rect 16393 22760 16405 22763
rect 15896 22732 16405 22760
rect 15896 22720 15902 22732
rect 16393 22729 16405 22732
rect 16439 22760 16451 22763
rect 16439 22732 17264 22760
rect 16439 22729 16451 22732
rect 16393 22723 16451 22729
rect 13909 22695 13967 22701
rect 13909 22661 13921 22695
rect 13955 22661 13967 22695
rect 15856 22692 15884 22720
rect 15134 22664 15884 22692
rect 17236 22692 17264 22732
rect 18414 22720 18420 22772
rect 18472 22760 18478 22772
rect 18601 22763 18659 22769
rect 18601 22760 18613 22763
rect 18472 22732 18613 22760
rect 18472 22720 18478 22732
rect 18601 22729 18613 22732
rect 18647 22729 18659 22763
rect 18601 22723 18659 22729
rect 19061 22763 19119 22769
rect 19061 22729 19073 22763
rect 19107 22729 19119 22763
rect 19061 22723 19119 22729
rect 17236 22664 17618 22692
rect 13909 22655 13967 22661
rect 1302 22584 1308 22636
rect 1360 22624 1366 22636
rect 1673 22627 1731 22633
rect 1673 22624 1685 22627
rect 1360 22596 1685 22624
rect 1360 22584 1366 22596
rect 1673 22593 1685 22596
rect 1719 22624 1731 22627
rect 2133 22627 2191 22633
rect 2133 22624 2145 22627
rect 1719 22596 2145 22624
rect 1719 22593 1731 22596
rect 1673 22587 1731 22593
rect 2133 22593 2145 22596
rect 2179 22593 2191 22627
rect 2133 22587 2191 22593
rect 2961 22627 3019 22633
rect 2961 22593 2973 22627
rect 3007 22624 3019 22627
rect 3786 22624 3792 22636
rect 3007 22596 3792 22624
rect 3007 22593 3019 22596
rect 2961 22587 3019 22593
rect 3786 22584 3792 22596
rect 3844 22584 3850 22636
rect 4801 22627 4859 22633
rect 4801 22593 4813 22627
rect 4847 22624 4859 22627
rect 4847 22596 5304 22624
rect 4847 22593 4859 22596
rect 4801 22587 4859 22593
rect 1857 22491 1915 22497
rect 1857 22457 1869 22491
rect 1903 22488 1915 22491
rect 5276 22488 5304 22596
rect 6638 22584 6644 22636
rect 6696 22584 6702 22636
rect 7561 22627 7619 22633
rect 7561 22593 7573 22627
rect 7607 22593 7619 22627
rect 7561 22587 7619 22593
rect 12161 22627 12219 22633
rect 12161 22593 12173 22627
rect 12207 22624 12219 22627
rect 12207 22596 12940 22624
rect 12207 22593 12219 22596
rect 12161 22587 12219 22593
rect 5350 22516 5356 22568
rect 5408 22556 5414 22568
rect 7576 22556 7604 22587
rect 5408 22528 7604 22556
rect 5408 22516 5414 22528
rect 9030 22516 9036 22568
rect 9088 22556 9094 22568
rect 9401 22559 9459 22565
rect 9401 22556 9413 22559
rect 9088 22528 9413 22556
rect 9088 22516 9094 22528
rect 9401 22525 9413 22528
rect 9447 22525 9459 22559
rect 9401 22519 9459 22525
rect 9677 22559 9735 22565
rect 9677 22525 9689 22559
rect 9723 22556 9735 22559
rect 12250 22556 12256 22568
rect 9723 22528 12256 22556
rect 9723 22525 9735 22528
rect 9677 22519 9735 22525
rect 12250 22516 12256 22528
rect 12308 22516 12314 22568
rect 12912 22556 12940 22596
rect 12986 22584 12992 22636
rect 13044 22584 13050 22636
rect 13630 22584 13636 22636
rect 13688 22584 13694 22636
rect 15746 22584 15752 22636
rect 15804 22624 15810 22636
rect 15933 22627 15991 22633
rect 15933 22624 15945 22627
rect 15804 22596 15945 22624
rect 15804 22584 15810 22596
rect 15933 22593 15945 22596
rect 15979 22593 15991 22627
rect 15933 22587 15991 22593
rect 16022 22584 16028 22636
rect 16080 22624 16086 22636
rect 16117 22627 16175 22633
rect 16117 22624 16129 22627
rect 16080 22596 16129 22624
rect 16080 22584 16086 22596
rect 16117 22593 16129 22596
rect 16163 22593 16175 22627
rect 16117 22587 16175 22593
rect 16574 22584 16580 22636
rect 16632 22624 16638 22636
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16632 22596 16865 22624
rect 16632 22584 16638 22596
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 17129 22559 17187 22565
rect 17129 22556 17141 22559
rect 12912 22528 15332 22556
rect 11330 22488 11336 22500
rect 1903 22460 2774 22488
rect 5276 22460 6868 22488
rect 1903 22457 1915 22460
rect 1857 22451 1915 22457
rect 2746 22420 2774 22460
rect 4062 22420 4068 22432
rect 2746 22392 4068 22420
rect 4062 22380 4068 22392
rect 4120 22380 4126 22432
rect 4154 22380 4160 22432
rect 4212 22420 4218 22432
rect 6733 22423 6791 22429
rect 6733 22420 6745 22423
rect 4212 22392 6745 22420
rect 4212 22380 4218 22392
rect 6733 22389 6745 22392
rect 6779 22389 6791 22423
rect 6840 22420 6868 22460
rect 10704 22460 11336 22488
rect 10704 22420 10732 22460
rect 11330 22448 11336 22460
rect 11388 22448 11394 22500
rect 11882 22448 11888 22500
rect 11940 22488 11946 22500
rect 12986 22488 12992 22500
rect 11940 22460 12992 22488
rect 11940 22448 11946 22460
rect 12986 22448 12992 22460
rect 13044 22448 13050 22500
rect 6840 22392 10732 22420
rect 6733 22383 6791 22389
rect 11146 22380 11152 22432
rect 11204 22380 11210 22432
rect 11238 22380 11244 22432
rect 11296 22420 11302 22432
rect 11701 22423 11759 22429
rect 11701 22420 11713 22423
rect 11296 22392 11713 22420
rect 11296 22380 11302 22392
rect 11701 22389 11713 22392
rect 11747 22389 11759 22423
rect 11701 22383 11759 22389
rect 13630 22380 13636 22432
rect 13688 22420 13694 22432
rect 14274 22420 14280 22432
rect 13688 22392 14280 22420
rect 13688 22380 13694 22392
rect 14274 22380 14280 22392
rect 14332 22380 14338 22432
rect 15304 22420 15332 22528
rect 16960 22528 17141 22556
rect 16482 22448 16488 22500
rect 16540 22488 16546 22500
rect 16960 22488 16988 22528
rect 17129 22525 17141 22528
rect 17175 22525 17187 22559
rect 17129 22519 17187 22525
rect 17770 22516 17776 22568
rect 17828 22556 17834 22568
rect 19076 22556 19104 22723
rect 19242 22720 19248 22772
rect 19300 22760 19306 22772
rect 20257 22763 20315 22769
rect 20257 22760 20269 22763
rect 19300 22732 20269 22760
rect 19300 22720 19306 22732
rect 20257 22729 20269 22732
rect 20303 22729 20315 22763
rect 20257 22723 20315 22729
rect 20530 22720 20536 22772
rect 20588 22760 20594 22772
rect 20588 22732 20944 22760
rect 20588 22720 20594 22732
rect 19702 22652 19708 22704
rect 19760 22692 19766 22704
rect 20438 22692 20444 22704
rect 19760 22664 20444 22692
rect 19760 22652 19766 22664
rect 20438 22652 20444 22664
rect 20496 22692 20502 22704
rect 20496 22664 20852 22692
rect 20496 22652 20502 22664
rect 19429 22627 19487 22633
rect 19429 22593 19441 22627
rect 19475 22624 19487 22627
rect 19794 22624 19800 22636
rect 19475 22596 19800 22624
rect 19475 22593 19487 22596
rect 19429 22587 19487 22593
rect 19794 22584 19800 22596
rect 19852 22584 19858 22636
rect 20162 22584 20168 22636
rect 20220 22624 20226 22636
rect 20625 22627 20683 22633
rect 20625 22624 20637 22627
rect 20220 22596 20637 22624
rect 20220 22584 20226 22596
rect 20625 22593 20637 22596
rect 20671 22593 20683 22627
rect 20625 22587 20683 22593
rect 17828 22528 19104 22556
rect 19521 22559 19579 22565
rect 17828 22516 17834 22528
rect 19521 22525 19533 22559
rect 19567 22525 19579 22559
rect 19521 22519 19579 22525
rect 19613 22559 19671 22565
rect 19613 22525 19625 22559
rect 19659 22525 19671 22559
rect 19613 22519 19671 22525
rect 16540 22460 16988 22488
rect 18524 22460 19380 22488
rect 16540 22448 16546 22460
rect 16574 22420 16580 22432
rect 15304 22392 16580 22420
rect 16574 22380 16580 22392
rect 16632 22380 16638 22432
rect 16666 22380 16672 22432
rect 16724 22420 16730 22432
rect 18524 22420 18552 22460
rect 16724 22392 18552 22420
rect 19352 22420 19380 22460
rect 19426 22448 19432 22500
rect 19484 22488 19490 22500
rect 19536 22488 19564 22519
rect 19484 22460 19564 22488
rect 19484 22448 19490 22460
rect 19628 22420 19656 22519
rect 19886 22516 19892 22568
rect 19944 22556 19950 22568
rect 20824 22565 20852 22664
rect 20717 22559 20775 22565
rect 20717 22556 20729 22559
rect 19944 22528 20729 22556
rect 19944 22516 19950 22528
rect 20717 22525 20729 22528
rect 20763 22525 20775 22559
rect 20717 22519 20775 22525
rect 20809 22559 20867 22565
rect 20809 22525 20821 22559
rect 20855 22525 20867 22559
rect 20916 22556 20944 22732
rect 21266 22720 21272 22772
rect 21324 22720 21330 22772
rect 23658 22720 23664 22772
rect 23716 22760 23722 22772
rect 24578 22760 24584 22772
rect 23716 22732 24584 22760
rect 23716 22720 23722 22732
rect 24578 22720 24584 22732
rect 24636 22760 24642 22772
rect 24636 22732 24900 22760
rect 24636 22720 24642 22732
rect 23566 22652 23572 22704
rect 23624 22652 23630 22704
rect 24872 22692 24900 22732
rect 25317 22695 25375 22701
rect 25317 22692 25329 22695
rect 24794 22664 25329 22692
rect 25317 22661 25329 22664
rect 25363 22661 25375 22695
rect 25317 22655 25375 22661
rect 21637 22627 21695 22633
rect 21637 22593 21649 22627
rect 21683 22624 21695 22627
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21683 22596 22017 22624
rect 21683 22593 21695 22596
rect 21637 22587 21695 22593
rect 22005 22593 22017 22596
rect 22051 22624 22063 22627
rect 22051 22596 23244 22624
rect 22051 22593 22063 22596
rect 22005 22587 22063 22593
rect 22186 22556 22192 22568
rect 20916 22528 22192 22556
rect 20809 22519 20867 22525
rect 22186 22516 22192 22528
rect 22244 22516 22250 22568
rect 22278 22516 22284 22568
rect 22336 22516 22342 22568
rect 23216 22556 23244 22596
rect 23290 22584 23296 22636
rect 23348 22584 23354 22636
rect 25038 22556 25044 22568
rect 23216 22528 25044 22556
rect 25038 22516 25044 22528
rect 25096 22516 25102 22568
rect 23198 22488 23204 22500
rect 20824 22460 23204 22488
rect 20824 22432 20852 22460
rect 23198 22448 23204 22460
rect 23256 22448 23262 22500
rect 19352 22392 19656 22420
rect 16724 22380 16730 22392
rect 20806 22380 20812 22432
rect 20864 22380 20870 22432
rect 21358 22380 21364 22432
rect 21416 22420 21422 22432
rect 22738 22420 22744 22432
rect 21416 22392 22744 22420
rect 21416 22380 21422 22392
rect 22738 22380 22744 22392
rect 22796 22380 22802 22432
rect 25041 22423 25099 22429
rect 25041 22389 25053 22423
rect 25087 22420 25099 22423
rect 25130 22420 25136 22432
rect 25087 22392 25136 22420
rect 25087 22389 25099 22392
rect 25041 22383 25099 22389
rect 25130 22380 25136 22392
rect 25188 22380 25194 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 7650 22176 7656 22228
rect 7708 22216 7714 22228
rect 12066 22216 12072 22228
rect 7708 22188 12072 22216
rect 7708 22176 7714 22188
rect 12066 22176 12072 22188
rect 12124 22176 12130 22228
rect 12158 22176 12164 22228
rect 12216 22216 12222 22228
rect 12526 22216 12532 22228
rect 12216 22188 12532 22216
rect 12216 22176 12222 22188
rect 12526 22176 12532 22188
rect 12584 22176 12590 22228
rect 14540 22219 14598 22225
rect 14540 22185 14552 22219
rect 14586 22216 14598 22219
rect 14642 22216 14648 22228
rect 14586 22188 14648 22216
rect 14586 22185 14598 22188
rect 14540 22179 14598 22185
rect 14642 22176 14648 22188
rect 14700 22176 14706 22228
rect 17034 22216 17040 22228
rect 15580 22188 17040 22216
rect 2406 22108 2412 22160
rect 2464 22148 2470 22160
rect 2774 22148 2780 22160
rect 2464 22120 2780 22148
rect 2464 22108 2470 22120
rect 2774 22108 2780 22120
rect 2832 22108 2838 22160
rect 2866 22040 2872 22092
rect 2924 22040 2930 22092
rect 6086 22040 6092 22092
rect 6144 22040 6150 22092
rect 8294 22040 8300 22092
rect 8352 22040 8358 22092
rect 9030 22040 9036 22092
rect 9088 22080 9094 22092
rect 10689 22083 10747 22089
rect 10689 22080 10701 22083
rect 9088 22052 10701 22080
rect 9088 22040 9094 22052
rect 10689 22049 10701 22052
rect 10735 22080 10747 22083
rect 11054 22080 11060 22092
rect 10735 22052 11060 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 11054 22040 11060 22052
rect 11112 22040 11118 22092
rect 11330 22040 11336 22092
rect 11388 22080 11394 22092
rect 11388 22052 12204 22080
rect 11388 22040 11394 22052
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 21981 2283 22015
rect 2225 21975 2283 21981
rect 2240 21944 2268 21975
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 22012 4307 22015
rect 4614 22012 4620 22024
rect 4295 21984 4620 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 4614 21972 4620 21984
rect 4672 21972 4678 22024
rect 5537 22015 5595 22021
rect 5537 21981 5549 22015
rect 5583 22012 5595 22015
rect 6362 22012 6368 22024
rect 5583 21984 6368 22012
rect 5583 21981 5595 21984
rect 5537 21975 5595 21981
rect 6362 21972 6368 21984
rect 6420 21972 6426 22024
rect 7374 21972 7380 22024
rect 7432 21972 7438 22024
rect 8941 22015 8999 22021
rect 8941 21981 8953 22015
rect 8987 22012 8999 22015
rect 9493 22015 9551 22021
rect 9493 22012 9505 22015
rect 8987 21984 9505 22012
rect 8987 21981 8999 21984
rect 8941 21975 8999 21981
rect 9493 21981 9505 21984
rect 9539 22012 9551 22015
rect 12176 22012 12204 22052
rect 12250 22040 12256 22092
rect 12308 22080 12314 22092
rect 12437 22083 12495 22089
rect 12437 22080 12449 22083
rect 12308 22052 12449 22080
rect 12308 22040 12314 22052
rect 12437 22049 12449 22052
rect 12483 22049 12495 22083
rect 12437 22043 12495 22049
rect 12618 22040 12624 22092
rect 12676 22080 12682 22092
rect 13630 22080 13636 22092
rect 12676 22052 13636 22080
rect 12676 22040 12682 22052
rect 13630 22040 13636 22052
rect 13688 22080 13694 22092
rect 15580 22080 15608 22188
rect 17034 22176 17040 22188
rect 17092 22176 17098 22228
rect 18414 22176 18420 22228
rect 18472 22216 18478 22228
rect 22830 22216 22836 22228
rect 18472 22188 22836 22216
rect 18472 22176 18478 22188
rect 22830 22176 22836 22188
rect 22888 22176 22894 22228
rect 23198 22176 23204 22228
rect 23256 22216 23262 22228
rect 23474 22216 23480 22228
rect 23256 22188 23480 22216
rect 23256 22176 23262 22188
rect 23474 22176 23480 22188
rect 23532 22216 23538 22228
rect 25314 22216 25320 22228
rect 23532 22188 25320 22216
rect 23532 22176 23538 22188
rect 25314 22176 25320 22188
rect 25372 22176 25378 22228
rect 15654 22108 15660 22160
rect 15712 22148 15718 22160
rect 16482 22148 16488 22160
rect 15712 22120 16488 22148
rect 15712 22108 15718 22120
rect 16482 22108 16488 22120
rect 16540 22148 16546 22160
rect 17770 22148 17776 22160
rect 16540 22120 17776 22148
rect 16540 22108 16546 22120
rect 17770 22108 17776 22120
rect 17828 22108 17834 22160
rect 17862 22108 17868 22160
rect 17920 22148 17926 22160
rect 19886 22148 19892 22160
rect 17920 22120 19892 22148
rect 17920 22108 17926 22120
rect 19886 22108 19892 22120
rect 19944 22108 19950 22160
rect 13688 22052 15608 22080
rect 13688 22040 13694 22052
rect 17034 22040 17040 22092
rect 17092 22040 17098 22092
rect 18046 22080 18052 22092
rect 17144 22052 18052 22080
rect 13725 22015 13783 22021
rect 13725 22012 13737 22015
rect 9539 21984 10272 22012
rect 12176 21984 13737 22012
rect 9539 21981 9551 21984
rect 9493 21975 9551 21981
rect 4890 21944 4896 21956
rect 2240 21916 4896 21944
rect 4890 21904 4896 21916
rect 4948 21904 4954 21956
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 10042 21836 10048 21888
rect 10100 21836 10106 21888
rect 10244 21876 10272 21984
rect 13725 21981 13737 21984
rect 13771 21981 13783 22015
rect 13725 21975 13783 21981
rect 14274 21972 14280 22024
rect 14332 21972 14338 22024
rect 15930 21972 15936 22024
rect 15988 22012 15994 22024
rect 16945 22015 17003 22021
rect 16945 22012 16957 22015
rect 15988 21984 16957 22012
rect 15988 21972 15994 21984
rect 16945 21981 16957 21984
rect 16991 22012 17003 22015
rect 17144 22012 17172 22052
rect 18046 22040 18052 22052
rect 18104 22040 18110 22092
rect 18233 22083 18291 22089
rect 18233 22049 18245 22083
rect 18279 22049 18291 22083
rect 18233 22043 18291 22049
rect 20625 22083 20683 22089
rect 20625 22049 20637 22083
rect 20671 22080 20683 22083
rect 20714 22080 20720 22092
rect 20671 22052 20720 22080
rect 20671 22049 20683 22052
rect 20625 22043 20683 22049
rect 18248 22012 18276 22043
rect 20714 22040 20720 22052
rect 20772 22040 20778 22092
rect 23474 22080 23480 22092
rect 23308 22052 23480 22080
rect 16991 21984 17172 22012
rect 17972 21984 18276 22012
rect 16991 21981 17003 21984
rect 16945 21975 17003 21981
rect 10962 21904 10968 21956
rect 11020 21904 11026 21956
rect 11422 21904 11428 21956
rect 11480 21904 11486 21956
rect 13538 21904 13544 21956
rect 13596 21904 13602 21956
rect 15838 21944 15844 21956
rect 15778 21916 15844 21944
rect 15838 21904 15844 21916
rect 15896 21904 15902 21956
rect 17972 21944 18000 21984
rect 19334 21972 19340 22024
rect 19392 22012 19398 22024
rect 20349 22015 20407 22021
rect 20349 22012 20361 22015
rect 19392 21984 20361 22012
rect 19392 21972 19398 21984
rect 20349 21981 20361 21984
rect 20395 21981 20407 22015
rect 20349 21975 20407 21981
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22462 22012 22468 22024
rect 22152 21984 22468 22012
rect 22152 21972 22158 21984
rect 22462 21972 22468 21984
rect 22520 21972 22526 22024
rect 22738 21972 22744 22024
rect 22796 21972 22802 22024
rect 23198 21972 23204 22024
rect 23256 21972 23262 22024
rect 16224 21916 18000 21944
rect 18049 21947 18107 21953
rect 16224 21888 16252 21916
rect 18049 21913 18061 21947
rect 18095 21944 18107 21947
rect 18598 21944 18604 21956
rect 18095 21916 18604 21944
rect 18095 21913 18107 21916
rect 18049 21907 18107 21913
rect 18598 21904 18604 21916
rect 18656 21904 18662 21956
rect 18690 21904 18696 21956
rect 18748 21904 18754 21956
rect 19426 21944 19432 21956
rect 18892 21916 19432 21944
rect 18892 21888 18920 21916
rect 19426 21904 19432 21916
rect 19484 21904 19490 21956
rect 19518 21904 19524 21956
rect 19576 21904 19582 21956
rect 21174 21904 21180 21956
rect 21232 21904 21238 21956
rect 23308 21944 23336 22052
rect 23474 22040 23480 22052
rect 23532 22040 23538 22092
rect 24854 22040 24860 22092
rect 24912 22080 24918 22092
rect 25041 22083 25099 22089
rect 25041 22080 25053 22083
rect 24912 22052 25053 22080
rect 24912 22040 24918 22052
rect 25041 22049 25053 22052
rect 25087 22049 25099 22083
rect 25041 22043 25099 22049
rect 25130 22040 25136 22092
rect 25188 22040 25194 22092
rect 21928 21916 23336 21944
rect 11974 21876 11980 21888
rect 10244 21848 11980 21876
rect 11974 21836 11980 21848
rect 12032 21836 12038 21888
rect 12250 21836 12256 21888
rect 12308 21876 12314 21888
rect 12713 21879 12771 21885
rect 12713 21876 12725 21879
rect 12308 21848 12725 21876
rect 12308 21836 12314 21848
rect 12713 21845 12725 21848
rect 12759 21845 12771 21879
rect 12713 21839 12771 21845
rect 16025 21879 16083 21885
rect 16025 21845 16037 21879
rect 16071 21876 16083 21879
rect 16206 21876 16212 21888
rect 16071 21848 16212 21876
rect 16071 21845 16083 21848
rect 16025 21839 16083 21845
rect 16206 21836 16212 21848
rect 16264 21836 16270 21888
rect 16485 21879 16543 21885
rect 16485 21845 16497 21879
rect 16531 21876 16543 21879
rect 16666 21876 16672 21888
rect 16531 21848 16672 21876
rect 16531 21845 16543 21848
rect 16485 21839 16543 21845
rect 16666 21836 16672 21848
rect 16724 21836 16730 21888
rect 16850 21836 16856 21888
rect 16908 21836 16914 21888
rect 17034 21836 17040 21888
rect 17092 21876 17098 21888
rect 17494 21876 17500 21888
rect 17092 21848 17500 21876
rect 17092 21836 17098 21848
rect 17494 21836 17500 21848
rect 17552 21836 17558 21888
rect 17678 21836 17684 21888
rect 17736 21836 17742 21888
rect 17862 21836 17868 21888
rect 17920 21876 17926 21888
rect 18141 21879 18199 21885
rect 18141 21876 18153 21879
rect 17920 21848 18153 21876
rect 17920 21836 17926 21848
rect 18141 21845 18153 21848
rect 18187 21845 18199 21879
rect 18141 21839 18199 21845
rect 18230 21836 18236 21888
rect 18288 21876 18294 21888
rect 18874 21876 18880 21888
rect 18288 21848 18880 21876
rect 18288 21836 18294 21848
rect 18874 21836 18880 21848
rect 18932 21836 18938 21888
rect 18966 21836 18972 21888
rect 19024 21876 19030 21888
rect 19613 21879 19671 21885
rect 19613 21876 19625 21879
rect 19024 21848 19625 21876
rect 19024 21836 19030 21848
rect 19613 21845 19625 21848
rect 19659 21845 19671 21879
rect 19613 21839 19671 21845
rect 20254 21836 20260 21888
rect 20312 21876 20318 21888
rect 21928 21876 21956 21916
rect 20312 21848 21956 21876
rect 20312 21836 20318 21848
rect 22002 21836 22008 21888
rect 22060 21876 22066 21888
rect 22097 21879 22155 21885
rect 22097 21876 22109 21879
rect 22060 21848 22109 21876
rect 22060 21836 22066 21848
rect 22097 21845 22109 21848
rect 22143 21845 22155 21879
rect 22097 21839 22155 21845
rect 22557 21879 22615 21885
rect 22557 21845 22569 21879
rect 22603 21876 22615 21879
rect 24210 21876 24216 21888
rect 22603 21848 24216 21876
rect 22603 21845 22615 21848
rect 22557 21839 22615 21845
rect 24210 21836 24216 21848
rect 24268 21836 24274 21888
rect 24578 21836 24584 21888
rect 24636 21836 24642 21888
rect 24670 21836 24676 21888
rect 24728 21876 24734 21888
rect 24949 21879 25007 21885
rect 24949 21876 24961 21879
rect 24728 21848 24961 21876
rect 24728 21836 24734 21848
rect 24949 21845 24961 21848
rect 24995 21845 25007 21879
rect 24949 21839 25007 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 2222 21632 2228 21684
rect 2280 21672 2286 21684
rect 9398 21672 9404 21684
rect 2280 21644 9404 21672
rect 2280 21632 2286 21644
rect 9398 21632 9404 21644
rect 9456 21632 9462 21684
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 12621 21675 12679 21681
rect 12621 21672 12633 21675
rect 10100 21644 12633 21672
rect 10100 21632 10106 21644
rect 12621 21641 12633 21644
rect 12667 21641 12679 21675
rect 12621 21635 12679 21641
rect 13170 21632 13176 21684
rect 13228 21672 13234 21684
rect 13354 21672 13360 21684
rect 13228 21644 13360 21672
rect 13228 21632 13234 21644
rect 13354 21632 13360 21644
rect 13412 21632 13418 21684
rect 14277 21675 14335 21681
rect 14277 21641 14289 21675
rect 14323 21672 14335 21675
rect 17678 21672 17684 21684
rect 14323 21644 17684 21672
rect 14323 21641 14335 21644
rect 14277 21635 14335 21641
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 17788 21644 21036 21672
rect 1673 21607 1731 21613
rect 1673 21573 1685 21607
rect 1719 21604 1731 21607
rect 2133 21607 2191 21613
rect 2133 21604 2145 21607
rect 1719 21576 2145 21604
rect 1719 21573 1731 21576
rect 1673 21567 1731 21573
rect 2133 21573 2145 21576
rect 2179 21604 2191 21607
rect 3418 21604 3424 21616
rect 2179 21576 3424 21604
rect 2179 21573 2191 21576
rect 2133 21567 2191 21573
rect 3418 21564 3424 21576
rect 3476 21564 3482 21616
rect 8478 21604 8484 21616
rect 4816 21576 8484 21604
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21536 3019 21539
rect 4154 21536 4160 21548
rect 3007 21508 4160 21536
rect 3007 21505 3019 21508
rect 2961 21499 3019 21505
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4816 21545 4844 21576
rect 8478 21564 8484 21576
rect 8536 21564 8542 21616
rect 12713 21607 12771 21613
rect 12713 21573 12725 21607
rect 12759 21604 12771 21607
rect 16482 21604 16488 21616
rect 12759 21576 16488 21604
rect 12759 21573 12771 21576
rect 12713 21567 12771 21573
rect 16482 21564 16488 21576
rect 16540 21564 16546 21616
rect 17788 21604 17816 21644
rect 16776 21576 17816 21604
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21505 4859 21539
rect 4801 21499 4859 21505
rect 6730 21496 6736 21548
rect 6788 21496 6794 21548
rect 7374 21496 7380 21548
rect 7432 21496 7438 21548
rect 9030 21496 9036 21548
rect 9088 21496 9094 21548
rect 10410 21496 10416 21548
rect 10468 21536 10474 21548
rect 11057 21539 11115 21545
rect 11057 21536 11069 21539
rect 10468 21508 11069 21536
rect 10468 21496 10474 21508
rect 11057 21505 11069 21508
rect 11103 21536 11115 21539
rect 11241 21539 11299 21545
rect 11241 21536 11253 21539
rect 11103 21508 11253 21536
rect 11103 21505 11115 21508
rect 11057 21499 11115 21505
rect 11241 21505 11253 21508
rect 11287 21536 11299 21539
rect 11422 21536 11428 21548
rect 11287 21508 11428 21536
rect 11287 21505 11299 21508
rect 11241 21499 11299 21505
rect 11422 21496 11428 21508
rect 11480 21536 11486 21548
rect 12250 21536 12256 21548
rect 11480 21508 12256 21536
rect 11480 21496 11486 21508
rect 12250 21496 12256 21508
rect 12308 21496 12314 21548
rect 12544 21508 14136 21536
rect 3510 21428 3516 21480
rect 3568 21428 3574 21480
rect 5074 21428 5080 21480
rect 5132 21428 5138 21480
rect 7282 21428 7288 21480
rect 7340 21468 7346 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7340 21440 7665 21468
rect 7340 21428 7346 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 7653 21431 7711 21437
rect 9306 21428 9312 21480
rect 9364 21428 9370 21480
rect 9398 21428 9404 21480
rect 9456 21468 9462 21480
rect 9456 21440 10456 21468
rect 9456 21428 9462 21440
rect 1857 21403 1915 21409
rect 1857 21369 1869 21403
rect 1903 21400 1915 21403
rect 10428 21400 10456 21440
rect 10686 21428 10692 21480
rect 10744 21468 10750 21480
rect 12544 21468 12572 21508
rect 10744 21440 12572 21468
rect 10744 21428 10750 21440
rect 12618 21428 12624 21480
rect 12676 21468 12682 21480
rect 12897 21471 12955 21477
rect 12897 21468 12909 21471
rect 12676 21440 12909 21468
rect 12676 21428 12682 21440
rect 12897 21437 12909 21440
rect 12943 21468 12955 21471
rect 13446 21468 13452 21480
rect 12943 21440 13452 21468
rect 12943 21437 12955 21440
rect 12897 21431 12955 21437
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 14108 21468 14136 21508
rect 14182 21496 14188 21548
rect 14240 21496 14246 21548
rect 15194 21536 15200 21548
rect 14292 21508 15200 21536
rect 14292 21468 14320 21508
rect 15194 21496 15200 21508
rect 15252 21536 15258 21548
rect 15381 21539 15439 21545
rect 15381 21536 15393 21539
rect 15252 21508 15393 21536
rect 15252 21496 15258 21508
rect 15381 21505 15393 21508
rect 15427 21505 15439 21539
rect 15381 21499 15439 21505
rect 15930 21496 15936 21548
rect 15988 21536 15994 21548
rect 16393 21539 16451 21545
rect 16393 21536 16405 21539
rect 15988 21508 16405 21536
rect 15988 21496 15994 21508
rect 16393 21505 16405 21508
rect 16439 21505 16451 21539
rect 16393 21499 16451 21505
rect 14108 21440 14320 21468
rect 14369 21471 14427 21477
rect 14369 21437 14381 21471
rect 14415 21468 14427 21471
rect 15102 21468 15108 21480
rect 14415 21440 15108 21468
rect 14415 21437 14427 21440
rect 14369 21431 14427 21437
rect 15102 21428 15108 21440
rect 15160 21428 15166 21480
rect 15470 21428 15476 21480
rect 15528 21428 15534 21480
rect 15654 21428 15660 21480
rect 15712 21428 15718 21480
rect 16298 21428 16304 21480
rect 16356 21468 16362 21480
rect 16776 21468 16804 21576
rect 19150 21564 19156 21616
rect 19208 21604 19214 21616
rect 21008 21604 21036 21644
rect 21082 21632 21088 21684
rect 21140 21672 21146 21684
rect 21140 21644 22876 21672
rect 21140 21632 21146 21644
rect 22738 21604 22744 21616
rect 19208 21576 20944 21604
rect 21008 21576 22744 21604
rect 19208 21564 19214 21576
rect 17402 21496 17408 21548
rect 17460 21496 17466 21548
rect 18233 21539 18291 21545
rect 18233 21505 18245 21539
rect 18279 21536 18291 21539
rect 18874 21536 18880 21548
rect 18279 21508 18880 21536
rect 18279 21505 18291 21508
rect 18233 21499 18291 21505
rect 18874 21496 18880 21508
rect 18932 21496 18938 21548
rect 19242 21496 19248 21548
rect 19300 21536 19306 21548
rect 19300 21508 19840 21536
rect 19300 21496 19306 21508
rect 16356 21440 16804 21468
rect 16356 21428 16362 21440
rect 16942 21428 16948 21480
rect 17000 21468 17006 21480
rect 17497 21471 17555 21477
rect 17497 21468 17509 21471
rect 17000 21440 17509 21468
rect 17000 21428 17006 21440
rect 17497 21437 17509 21440
rect 17543 21437 17555 21471
rect 17497 21431 17555 21437
rect 17589 21471 17647 21477
rect 17589 21437 17601 21471
rect 17635 21437 17647 21471
rect 19702 21468 19708 21480
rect 17589 21431 17647 21437
rect 18248 21440 19708 21468
rect 14458 21400 14464 21412
rect 1903 21372 7604 21400
rect 10428 21372 14464 21400
rect 1903 21369 1915 21372
rect 1857 21363 1915 21369
rect 6546 21292 6552 21344
rect 6604 21292 6610 21344
rect 7576 21332 7604 21372
rect 14458 21360 14464 21372
rect 14516 21360 14522 21412
rect 15013 21403 15071 21409
rect 15013 21369 15025 21403
rect 15059 21400 15071 21403
rect 17126 21400 17132 21412
rect 15059 21372 17132 21400
rect 15059 21369 15071 21372
rect 15013 21363 15071 21369
rect 17126 21360 17132 21372
rect 17184 21360 17190 21412
rect 17310 21360 17316 21412
rect 17368 21400 17374 21412
rect 17604 21400 17632 21431
rect 17368 21372 17632 21400
rect 17368 21360 17374 21372
rect 10686 21332 10692 21344
rect 7576 21304 10692 21332
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 10778 21292 10784 21344
rect 10836 21292 10842 21344
rect 10870 21292 10876 21344
rect 10928 21332 10934 21344
rect 12253 21335 12311 21341
rect 12253 21332 12265 21335
rect 10928 21304 12265 21332
rect 10928 21292 10934 21304
rect 12253 21301 12265 21304
rect 12299 21301 12311 21335
rect 12253 21295 12311 21301
rect 12802 21292 12808 21344
rect 12860 21332 12866 21344
rect 13817 21335 13875 21341
rect 13817 21332 13829 21335
rect 12860 21304 13829 21332
rect 12860 21292 12866 21304
rect 13817 21301 13829 21304
rect 13863 21301 13875 21335
rect 13817 21295 13875 21301
rect 16022 21292 16028 21344
rect 16080 21332 16086 21344
rect 16117 21335 16175 21341
rect 16117 21332 16129 21335
rect 16080 21304 16129 21332
rect 16080 21292 16086 21304
rect 16117 21301 16129 21304
rect 16163 21301 16175 21335
rect 16117 21295 16175 21301
rect 17037 21335 17095 21341
rect 17037 21301 17049 21335
rect 17083 21332 17095 21335
rect 18248 21332 18276 21440
rect 19702 21428 19708 21440
rect 19760 21428 19766 21480
rect 19812 21468 19840 21508
rect 20254 21496 20260 21548
rect 20312 21536 20318 21548
rect 20809 21539 20867 21545
rect 20809 21536 20821 21539
rect 20312 21508 20821 21536
rect 20312 21496 20318 21508
rect 20809 21505 20821 21508
rect 20855 21505 20867 21539
rect 20916 21536 20944 21576
rect 22738 21564 22744 21576
rect 22796 21564 22802 21616
rect 21910 21536 21916 21548
rect 20916 21508 21916 21536
rect 20809 21499 20867 21505
rect 21910 21496 21916 21508
rect 21968 21496 21974 21548
rect 22186 21496 22192 21548
rect 22244 21536 22250 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22244 21508 22385 21536
rect 22244 21496 22250 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22848 21536 22876 21644
rect 23109 21607 23167 21613
rect 23109 21573 23121 21607
rect 23155 21604 23167 21607
rect 23658 21604 23664 21616
rect 23155 21576 23664 21604
rect 23155 21573 23167 21576
rect 23109 21567 23167 21573
rect 23658 21564 23664 21576
rect 23716 21564 23722 21616
rect 25222 21604 25228 21616
rect 24886 21576 25228 21604
rect 25222 21564 25228 21576
rect 25280 21604 25286 21616
rect 25409 21607 25467 21613
rect 25409 21604 25421 21607
rect 25280 21576 25421 21604
rect 25280 21564 25286 21576
rect 25409 21573 25421 21576
rect 25455 21573 25467 21607
rect 25409 21567 25467 21573
rect 22373 21499 22431 21505
rect 22664 21508 22876 21536
rect 20901 21471 20959 21477
rect 20901 21468 20913 21471
rect 19812 21440 20913 21468
rect 20901 21437 20913 21440
rect 20947 21437 20959 21471
rect 20901 21431 20959 21437
rect 21085 21471 21143 21477
rect 21085 21437 21097 21471
rect 21131 21468 21143 21471
rect 21266 21468 21272 21480
rect 21131 21440 21272 21468
rect 21131 21437 21143 21440
rect 21085 21431 21143 21437
rect 21266 21428 21272 21440
rect 21324 21428 21330 21480
rect 21450 21428 21456 21480
rect 21508 21468 21514 21480
rect 22664 21477 22692 21508
rect 23290 21496 23296 21548
rect 23348 21536 23354 21548
rect 23385 21539 23443 21545
rect 23385 21536 23397 21539
rect 23348 21508 23397 21536
rect 23348 21496 23354 21508
rect 23385 21505 23397 21508
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 21545 21471 21603 21477
rect 21545 21468 21557 21471
rect 21508 21440 21557 21468
rect 21508 21428 21514 21440
rect 21545 21437 21557 21440
rect 21591 21468 21603 21471
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 21591 21440 22477 21468
rect 21591 21437 21603 21440
rect 21545 21431 21603 21437
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21437 22707 21471
rect 22649 21431 22707 21437
rect 23661 21471 23719 21477
rect 23661 21437 23673 21471
rect 23707 21468 23719 21471
rect 25130 21468 25136 21480
rect 23707 21440 25136 21468
rect 23707 21437 23719 21440
rect 23661 21431 23719 21437
rect 25130 21428 25136 21440
rect 25188 21428 25194 21480
rect 18322 21360 18328 21412
rect 18380 21400 18386 21412
rect 22005 21403 22063 21409
rect 22005 21400 22017 21403
rect 18380 21372 22017 21400
rect 18380 21360 18386 21372
rect 22005 21369 22017 21372
rect 22051 21369 22063 21403
rect 22005 21363 22063 21369
rect 17083 21304 18276 21332
rect 17083 21301 17095 21304
rect 17037 21295 17095 21301
rect 19334 21292 19340 21344
rect 19392 21332 19398 21344
rect 19521 21335 19579 21341
rect 19521 21332 19533 21335
rect 19392 21304 19533 21332
rect 19392 21292 19398 21304
rect 19521 21301 19533 21304
rect 19567 21301 19579 21335
rect 19521 21295 19579 21301
rect 19978 21292 19984 21344
rect 20036 21332 20042 21344
rect 20441 21335 20499 21341
rect 20441 21332 20453 21335
rect 20036 21304 20453 21332
rect 20036 21292 20042 21304
rect 20441 21301 20453 21304
rect 20487 21301 20499 21335
rect 20441 21295 20499 21301
rect 23750 21292 23756 21344
rect 23808 21332 23814 21344
rect 25133 21335 25191 21341
rect 25133 21332 25145 21335
rect 23808 21304 25145 21332
rect 23808 21292 23814 21304
rect 25133 21301 25145 21304
rect 25179 21301 25191 21335
rect 25133 21295 25191 21301
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 3970 21088 3976 21140
rect 4028 21128 4034 21140
rect 6365 21131 6423 21137
rect 6365 21128 6377 21131
rect 4028 21100 6377 21128
rect 4028 21088 4034 21100
rect 6365 21097 6377 21100
rect 6411 21128 6423 21131
rect 9214 21128 9220 21140
rect 6411 21100 9220 21128
rect 6411 21097 6423 21100
rect 6365 21091 6423 21097
rect 9214 21088 9220 21100
rect 9272 21088 9278 21140
rect 10410 21088 10416 21140
rect 10468 21128 10474 21140
rect 12897 21131 12955 21137
rect 10468 21100 12848 21128
rect 10468 21088 10474 21100
rect 3418 21020 3424 21072
rect 3476 21060 3482 21072
rect 3476 21032 7512 21060
rect 3476 21020 3482 21032
rect 2774 20952 2780 21004
rect 2832 20952 2838 21004
rect 4246 20952 4252 21004
rect 4304 20992 4310 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4304 20964 4445 20992
rect 4304 20952 4310 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 7006 20952 7012 21004
rect 7064 20992 7070 21004
rect 7377 20995 7435 21001
rect 7377 20992 7389 20995
rect 7064 20964 7389 20992
rect 7064 20952 7070 20964
rect 7377 20961 7389 20964
rect 7423 20961 7435 20995
rect 7484 20992 7512 21032
rect 8478 21020 8484 21072
rect 8536 21060 8542 21072
rect 9953 21063 10011 21069
rect 9953 21060 9965 21063
rect 8536 21032 9965 21060
rect 8536 21020 8542 21032
rect 9953 21029 9965 21032
rect 9999 21029 10011 21063
rect 9953 21023 10011 21029
rect 10042 21020 10048 21072
rect 10100 21060 10106 21072
rect 10778 21060 10784 21072
rect 10100 21032 10784 21060
rect 10100 21020 10106 21032
rect 10502 20992 10508 21004
rect 7484 20964 10508 20992
rect 7377 20955 7435 20961
rect 10502 20952 10508 20964
rect 10560 20952 10566 21004
rect 10612 21001 10640 21032
rect 10778 21020 10784 21032
rect 10836 21020 10842 21072
rect 12434 21020 12440 21072
rect 12492 21060 12498 21072
rect 12820 21060 12848 21100
rect 12897 21097 12909 21131
rect 12943 21128 12955 21131
rect 13630 21128 13636 21140
rect 12943 21100 13636 21128
rect 12943 21097 12955 21100
rect 12897 21091 12955 21097
rect 13630 21088 13636 21100
rect 13688 21088 13694 21140
rect 14458 21088 14464 21140
rect 14516 21088 14522 21140
rect 17954 21128 17960 21140
rect 15948 21100 17960 21128
rect 15473 21063 15531 21069
rect 15473 21060 15485 21063
rect 12492 21032 12572 21060
rect 12820 21032 15485 21060
rect 12492 21020 12498 21032
rect 10597 20995 10655 21001
rect 10597 20961 10609 20995
rect 10643 20961 10655 20995
rect 10597 20955 10655 20961
rect 11054 20952 11060 21004
rect 11112 20992 11118 21004
rect 11149 20995 11207 21001
rect 11149 20992 11161 20995
rect 11112 20964 11161 20992
rect 11112 20952 11118 20964
rect 11149 20961 11161 20964
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 11425 20995 11483 21001
rect 11425 20961 11437 20995
rect 11471 20992 11483 20995
rect 12544 20992 12572 21032
rect 15473 21029 15485 21032
rect 15519 21029 15531 21063
rect 15473 21023 15531 21029
rect 13725 20995 13783 21001
rect 13725 20992 13737 20995
rect 11471 20964 12480 20992
rect 12544 20964 13737 20992
rect 11471 20961 11483 20964
rect 11425 20955 11483 20961
rect 12452 20936 12480 20964
rect 13725 20961 13737 20964
rect 13771 20961 13783 20995
rect 13725 20955 13783 20961
rect 14734 20952 14740 21004
rect 14792 20992 14798 21004
rect 15948 21001 15976 21100
rect 17954 21088 17960 21100
rect 18012 21088 18018 21140
rect 18506 21088 18512 21140
rect 18564 21128 18570 21140
rect 18690 21128 18696 21140
rect 18564 21100 18696 21128
rect 18564 21088 18570 21100
rect 18690 21088 18696 21100
rect 18748 21128 18754 21140
rect 18877 21131 18935 21137
rect 18877 21128 18889 21131
rect 18748 21100 18889 21128
rect 18748 21088 18754 21100
rect 18877 21097 18889 21100
rect 18923 21097 18935 21131
rect 18877 21091 18935 21097
rect 20438 21088 20444 21140
rect 20496 21128 20502 21140
rect 21177 21131 21235 21137
rect 21177 21128 21189 21131
rect 20496 21100 21189 21128
rect 20496 21088 20502 21100
rect 21177 21097 21189 21100
rect 21223 21097 21235 21131
rect 21177 21091 21235 21097
rect 21910 21088 21916 21140
rect 21968 21128 21974 21140
rect 22646 21128 22652 21140
rect 21968 21100 22652 21128
rect 21968 21088 21974 21100
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 22738 21088 22744 21140
rect 22796 21128 22802 21140
rect 24029 21131 24087 21137
rect 24029 21128 24041 21131
rect 22796 21100 24041 21128
rect 22796 21088 22802 21100
rect 24029 21097 24041 21100
rect 24075 21097 24087 21131
rect 24029 21091 24087 21097
rect 16669 21063 16727 21069
rect 16669 21029 16681 21063
rect 16715 21029 16727 21063
rect 17402 21060 17408 21072
rect 16669 21023 16727 21029
rect 17236 21032 17408 21060
rect 15933 20995 15991 21001
rect 15933 20992 15945 20995
rect 14792 20964 15945 20992
rect 14792 20952 14798 20964
rect 15933 20961 15945 20964
rect 15979 20961 15991 20995
rect 15933 20955 15991 20961
rect 16025 20995 16083 21001
rect 16025 20961 16037 20995
rect 16071 20961 16083 20995
rect 16025 20955 16083 20961
rect 2222 20884 2228 20936
rect 2280 20884 2286 20936
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20924 4215 20927
rect 5718 20924 5724 20936
rect 4203 20896 5724 20924
rect 4203 20893 4215 20896
rect 4157 20887 4215 20893
rect 5718 20884 5724 20896
rect 5776 20884 5782 20936
rect 5997 20927 6055 20933
rect 5997 20893 6009 20927
rect 6043 20924 6055 20927
rect 6270 20924 6276 20936
rect 6043 20896 6276 20924
rect 6043 20893 6055 20896
rect 5997 20887 6055 20893
rect 6270 20884 6276 20896
rect 6328 20884 6334 20936
rect 6914 20884 6920 20936
rect 6972 20884 6978 20936
rect 9306 20884 9312 20936
rect 9364 20924 9370 20936
rect 9364 20896 11192 20924
rect 9364 20884 9370 20896
rect 11164 20868 11192 20896
rect 12434 20884 12440 20936
rect 12492 20884 12498 20936
rect 12986 20884 12992 20936
rect 13044 20924 13050 20936
rect 13541 20927 13599 20933
rect 13541 20924 13553 20927
rect 13044 20896 13553 20924
rect 13044 20884 13050 20896
rect 13541 20893 13553 20896
rect 13587 20893 13599 20927
rect 15470 20924 15476 20936
rect 13541 20887 13599 20893
rect 13924 20896 15476 20924
rect 6730 20816 6736 20868
rect 6788 20856 6794 20868
rect 10962 20856 10968 20868
rect 6788 20828 10968 20856
rect 6788 20816 6794 20828
rect 10962 20816 10968 20828
rect 11020 20816 11026 20868
rect 11146 20816 11152 20868
rect 11204 20816 11210 20868
rect 11422 20816 11428 20868
rect 11480 20856 11486 20868
rect 11480 20828 11914 20856
rect 11480 20816 11486 20828
rect 13262 20816 13268 20868
rect 13320 20856 13326 20868
rect 13924 20856 13952 20896
rect 15470 20884 15476 20896
rect 15528 20884 15534 20936
rect 13320 20828 13952 20856
rect 13320 20816 13326 20828
rect 13998 20816 14004 20868
rect 14056 20856 14062 20868
rect 14369 20859 14427 20865
rect 14369 20856 14381 20859
rect 14056 20828 14381 20856
rect 14056 20816 14062 20828
rect 14369 20825 14381 20828
rect 14415 20825 14427 20859
rect 14369 20819 14427 20825
rect 15838 20816 15844 20868
rect 15896 20816 15902 20868
rect 15930 20816 15936 20868
rect 15988 20856 15994 20868
rect 16040 20856 16068 20955
rect 16482 20884 16488 20936
rect 16540 20924 16546 20936
rect 16684 20924 16712 21023
rect 17236 21001 17264 21032
rect 17402 21020 17408 21032
rect 17460 21020 17466 21072
rect 17678 21020 17684 21072
rect 17736 21060 17742 21072
rect 17865 21063 17923 21069
rect 17865 21060 17877 21063
rect 17736 21032 17877 21060
rect 17736 21020 17742 21032
rect 17865 21029 17877 21032
rect 17911 21029 17923 21063
rect 17865 21023 17923 21029
rect 22002 21020 22008 21072
rect 22060 21060 22066 21072
rect 22060 21032 23428 21060
rect 22060 21020 22066 21032
rect 17221 20995 17279 21001
rect 17221 20961 17233 20995
rect 17267 20961 17279 20995
rect 17221 20955 17279 20961
rect 18322 20952 18328 21004
rect 18380 20952 18386 21004
rect 18509 20995 18567 21001
rect 18509 20961 18521 20995
rect 18555 20992 18567 20995
rect 18690 20992 18696 21004
rect 18555 20964 18696 20992
rect 18555 20961 18567 20964
rect 18509 20955 18567 20961
rect 18690 20952 18696 20964
rect 18748 20992 18754 21004
rect 19705 20995 19763 21001
rect 19705 20992 19717 20995
rect 18748 20964 19717 20992
rect 18748 20952 18754 20964
rect 19705 20961 19717 20964
rect 19751 20961 19763 20995
rect 19705 20955 19763 20961
rect 20898 20952 20904 21004
rect 20956 20992 20962 21004
rect 21818 20992 21824 21004
rect 20956 20964 21824 20992
rect 20956 20952 20962 20964
rect 21818 20952 21824 20964
rect 21876 20952 21882 21004
rect 21910 20952 21916 21004
rect 21968 20992 21974 21004
rect 23400 21001 23428 21032
rect 22189 20995 22247 21001
rect 22189 20992 22201 20995
rect 21968 20964 22201 20992
rect 21968 20952 21974 20964
rect 22189 20961 22201 20964
rect 22235 20961 22247 20995
rect 22189 20955 22247 20961
rect 23385 20995 23443 21001
rect 23385 20961 23397 20995
rect 23431 20961 23443 20995
rect 23385 20955 23443 20961
rect 25038 20952 25044 21004
rect 25096 20992 25102 21004
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 25096 20964 25145 20992
rect 25096 20952 25102 20964
rect 25133 20961 25145 20964
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 16540 20896 16712 20924
rect 16540 20884 16546 20896
rect 17678 20884 17684 20936
rect 17736 20924 17742 20936
rect 17736 20896 19196 20924
rect 17736 20884 17742 20896
rect 15988 20828 16068 20856
rect 16132 20828 16804 20856
rect 15988 20816 15994 20828
rect 5810 20748 5816 20800
rect 5868 20748 5874 20800
rect 9306 20748 9312 20800
rect 9364 20748 9370 20800
rect 10318 20748 10324 20800
rect 10376 20748 10382 20800
rect 10410 20748 10416 20800
rect 10468 20748 10474 20800
rect 10502 20748 10508 20800
rect 10560 20788 10566 20800
rect 10870 20788 10876 20800
rect 10560 20760 10876 20788
rect 10560 20748 10566 20760
rect 10870 20748 10876 20760
rect 10928 20748 10934 20800
rect 13630 20748 13636 20800
rect 13688 20788 13694 20800
rect 14090 20788 14096 20800
rect 13688 20760 14096 20788
rect 13688 20748 13694 20760
rect 14090 20748 14096 20760
rect 14148 20748 14154 20800
rect 15470 20748 15476 20800
rect 15528 20788 15534 20800
rect 16132 20788 16160 20828
rect 15528 20760 16160 20788
rect 16776 20788 16804 20828
rect 17034 20816 17040 20868
rect 17092 20816 17098 20868
rect 18233 20859 18291 20865
rect 18233 20825 18245 20859
rect 18279 20856 18291 20859
rect 19058 20856 19064 20868
rect 18279 20828 19064 20856
rect 18279 20825 18291 20828
rect 18233 20819 18291 20825
rect 19058 20816 19064 20828
rect 19116 20816 19122 20868
rect 17129 20791 17187 20797
rect 17129 20788 17141 20791
rect 16776 20760 17141 20788
rect 15528 20748 15534 20760
rect 17129 20757 17141 20760
rect 17175 20757 17187 20791
rect 17129 20751 17187 20757
rect 17402 20748 17408 20800
rect 17460 20788 17466 20800
rect 17586 20788 17592 20800
rect 17460 20760 17592 20788
rect 17460 20748 17466 20760
rect 17586 20748 17592 20760
rect 17644 20748 17650 20800
rect 19168 20788 19196 20896
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 19429 20927 19487 20933
rect 19429 20924 19441 20927
rect 19392 20896 19441 20924
rect 19392 20884 19398 20896
rect 19429 20893 19441 20896
rect 19475 20893 19487 20927
rect 21836 20924 21864 20952
rect 22005 20927 22063 20933
rect 22005 20924 22017 20927
rect 21836 20896 22017 20924
rect 19429 20887 19487 20893
rect 22005 20893 22017 20896
rect 22051 20893 22063 20927
rect 22005 20887 22063 20893
rect 23474 20884 23480 20936
rect 23532 20924 23538 20936
rect 24949 20927 25007 20933
rect 24949 20924 24961 20927
rect 23532 20896 24961 20924
rect 23532 20884 23538 20896
rect 24949 20893 24961 20896
rect 24995 20893 25007 20927
rect 24949 20887 25007 20893
rect 20254 20816 20260 20868
rect 20312 20816 20318 20868
rect 20990 20816 20996 20868
rect 21048 20856 21054 20868
rect 22097 20859 22155 20865
rect 22097 20856 22109 20859
rect 21048 20828 22109 20856
rect 21048 20816 21054 20828
rect 22097 20825 22109 20828
rect 22143 20825 22155 20859
rect 22097 20819 22155 20825
rect 22646 20816 22652 20868
rect 22704 20856 22710 20868
rect 23201 20859 23259 20865
rect 23201 20856 23213 20859
rect 22704 20828 23213 20856
rect 22704 20816 22710 20828
rect 23201 20825 23213 20828
rect 23247 20825 23259 20859
rect 23201 20819 23259 20825
rect 23293 20859 23351 20865
rect 23293 20825 23305 20859
rect 23339 20856 23351 20859
rect 23382 20856 23388 20868
rect 23339 20828 23388 20856
rect 23339 20825 23351 20828
rect 23293 20819 23351 20825
rect 23382 20816 23388 20828
rect 23440 20816 23446 20868
rect 23658 20816 23664 20868
rect 23716 20856 23722 20868
rect 23842 20856 23848 20868
rect 23716 20828 23848 20856
rect 23716 20816 23722 20828
rect 23842 20816 23848 20828
rect 23900 20856 23906 20868
rect 23937 20859 23995 20865
rect 23937 20856 23949 20859
rect 23900 20828 23949 20856
rect 23900 20816 23906 20828
rect 23937 20825 23949 20828
rect 23983 20856 23995 20859
rect 25222 20856 25228 20868
rect 23983 20828 25228 20856
rect 23983 20825 23995 20828
rect 23937 20819 23995 20825
rect 25222 20816 25228 20828
rect 25280 20816 25286 20868
rect 21082 20788 21088 20800
rect 19168 20760 21088 20788
rect 21082 20748 21088 20760
rect 21140 20748 21146 20800
rect 21634 20748 21640 20800
rect 21692 20748 21698 20800
rect 22830 20748 22836 20800
rect 22888 20748 22894 20800
rect 24578 20748 24584 20800
rect 24636 20748 24642 20800
rect 24854 20748 24860 20800
rect 24912 20788 24918 20800
rect 25041 20791 25099 20797
rect 25041 20788 25053 20791
rect 24912 20760 25053 20788
rect 24912 20748 24918 20760
rect 25041 20757 25053 20760
rect 25087 20757 25099 20791
rect 25041 20751 25099 20757
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 2225 20587 2283 20593
rect 2225 20553 2237 20587
rect 2271 20584 2283 20587
rect 4982 20584 4988 20596
rect 2271 20556 4988 20584
rect 2271 20553 2283 20556
rect 2225 20547 2283 20553
rect 4982 20544 4988 20556
rect 5040 20544 5046 20596
rect 5077 20587 5135 20593
rect 5077 20553 5089 20587
rect 5123 20584 5135 20587
rect 5166 20584 5172 20596
rect 5123 20556 5172 20584
rect 5123 20553 5135 20556
rect 5077 20547 5135 20553
rect 5166 20544 5172 20556
rect 5224 20544 5230 20596
rect 7745 20587 7803 20593
rect 7745 20553 7757 20587
rect 7791 20584 7803 20587
rect 10318 20584 10324 20596
rect 7791 20556 10324 20584
rect 7791 20553 7803 20556
rect 7745 20547 7803 20553
rect 10318 20544 10324 20556
rect 10376 20544 10382 20596
rect 10962 20544 10968 20596
rect 11020 20584 11026 20596
rect 12069 20587 12127 20593
rect 12069 20584 12081 20587
rect 11020 20556 12081 20584
rect 11020 20544 11026 20556
rect 12069 20553 12081 20556
rect 12115 20553 12127 20587
rect 12069 20547 12127 20553
rect 12434 20544 12440 20596
rect 12492 20544 12498 20596
rect 12526 20544 12532 20596
rect 12584 20544 12590 20596
rect 12710 20544 12716 20596
rect 12768 20584 12774 20596
rect 17586 20584 17592 20596
rect 12768 20556 17592 20584
rect 12768 20544 12774 20556
rect 17586 20544 17592 20556
rect 17644 20544 17650 20596
rect 18690 20544 18696 20596
rect 18748 20544 18754 20596
rect 20254 20584 20260 20596
rect 19904 20556 20260 20584
rect 1780 20488 2774 20516
rect 1780 20457 1808 20488
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20417 1823 20451
rect 1765 20411 1823 20417
rect 2409 20451 2467 20457
rect 2409 20417 2421 20451
rect 2455 20417 2467 20451
rect 2409 20411 2467 20417
rect 1578 20204 1584 20256
rect 1636 20204 1642 20256
rect 2424 20244 2452 20411
rect 2746 20312 2774 20488
rect 4706 20476 4712 20528
rect 4764 20516 4770 20528
rect 4893 20519 4951 20525
rect 4893 20516 4905 20519
rect 4764 20488 4905 20516
rect 4764 20476 4770 20488
rect 4893 20485 4905 20488
rect 4939 20516 4951 20519
rect 5258 20516 5264 20528
rect 4939 20488 5264 20516
rect 4939 20485 4951 20488
rect 4893 20479 4951 20485
rect 5258 20476 5264 20488
rect 5316 20476 5322 20528
rect 11149 20519 11207 20525
rect 11149 20516 11161 20519
rect 10534 20488 11161 20516
rect 11149 20485 11161 20488
rect 11195 20516 11207 20519
rect 11422 20516 11428 20528
rect 11195 20488 11428 20516
rect 11195 20485 11207 20488
rect 11149 20479 11207 20485
rect 11422 20476 11428 20488
rect 11480 20516 11486 20528
rect 12158 20516 12164 20528
rect 11480 20488 12164 20516
rect 11480 20476 11486 20488
rect 12158 20476 12164 20488
rect 12216 20516 12222 20528
rect 13081 20519 13139 20525
rect 13081 20516 13093 20519
rect 12216 20488 13093 20516
rect 12216 20476 12222 20488
rect 13081 20485 13093 20488
rect 13127 20516 13139 20519
rect 13538 20516 13544 20528
rect 13127 20488 13544 20516
rect 13127 20485 13139 20488
rect 13081 20479 13139 20485
rect 13538 20476 13544 20488
rect 13596 20516 13602 20528
rect 18506 20516 18512 20528
rect 13596 20488 14306 20516
rect 18446 20488 18512 20516
rect 13596 20476 13602 20488
rect 18506 20476 18512 20488
rect 18564 20516 18570 20528
rect 19150 20516 19156 20528
rect 18564 20488 19156 20516
rect 18564 20476 18570 20488
rect 19150 20476 19156 20488
rect 19208 20516 19214 20528
rect 19904 20516 19932 20556
rect 20254 20544 20260 20556
rect 20312 20544 20318 20596
rect 20806 20544 20812 20596
rect 20864 20584 20870 20596
rect 20993 20587 21051 20593
rect 20993 20584 21005 20587
rect 20864 20556 21005 20584
rect 20864 20544 20870 20556
rect 20993 20553 21005 20556
rect 21039 20553 21051 20587
rect 20993 20547 21051 20553
rect 22097 20587 22155 20593
rect 22097 20553 22109 20587
rect 22143 20584 22155 20587
rect 23658 20584 23664 20596
rect 22143 20556 23664 20584
rect 22143 20553 22155 20556
rect 22097 20547 22155 20553
rect 23658 20544 23664 20556
rect 23716 20544 23722 20596
rect 19208 20488 20010 20516
rect 19208 20476 19214 20488
rect 22186 20476 22192 20528
rect 22244 20516 22250 20528
rect 22465 20519 22523 20525
rect 22465 20516 22477 20519
rect 22244 20488 22477 20516
rect 22244 20476 22250 20488
rect 22465 20485 22477 20488
rect 22511 20516 22523 20519
rect 22554 20516 22560 20528
rect 22511 20488 22560 20516
rect 22511 20485 22523 20488
rect 22465 20479 22523 20485
rect 22554 20476 22560 20488
rect 22612 20476 22618 20528
rect 22738 20476 22744 20528
rect 22796 20516 22802 20528
rect 23750 20516 23756 20528
rect 22796 20488 23756 20516
rect 22796 20476 22802 20488
rect 23750 20476 23756 20488
rect 23808 20476 23814 20528
rect 25222 20516 25228 20528
rect 24978 20488 25228 20516
rect 25222 20476 25228 20488
rect 25280 20476 25286 20528
rect 3053 20451 3111 20457
rect 3053 20417 3065 20451
rect 3099 20448 3111 20451
rect 5534 20448 5540 20460
rect 3099 20420 5540 20448
rect 3099 20417 3111 20420
rect 3053 20411 3111 20417
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 5997 20451 6055 20457
rect 5997 20417 6009 20451
rect 6043 20448 6055 20451
rect 7190 20448 7196 20460
rect 6043 20420 7196 20448
rect 6043 20417 6055 20420
rect 5997 20411 6055 20417
rect 7190 20408 7196 20420
rect 7248 20408 7254 20460
rect 7282 20408 7288 20460
rect 7340 20408 7346 20460
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20417 8631 20451
rect 8573 20411 8631 20417
rect 3326 20340 3332 20392
rect 3384 20340 3390 20392
rect 8588 20380 8616 20411
rect 9030 20408 9036 20460
rect 9088 20408 9094 20460
rect 12802 20408 12808 20460
rect 12860 20448 12866 20460
rect 12860 20420 13032 20448
rect 12860 20408 12866 20420
rect 9309 20383 9367 20389
rect 8588 20352 9168 20380
rect 8846 20312 8852 20324
rect 2746 20284 8852 20312
rect 8846 20272 8852 20284
rect 8904 20272 8910 20324
rect 4062 20244 4068 20256
rect 2424 20216 4068 20244
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 4154 20204 4160 20256
rect 4212 20244 4218 20256
rect 5813 20247 5871 20253
rect 5813 20244 5825 20247
rect 4212 20216 5825 20244
rect 4212 20204 4218 20216
rect 5813 20213 5825 20216
rect 5859 20213 5871 20247
rect 5813 20207 5871 20213
rect 6086 20204 6092 20256
rect 6144 20244 6150 20256
rect 7101 20247 7159 20253
rect 7101 20244 7113 20247
rect 6144 20216 7113 20244
rect 6144 20204 6150 20216
rect 7101 20213 7113 20216
rect 7147 20213 7159 20247
rect 7101 20207 7159 20213
rect 8386 20204 8392 20256
rect 8444 20204 8450 20256
rect 9140 20244 9168 20352
rect 9309 20349 9321 20383
rect 9355 20380 9367 20383
rect 10042 20380 10048 20392
rect 9355 20352 10048 20380
rect 9355 20349 9367 20352
rect 9309 20343 9367 20349
rect 10042 20340 10048 20352
rect 10100 20340 10106 20392
rect 12621 20383 12679 20389
rect 12621 20349 12633 20383
rect 12667 20349 12679 20383
rect 12621 20343 12679 20349
rect 10704 20284 10916 20312
rect 10704 20244 10732 20284
rect 9140 20216 10732 20244
rect 10778 20204 10784 20256
rect 10836 20204 10842 20256
rect 10888 20244 10916 20284
rect 12434 20272 12440 20324
rect 12492 20312 12498 20324
rect 12636 20312 12664 20343
rect 12492 20284 12664 20312
rect 12492 20272 12498 20284
rect 13004 20244 13032 20420
rect 15838 20408 15844 20460
rect 15896 20408 15902 20460
rect 16482 20408 16488 20460
rect 16540 20448 16546 20460
rect 16945 20451 17003 20457
rect 16945 20448 16957 20451
rect 16540 20420 16957 20448
rect 16540 20408 16546 20420
rect 16945 20417 16957 20420
rect 16991 20417 17003 20451
rect 16945 20411 17003 20417
rect 23290 20408 23296 20460
rect 23348 20448 23354 20460
rect 23477 20451 23535 20457
rect 23477 20448 23489 20451
rect 23348 20420 23489 20448
rect 23348 20408 23354 20420
rect 23477 20417 23489 20420
rect 23523 20417 23535 20451
rect 23477 20411 23535 20417
rect 13541 20383 13599 20389
rect 13541 20349 13553 20383
rect 13587 20380 13599 20383
rect 13817 20383 13875 20389
rect 13587 20352 13676 20380
rect 13587 20349 13599 20352
rect 13541 20343 13599 20349
rect 10888 20216 13032 20244
rect 13648 20244 13676 20352
rect 13817 20349 13829 20383
rect 13863 20380 13875 20383
rect 17221 20383 17279 20389
rect 13863 20352 14964 20380
rect 13863 20349 13875 20352
rect 13817 20343 13875 20349
rect 14936 20312 14964 20352
rect 17221 20349 17233 20383
rect 17267 20380 17279 20383
rect 17678 20380 17684 20392
rect 17267 20352 17684 20380
rect 17267 20349 17279 20352
rect 17221 20343 17279 20349
rect 17678 20340 17684 20352
rect 17736 20340 17742 20392
rect 19242 20340 19248 20392
rect 19300 20340 19306 20392
rect 19521 20383 19579 20389
rect 19521 20349 19533 20383
rect 19567 20380 19579 20383
rect 19886 20380 19892 20392
rect 19567 20352 19892 20380
rect 19567 20349 19579 20352
rect 19521 20343 19579 20349
rect 19886 20340 19892 20352
rect 19944 20340 19950 20392
rect 21450 20340 21456 20392
rect 21508 20380 21514 20392
rect 22370 20380 22376 20392
rect 21508 20352 22376 20380
rect 21508 20340 21514 20352
rect 22370 20340 22376 20352
rect 22428 20340 22434 20392
rect 22554 20340 22560 20392
rect 22612 20340 22618 20392
rect 22646 20340 22652 20392
rect 22704 20340 22710 20392
rect 23201 20383 23259 20389
rect 23201 20349 23213 20383
rect 23247 20380 23259 20383
rect 23842 20380 23848 20392
rect 23247 20352 23848 20380
rect 23247 20349 23259 20352
rect 23201 20343 23259 20349
rect 16206 20312 16212 20324
rect 14936 20284 16212 20312
rect 16206 20272 16212 20284
rect 16264 20272 16270 20324
rect 21542 20272 21548 20324
rect 21600 20312 21606 20324
rect 22278 20312 22284 20324
rect 21600 20284 22284 20312
rect 21600 20272 21606 20284
rect 22278 20272 22284 20284
rect 22336 20272 22342 20324
rect 13814 20244 13820 20256
rect 13648 20216 13820 20244
rect 13814 20204 13820 20216
rect 13872 20244 13878 20256
rect 14274 20244 14280 20256
rect 13872 20216 14280 20244
rect 13872 20204 13878 20216
rect 14274 20204 14280 20216
rect 14332 20204 14338 20256
rect 15102 20204 15108 20256
rect 15160 20244 15166 20256
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 15160 20216 15301 20244
rect 15160 20204 15166 20216
rect 15289 20213 15301 20216
rect 15335 20213 15347 20247
rect 15289 20207 15347 20213
rect 15930 20204 15936 20256
rect 15988 20204 15994 20256
rect 16022 20204 16028 20256
rect 16080 20244 16086 20256
rect 16301 20247 16359 20253
rect 16301 20244 16313 20247
rect 16080 20216 16313 20244
rect 16080 20204 16086 20216
rect 16301 20213 16313 20216
rect 16347 20213 16359 20247
rect 16301 20207 16359 20213
rect 16390 20204 16396 20256
rect 16448 20244 16454 20256
rect 20806 20244 20812 20256
rect 16448 20216 20812 20244
rect 16448 20204 16454 20216
rect 20806 20204 20812 20216
rect 20864 20204 20870 20256
rect 21174 20204 21180 20256
rect 21232 20244 21238 20256
rect 21269 20247 21327 20253
rect 21269 20244 21281 20247
rect 21232 20216 21281 20244
rect 21232 20204 21238 20216
rect 21269 20213 21281 20216
rect 21315 20244 21327 20247
rect 21453 20247 21511 20253
rect 21453 20244 21465 20247
rect 21315 20216 21465 20244
rect 21315 20213 21327 20216
rect 21269 20207 21327 20213
rect 21453 20213 21465 20216
rect 21499 20244 21511 20247
rect 21818 20244 21824 20256
rect 21499 20216 21824 20244
rect 21499 20213 21511 20216
rect 21453 20207 21511 20213
rect 21818 20204 21824 20216
rect 21876 20244 21882 20256
rect 23216 20244 23244 20343
rect 23842 20340 23848 20352
rect 23900 20340 23906 20392
rect 21876 20216 23244 20244
rect 21876 20204 21882 20216
rect 25222 20204 25228 20256
rect 25280 20204 25286 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 1578 20000 1584 20052
rect 1636 20040 1642 20052
rect 1636 20012 2774 20040
rect 1636 20000 1642 20012
rect 2746 19972 2774 20012
rect 3970 20000 3976 20052
rect 4028 20040 4034 20052
rect 6730 20040 6736 20052
rect 4028 20012 6736 20040
rect 4028 20000 4034 20012
rect 6730 20000 6736 20012
rect 6788 20000 6794 20052
rect 7190 20000 7196 20052
rect 7248 20040 7254 20052
rect 10413 20043 10471 20049
rect 10413 20040 10425 20043
rect 7248 20012 10425 20040
rect 7248 20000 7254 20012
rect 10413 20009 10425 20012
rect 10459 20009 10471 20043
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 10413 20003 10471 20009
rect 10980 20012 14933 20040
rect 5074 19972 5080 19984
rect 2746 19944 5080 19972
rect 5074 19932 5080 19944
rect 5132 19932 5138 19984
rect 10980 19972 11008 20012
rect 14921 20009 14933 20012
rect 14967 20009 14979 20043
rect 14921 20003 14979 20009
rect 15286 20000 15292 20052
rect 15344 20040 15350 20052
rect 16942 20040 16948 20052
rect 15344 20012 16948 20040
rect 15344 20000 15350 20012
rect 16942 20000 16948 20012
rect 17000 20040 17006 20052
rect 17313 20043 17371 20049
rect 17313 20040 17325 20043
rect 17000 20012 17325 20040
rect 17000 20000 17006 20012
rect 17313 20009 17325 20012
rect 17359 20009 17371 20043
rect 17313 20003 17371 20009
rect 17586 20000 17592 20052
rect 17644 20040 17650 20052
rect 17681 20043 17739 20049
rect 17681 20040 17693 20043
rect 17644 20012 17693 20040
rect 17644 20000 17650 20012
rect 17681 20009 17693 20012
rect 17727 20009 17739 20043
rect 17681 20003 17739 20009
rect 18877 20043 18935 20049
rect 18877 20009 18889 20043
rect 18923 20040 18935 20043
rect 19150 20040 19156 20052
rect 18923 20012 19156 20040
rect 18923 20009 18935 20012
rect 18877 20003 18935 20009
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 20254 20000 20260 20052
rect 20312 20040 20318 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20312 20012 20729 20040
rect 20312 20000 20318 20012
rect 20717 20009 20729 20012
rect 20763 20040 20775 20043
rect 21082 20040 21088 20052
rect 20763 20012 21088 20040
rect 20763 20009 20775 20012
rect 20717 20003 20775 20009
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 21910 20000 21916 20052
rect 21968 20040 21974 20052
rect 22833 20043 22891 20049
rect 22833 20040 22845 20043
rect 21968 20012 22845 20040
rect 21968 20000 21974 20012
rect 22833 20009 22845 20012
rect 22879 20009 22891 20043
rect 22833 20003 22891 20009
rect 24581 20043 24639 20049
rect 24581 20009 24593 20043
rect 24627 20040 24639 20043
rect 24670 20040 24676 20052
rect 24627 20012 24676 20040
rect 24627 20009 24639 20012
rect 24581 20003 24639 20009
rect 24670 20000 24676 20012
rect 24728 20000 24734 20052
rect 6564 19944 10732 19972
rect 2038 19864 2044 19916
rect 2096 19904 2102 19916
rect 2501 19907 2559 19913
rect 2501 19904 2513 19907
rect 2096 19876 2513 19904
rect 2096 19864 2102 19876
rect 2501 19873 2513 19876
rect 2547 19873 2559 19907
rect 2501 19867 2559 19873
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19836 2283 19839
rect 2314 19836 2320 19848
rect 2271 19808 2320 19836
rect 2271 19805 2283 19808
rect 2225 19799 2283 19805
rect 2314 19796 2320 19808
rect 2372 19796 2378 19848
rect 4706 19796 4712 19848
rect 4764 19796 4770 19848
rect 5166 19796 5172 19848
rect 5224 19796 5230 19848
rect 5445 19839 5503 19845
rect 5445 19805 5457 19839
rect 5491 19805 5503 19839
rect 6564 19836 6592 19944
rect 6641 19839 6699 19845
rect 6641 19836 6653 19839
rect 6564 19808 6653 19836
rect 5445 19799 5503 19805
rect 6641 19805 6653 19808
rect 6687 19805 6699 19839
rect 6641 19799 6699 19805
rect 5460 19768 5488 19799
rect 6730 19796 6736 19848
rect 6788 19836 6794 19848
rect 7101 19839 7159 19845
rect 7101 19836 7113 19839
rect 6788 19808 7113 19836
rect 6788 19796 6794 19808
rect 7101 19805 7113 19808
rect 7147 19805 7159 19839
rect 7101 19799 7159 19805
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19836 7435 19839
rect 9490 19836 9496 19848
rect 7423 19808 9496 19836
rect 7423 19805 7435 19808
rect 7377 19799 7435 19805
rect 9490 19796 9496 19808
rect 9548 19796 9554 19848
rect 10704 19836 10732 19944
rect 10888 19944 11008 19972
rect 13357 19975 13415 19981
rect 10888 19913 10916 19944
rect 13357 19941 13369 19975
rect 13403 19972 13415 19975
rect 13446 19972 13452 19984
rect 13403 19944 13452 19972
rect 13403 19941 13415 19944
rect 13357 19935 13415 19941
rect 13446 19932 13452 19944
rect 13504 19932 13510 19984
rect 13538 19932 13544 19984
rect 13596 19972 13602 19984
rect 13633 19975 13691 19981
rect 13633 19972 13645 19975
rect 13596 19944 13645 19972
rect 13596 19932 13602 19944
rect 13633 19941 13645 19944
rect 13679 19972 13691 19975
rect 13817 19975 13875 19981
rect 13817 19972 13829 19975
rect 13679 19944 13829 19972
rect 13679 19941 13691 19944
rect 13633 19935 13691 19941
rect 13817 19941 13829 19944
rect 13863 19972 13875 19975
rect 14090 19972 14096 19984
rect 13863 19944 14096 19972
rect 13863 19941 13875 19944
rect 13817 19935 13875 19941
rect 14090 19932 14096 19944
rect 14148 19932 14154 19984
rect 14550 19932 14556 19984
rect 14608 19972 14614 19984
rect 16390 19972 16396 19984
rect 14608 19944 16396 19972
rect 14608 19932 14614 19944
rect 16390 19932 16396 19944
rect 16448 19932 16454 19984
rect 16853 19975 16911 19981
rect 16853 19941 16865 19975
rect 16899 19972 16911 19975
rect 18506 19972 18512 19984
rect 16899 19944 18512 19972
rect 16899 19941 16911 19944
rect 16853 19935 16911 19941
rect 18506 19932 18512 19944
rect 18564 19932 18570 19984
rect 18785 19975 18843 19981
rect 18785 19972 18797 19975
rect 18616 19944 18797 19972
rect 10873 19907 10931 19913
rect 10873 19873 10885 19907
rect 10919 19873 10931 19907
rect 10873 19867 10931 19873
rect 10962 19864 10968 19916
rect 11020 19864 11026 19916
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 11112 19876 15485 19904
rect 11112 19864 11118 19876
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 18233 19907 18291 19913
rect 18233 19904 18245 19907
rect 15473 19867 15531 19873
rect 15580 19876 18245 19904
rect 11238 19836 11244 19848
rect 10704 19808 11244 19836
rect 11238 19796 11244 19808
rect 11296 19796 11302 19848
rect 11606 19796 11612 19848
rect 11664 19796 11670 19848
rect 13906 19836 13912 19848
rect 13188 19808 13912 19836
rect 7834 19768 7840 19780
rect 5460 19740 7840 19768
rect 7834 19728 7840 19740
rect 7892 19728 7898 19780
rect 8389 19771 8447 19777
rect 8389 19737 8401 19771
rect 8435 19768 8447 19771
rect 10781 19771 10839 19777
rect 10781 19768 10793 19771
rect 8435 19740 10793 19768
rect 8435 19737 8447 19740
rect 8389 19731 8447 19737
rect 10781 19737 10793 19740
rect 10827 19737 10839 19771
rect 10781 19731 10839 19737
rect 11885 19771 11943 19777
rect 11885 19737 11897 19771
rect 11931 19737 11943 19771
rect 11885 19731 11943 19737
rect 4522 19660 4528 19712
rect 4580 19660 4586 19712
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 6457 19703 6515 19709
rect 6457 19700 6469 19703
rect 5592 19672 6469 19700
rect 5592 19660 5598 19672
rect 6457 19669 6469 19672
rect 6503 19669 6515 19703
rect 6457 19663 6515 19669
rect 6638 19660 6644 19712
rect 6696 19700 6702 19712
rect 8294 19700 8300 19712
rect 6696 19672 8300 19700
rect 6696 19660 6702 19672
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 9122 19660 9128 19712
rect 9180 19660 9186 19712
rect 9769 19703 9827 19709
rect 9769 19669 9781 19703
rect 9815 19700 9827 19703
rect 10870 19700 10876 19712
rect 9815 19672 10876 19700
rect 9815 19669 9827 19672
rect 9769 19663 9827 19669
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 11900 19700 11928 19731
rect 12158 19728 12164 19780
rect 12216 19768 12222 19780
rect 12216 19740 12374 19768
rect 12216 19728 12222 19740
rect 13188 19700 13216 19808
rect 13906 19796 13912 19808
rect 13964 19796 13970 19848
rect 14182 19796 14188 19848
rect 14240 19836 14246 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 14240 19808 14289 19836
rect 14240 19796 14246 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 15580 19836 15608 19876
rect 18233 19873 18245 19876
rect 18279 19873 18291 19907
rect 18233 19867 18291 19873
rect 14277 19799 14335 19805
rect 14384 19808 15608 19836
rect 13446 19728 13452 19780
rect 13504 19768 13510 19780
rect 14384 19768 14412 19808
rect 16942 19796 16948 19848
rect 17000 19836 17006 19848
rect 17037 19839 17095 19845
rect 17037 19836 17049 19839
rect 17000 19808 17049 19836
rect 17000 19796 17006 19808
rect 17037 19805 17049 19808
rect 17083 19805 17095 19839
rect 17037 19799 17095 19805
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19836 18199 19839
rect 18616 19836 18644 19944
rect 18785 19941 18797 19944
rect 18831 19972 18843 19975
rect 18966 19972 18972 19984
rect 18831 19944 18972 19972
rect 18831 19941 18843 19944
rect 18785 19935 18843 19941
rect 18966 19932 18972 19944
rect 19024 19932 19030 19984
rect 23566 19932 23572 19984
rect 23624 19972 23630 19984
rect 23624 19944 25176 19972
rect 23624 19932 23630 19944
rect 18690 19864 18696 19916
rect 18748 19904 18754 19916
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 18748 19876 19993 19904
rect 18748 19864 18754 19876
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 19981 19867 20039 19873
rect 21085 19907 21143 19913
rect 21085 19873 21097 19907
rect 21131 19904 21143 19907
rect 23290 19904 23296 19916
rect 21131 19876 23296 19904
rect 21131 19873 21143 19876
rect 21085 19867 21143 19873
rect 23290 19864 23296 19876
rect 23348 19864 23354 19916
rect 23937 19907 23995 19913
rect 23937 19873 23949 19907
rect 23983 19904 23995 19907
rect 24118 19904 24124 19916
rect 23983 19876 24124 19904
rect 23983 19873 23995 19876
rect 23937 19867 23995 19873
rect 24118 19864 24124 19876
rect 24176 19864 24182 19916
rect 25148 19913 25176 19944
rect 25133 19907 25191 19913
rect 25133 19873 25145 19907
rect 25179 19873 25191 19907
rect 25133 19867 25191 19873
rect 18187 19808 18644 19836
rect 18187 19805 18199 19808
rect 18141 19799 18199 19805
rect 22922 19796 22928 19848
rect 22980 19836 22986 19848
rect 25041 19839 25099 19845
rect 25041 19836 25053 19839
rect 22980 19808 25053 19836
rect 22980 19796 22986 19808
rect 25041 19805 25053 19808
rect 25087 19805 25099 19839
rect 25041 19799 25099 19805
rect 13504 19740 14412 19768
rect 13504 19728 13510 19740
rect 15194 19728 15200 19780
rect 15252 19768 15258 19780
rect 15381 19771 15439 19777
rect 15381 19768 15393 19771
rect 15252 19740 15393 19768
rect 15252 19728 15258 19740
rect 15381 19737 15393 19740
rect 15427 19737 15439 19771
rect 15381 19731 15439 19737
rect 16206 19728 16212 19780
rect 16264 19728 16270 19780
rect 16390 19728 16396 19780
rect 16448 19768 16454 19780
rect 19797 19771 19855 19777
rect 16448 19740 19472 19768
rect 16448 19728 16454 19740
rect 11900 19672 13216 19700
rect 15286 19660 15292 19712
rect 15344 19660 15350 19712
rect 16298 19660 16304 19712
rect 16356 19660 16362 19712
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 19444 19709 19472 19740
rect 19797 19737 19809 19771
rect 19843 19768 19855 19771
rect 20070 19768 20076 19780
rect 19843 19740 20076 19768
rect 19843 19737 19855 19740
rect 19797 19731 19855 19737
rect 20070 19728 20076 19740
rect 20128 19728 20134 19780
rect 21358 19728 21364 19780
rect 21416 19728 21422 19780
rect 21818 19728 21824 19780
rect 21876 19728 21882 19780
rect 23753 19771 23811 19777
rect 23753 19768 23765 19771
rect 23124 19740 23765 19768
rect 23124 19712 23152 19740
rect 23753 19737 23765 19740
rect 23799 19737 23811 19771
rect 23753 19731 23811 19737
rect 24949 19771 25007 19777
rect 24949 19737 24961 19771
rect 24995 19768 25007 19771
rect 26050 19768 26056 19780
rect 24995 19740 26056 19768
rect 24995 19737 25007 19740
rect 24949 19731 25007 19737
rect 26050 19728 26056 19740
rect 26108 19728 26114 19780
rect 18049 19703 18107 19709
rect 18049 19700 18061 19703
rect 16632 19672 18061 19700
rect 16632 19660 16638 19672
rect 18049 19669 18061 19672
rect 18095 19669 18107 19703
rect 18049 19663 18107 19669
rect 19429 19703 19487 19709
rect 19429 19669 19441 19703
rect 19475 19669 19487 19703
rect 19429 19663 19487 19669
rect 19610 19660 19616 19712
rect 19668 19700 19674 19712
rect 19889 19703 19947 19709
rect 19889 19700 19901 19703
rect 19668 19672 19901 19700
rect 19668 19660 19674 19672
rect 19889 19669 19901 19672
rect 19935 19669 19947 19703
rect 19889 19663 19947 19669
rect 20806 19660 20812 19712
rect 20864 19700 20870 19712
rect 23014 19700 23020 19712
rect 20864 19672 23020 19700
rect 20864 19660 20870 19672
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 23106 19660 23112 19712
rect 23164 19660 23170 19712
rect 23293 19703 23351 19709
rect 23293 19669 23305 19703
rect 23339 19700 23351 19703
rect 23382 19700 23388 19712
rect 23339 19672 23388 19700
rect 23339 19669 23351 19672
rect 23293 19663 23351 19669
rect 23382 19660 23388 19672
rect 23440 19660 23446 19712
rect 23474 19660 23480 19712
rect 23532 19700 23538 19712
rect 23661 19703 23719 19709
rect 23661 19700 23673 19703
rect 23532 19672 23673 19700
rect 23532 19660 23538 19672
rect 23661 19669 23673 19672
rect 23707 19669 23719 19703
rect 23661 19663 23719 19669
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 3878 19456 3884 19508
rect 3936 19456 3942 19508
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 5813 19499 5871 19505
rect 5813 19496 5825 19499
rect 5224 19468 5825 19496
rect 5224 19456 5230 19468
rect 5813 19465 5825 19468
rect 5859 19465 5871 19499
rect 5813 19459 5871 19465
rect 7101 19499 7159 19505
rect 7101 19465 7113 19499
rect 7147 19496 7159 19499
rect 9214 19496 9220 19508
rect 7147 19468 9220 19496
rect 7147 19465 7159 19468
rect 7101 19459 7159 19465
rect 9214 19456 9220 19468
rect 9272 19456 9278 19508
rect 10778 19496 10784 19508
rect 9324 19468 10784 19496
rect 8202 19428 8208 19440
rect 4080 19400 8208 19428
rect 1949 19363 2007 19369
rect 1949 19329 1961 19363
rect 1995 19360 2007 19363
rect 3602 19360 3608 19372
rect 1995 19332 3608 19360
rect 1995 19329 2007 19332
rect 1949 19323 2007 19329
rect 3602 19320 3608 19332
rect 3660 19320 3666 19372
rect 4080 19369 4108 19400
rect 8202 19388 8208 19400
rect 8260 19388 8266 19440
rect 9324 19437 9352 19468
rect 10778 19456 10784 19468
rect 10836 19456 10842 19508
rect 11057 19499 11115 19505
rect 11057 19465 11069 19499
rect 11103 19496 11115 19499
rect 11609 19499 11667 19505
rect 11609 19496 11621 19499
rect 11103 19468 11621 19496
rect 11103 19465 11115 19468
rect 11057 19459 11115 19465
rect 11609 19465 11621 19468
rect 11655 19496 11667 19499
rect 11701 19499 11759 19505
rect 11701 19496 11713 19499
rect 11655 19468 11713 19496
rect 11655 19465 11667 19468
rect 11609 19459 11667 19465
rect 11701 19465 11713 19468
rect 11747 19496 11759 19499
rect 12158 19496 12164 19508
rect 11747 19468 12164 19496
rect 11747 19465 11759 19468
rect 11701 19459 11759 19465
rect 9309 19431 9367 19437
rect 9309 19397 9321 19431
rect 9355 19397 9367 19431
rect 11072 19428 11100 19459
rect 12158 19456 12164 19468
rect 12216 19456 12222 19508
rect 13814 19496 13820 19508
rect 12544 19468 13820 19496
rect 10534 19400 11100 19428
rect 9309 19391 9367 19397
rect 4065 19363 4123 19369
rect 4065 19329 4077 19363
rect 4111 19329 4123 19363
rect 4065 19323 4123 19329
rect 4801 19363 4859 19369
rect 4801 19329 4813 19363
rect 4847 19360 4859 19363
rect 5442 19360 5448 19372
rect 4847 19332 5448 19360
rect 4847 19329 4859 19332
rect 4801 19323 4859 19329
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 5994 19320 6000 19372
rect 6052 19320 6058 19372
rect 7285 19363 7343 19369
rect 7285 19360 7297 19363
rect 6748 19332 7297 19360
rect 1670 19252 1676 19304
rect 1728 19292 1734 19304
rect 2225 19295 2283 19301
rect 2225 19292 2237 19295
rect 1728 19264 2237 19292
rect 1728 19252 1734 19264
rect 2225 19261 2237 19264
rect 2271 19261 2283 19295
rect 2225 19255 2283 19261
rect 4522 19252 4528 19304
rect 4580 19252 4586 19304
rect 6454 19252 6460 19304
rect 6512 19252 6518 19304
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19292 6699 19295
rect 6748 19292 6776 19332
rect 7285 19329 7297 19332
rect 7331 19360 7343 19363
rect 7558 19360 7564 19372
rect 7331 19332 7564 19360
rect 7331 19329 7343 19332
rect 7285 19323 7343 19329
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 7834 19320 7840 19372
rect 7892 19360 7898 19372
rect 7929 19363 7987 19369
rect 7929 19360 7941 19363
rect 7892 19332 7941 19360
rect 7892 19320 7898 19332
rect 7929 19329 7941 19332
rect 7975 19329 7987 19363
rect 7929 19323 7987 19329
rect 8294 19320 8300 19372
rect 8352 19360 8358 19372
rect 8352 19332 8432 19360
rect 8352 19320 8358 19332
rect 6687 19264 6776 19292
rect 6825 19295 6883 19301
rect 6687 19261 6699 19264
rect 6641 19255 6699 19261
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 7098 19292 7104 19304
rect 6871 19264 7104 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 7098 19252 7104 19264
rect 7156 19252 7162 19304
rect 6914 19184 6920 19236
rect 6972 19224 6978 19236
rect 8404 19233 8432 19332
rect 8570 19320 8576 19372
rect 8628 19320 8634 19372
rect 9030 19320 9036 19372
rect 9088 19320 9094 19372
rect 11606 19320 11612 19372
rect 11664 19360 11670 19372
rect 12544 19360 12572 19468
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 13906 19456 13912 19508
rect 13964 19496 13970 19508
rect 14458 19496 14464 19508
rect 13964 19468 14464 19496
rect 13964 19456 13970 19468
rect 14458 19456 14464 19468
rect 14516 19456 14522 19508
rect 14826 19456 14832 19508
rect 14884 19496 14890 19508
rect 14921 19499 14979 19505
rect 14921 19496 14933 19499
rect 14884 19468 14933 19496
rect 14884 19456 14890 19468
rect 14921 19465 14933 19468
rect 14967 19465 14979 19499
rect 14921 19459 14979 19465
rect 15289 19499 15347 19505
rect 15289 19465 15301 19499
rect 15335 19496 15347 19499
rect 16390 19496 16396 19508
rect 15335 19468 16396 19496
rect 15335 19465 15347 19468
rect 15289 19459 15347 19465
rect 16390 19456 16396 19468
rect 16448 19456 16454 19508
rect 18690 19496 18696 19508
rect 16500 19468 18696 19496
rect 13538 19388 13544 19440
rect 13596 19388 13602 19440
rect 14274 19388 14280 19440
rect 14332 19428 14338 19440
rect 15381 19431 15439 19437
rect 15381 19428 15393 19431
rect 14332 19400 15393 19428
rect 14332 19388 14338 19400
rect 15381 19397 15393 19400
rect 15427 19397 15439 19431
rect 16500 19428 16528 19468
rect 18690 19456 18696 19468
rect 18748 19456 18754 19508
rect 18785 19499 18843 19505
rect 18785 19465 18797 19499
rect 18831 19465 18843 19499
rect 18785 19459 18843 19465
rect 19613 19499 19671 19505
rect 19613 19465 19625 19499
rect 19659 19496 19671 19499
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 19659 19468 20453 19496
rect 19659 19465 19671 19468
rect 19613 19459 19671 19465
rect 20441 19465 20453 19468
rect 20487 19465 20499 19499
rect 20441 19459 20499 19465
rect 20809 19499 20867 19505
rect 20809 19465 20821 19499
rect 20855 19496 20867 19499
rect 20855 19468 21220 19496
rect 20855 19465 20867 19468
rect 20809 19459 20867 19465
rect 15381 19391 15439 19397
rect 15488 19400 16528 19428
rect 18800 19428 18828 19459
rect 19886 19428 19892 19440
rect 18800 19400 19892 19428
rect 12713 19363 12771 19369
rect 12713 19360 12725 19363
rect 11664 19332 12725 19360
rect 11664 19320 11670 19332
rect 12713 19329 12725 19332
rect 12759 19329 12771 19363
rect 12713 19323 12771 19329
rect 14918 19320 14924 19372
rect 14976 19360 14982 19372
rect 15488 19360 15516 19400
rect 19886 19388 19892 19400
rect 19944 19388 19950 19440
rect 20901 19431 20959 19437
rect 20901 19397 20913 19431
rect 20947 19428 20959 19431
rect 20990 19428 20996 19440
rect 20947 19400 20996 19428
rect 20947 19397 20959 19400
rect 20901 19391 20959 19397
rect 20990 19388 20996 19400
rect 21048 19428 21054 19440
rect 21048 19400 21128 19428
rect 21048 19388 21054 19400
rect 14976 19332 15516 19360
rect 16301 19363 16359 19369
rect 14976 19320 14982 19332
rect 16301 19329 16313 19363
rect 16347 19360 16359 19363
rect 16347 19332 16436 19360
rect 16347 19329 16359 19332
rect 16301 19323 16359 19329
rect 9398 19252 9404 19304
rect 9456 19292 9462 19304
rect 11974 19292 11980 19304
rect 9456 19264 11980 19292
rect 9456 19252 9462 19264
rect 11974 19252 11980 19264
rect 12032 19252 12038 19304
rect 12066 19252 12072 19304
rect 12124 19252 12130 19304
rect 12989 19295 13047 19301
rect 12989 19261 13001 19295
rect 13035 19292 13047 19295
rect 15102 19292 15108 19304
rect 13035 19264 15108 19292
rect 13035 19261 13047 19264
rect 12989 19255 13047 19261
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 16022 19292 16028 19304
rect 15611 19264 16028 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 16408 19292 16436 19332
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 16540 19332 17049 19360
rect 16540 19320 16546 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 19150 19360 19156 19372
rect 18380 19332 19156 19360
rect 18380 19320 18386 19332
rect 19150 19320 19156 19332
rect 19208 19320 19214 19372
rect 19702 19320 19708 19372
rect 19760 19320 19766 19372
rect 16758 19292 16764 19304
rect 16408 19264 16764 19292
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 17310 19252 17316 19304
rect 17368 19292 17374 19304
rect 17368 19264 19840 19292
rect 17368 19252 17374 19264
rect 7745 19227 7803 19233
rect 7745 19224 7757 19227
rect 6972 19196 7757 19224
rect 6972 19184 6978 19196
rect 7745 19193 7757 19196
rect 7791 19193 7803 19227
rect 7745 19187 7803 19193
rect 8389 19227 8447 19233
rect 8389 19193 8401 19227
rect 8435 19193 8447 19227
rect 12158 19224 12164 19236
rect 8389 19187 8447 19193
rect 10336 19196 12164 19224
rect 2866 19116 2872 19168
rect 2924 19156 2930 19168
rect 10336 19156 10364 19196
rect 12158 19184 12164 19196
rect 12216 19184 12222 19236
rect 19702 19224 19708 19236
rect 18340 19196 19708 19224
rect 2924 19128 10364 19156
rect 2924 19116 2930 19128
rect 10778 19116 10784 19168
rect 10836 19156 10842 19168
rect 10962 19156 10968 19168
rect 10836 19128 10968 19156
rect 10836 19116 10842 19128
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 11146 19116 11152 19168
rect 11204 19156 11210 19168
rect 11241 19159 11299 19165
rect 11241 19156 11253 19159
rect 11204 19128 11253 19156
rect 11204 19116 11210 19128
rect 11241 19125 11253 19128
rect 11287 19125 11299 19159
rect 11241 19119 11299 19125
rect 12250 19116 12256 19168
rect 12308 19156 12314 19168
rect 13446 19156 13452 19168
rect 12308 19128 13452 19156
rect 12308 19116 12314 19128
rect 13446 19116 13452 19128
rect 13504 19116 13510 19168
rect 16117 19159 16175 19165
rect 16117 19125 16129 19159
rect 16163 19156 16175 19159
rect 16298 19156 16304 19168
rect 16163 19128 16304 19156
rect 16163 19125 16175 19128
rect 16117 19119 16175 19125
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 18340 19156 18368 19196
rect 19702 19184 19708 19196
rect 19760 19184 19766 19236
rect 19812 19224 19840 19264
rect 19886 19252 19892 19304
rect 19944 19252 19950 19304
rect 20993 19295 21051 19301
rect 20993 19261 21005 19295
rect 21039 19261 21051 19295
rect 21100 19292 21128 19400
rect 21192 19360 21220 19468
rect 21818 19456 21824 19508
rect 21876 19496 21882 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21876 19468 22017 19496
rect 21876 19456 21882 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 22186 19456 22192 19508
rect 22244 19496 22250 19508
rect 22373 19499 22431 19505
rect 22373 19496 22385 19499
rect 22244 19468 22385 19496
rect 22244 19456 22250 19468
rect 22373 19465 22385 19468
rect 22419 19465 22431 19499
rect 22373 19459 22431 19465
rect 22462 19456 22468 19508
rect 22520 19456 22526 19508
rect 23934 19456 23940 19508
rect 23992 19456 23998 19508
rect 25038 19456 25044 19508
rect 25096 19456 25102 19508
rect 21358 19388 21364 19440
rect 21416 19428 21422 19440
rect 23842 19428 23848 19440
rect 21416 19400 23848 19428
rect 21416 19388 21422 19400
rect 23842 19388 23848 19400
rect 23900 19388 23906 19440
rect 23952 19428 23980 19456
rect 23952 19400 24058 19428
rect 22278 19360 22284 19372
rect 21192 19332 22284 19360
rect 22278 19320 22284 19332
rect 22336 19320 22342 19372
rect 22922 19360 22928 19372
rect 22480 19332 22928 19360
rect 21542 19292 21548 19304
rect 21100 19264 21548 19292
rect 20993 19255 21051 19261
rect 21008 19224 21036 19255
rect 21542 19252 21548 19264
rect 21600 19292 21606 19304
rect 22480 19292 22508 19332
rect 22922 19320 22928 19332
rect 22980 19320 22986 19372
rect 23290 19320 23296 19372
rect 23348 19320 23354 19372
rect 21600 19264 22508 19292
rect 22557 19295 22615 19301
rect 21600 19252 21606 19264
rect 22557 19261 22569 19295
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 23569 19295 23627 19301
rect 23569 19261 23581 19295
rect 23615 19292 23627 19295
rect 25222 19292 25228 19304
rect 23615 19264 25228 19292
rect 23615 19261 23627 19264
rect 23569 19255 23627 19261
rect 19812 19196 21036 19224
rect 21818 19184 21824 19236
rect 21876 19224 21882 19236
rect 22572 19224 22600 19255
rect 25222 19252 25228 19264
rect 25280 19252 25286 19304
rect 25314 19252 25320 19304
rect 25372 19252 25378 19304
rect 21876 19196 22600 19224
rect 21876 19184 21882 19196
rect 16448 19128 18368 19156
rect 16448 19116 16454 19128
rect 19150 19116 19156 19168
rect 19208 19156 19214 19168
rect 19245 19159 19303 19165
rect 19245 19156 19257 19159
rect 19208 19128 19257 19156
rect 19208 19116 19214 19128
rect 19245 19125 19257 19128
rect 19291 19125 19303 19159
rect 19245 19119 19303 19125
rect 21082 19116 21088 19168
rect 21140 19156 21146 19168
rect 21545 19159 21603 19165
rect 21545 19156 21557 19159
rect 21140 19128 21557 19156
rect 21140 19116 21146 19128
rect 21545 19125 21557 19128
rect 21591 19125 21603 19159
rect 21545 19119 21603 19125
rect 21726 19116 21732 19168
rect 21784 19156 21790 19168
rect 23382 19156 23388 19168
rect 21784 19128 23388 19156
rect 21784 19116 21790 19128
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 1946 18912 1952 18964
rect 2004 18912 2010 18964
rect 3694 18912 3700 18964
rect 3752 18952 3758 18964
rect 3789 18955 3847 18961
rect 3789 18952 3801 18955
rect 3752 18924 3801 18952
rect 3752 18912 3758 18924
rect 3789 18921 3801 18924
rect 3835 18921 3847 18955
rect 3789 18915 3847 18921
rect 4249 18955 4307 18961
rect 4249 18921 4261 18955
rect 4295 18952 4307 18955
rect 4798 18952 4804 18964
rect 4295 18924 4804 18952
rect 4295 18921 4307 18924
rect 4249 18915 4307 18921
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 5813 18955 5871 18961
rect 5813 18921 5825 18955
rect 5859 18952 5871 18955
rect 5902 18952 5908 18964
rect 5859 18924 5908 18952
rect 5859 18921 5871 18924
rect 5813 18915 5871 18921
rect 5902 18912 5908 18924
rect 5960 18912 5966 18964
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 8389 18955 8447 18961
rect 8389 18952 8401 18955
rect 8260 18924 8401 18952
rect 8260 18912 8266 18924
rect 8389 18921 8401 18924
rect 8435 18921 8447 18955
rect 8389 18915 8447 18921
rect 8846 18912 8852 18964
rect 8904 18952 8910 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 8904 18924 9229 18952
rect 8904 18912 8910 18924
rect 9217 18921 9229 18924
rect 9263 18921 9275 18955
rect 9217 18915 9275 18921
rect 9766 18912 9772 18964
rect 9824 18952 9830 18964
rect 10318 18952 10324 18964
rect 9824 18924 10324 18952
rect 9824 18912 9830 18924
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 11238 18912 11244 18964
rect 11296 18952 11302 18964
rect 12989 18955 13047 18961
rect 12989 18952 13001 18955
rect 11296 18924 13001 18952
rect 11296 18912 11302 18924
rect 12989 18921 13001 18924
rect 13035 18921 13047 18955
rect 12989 18915 13047 18921
rect 14274 18912 14280 18964
rect 14332 18912 14338 18964
rect 15470 18952 15476 18964
rect 14752 18924 15476 18952
rect 2593 18887 2651 18893
rect 2593 18853 2605 18887
rect 2639 18884 2651 18887
rect 2639 18856 3832 18884
rect 2639 18853 2651 18856
rect 2593 18847 2651 18853
rect 3694 18816 3700 18828
rect 2792 18788 3700 18816
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 2130 18748 2136 18760
rect 1719 18720 2136 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 2792 18757 2820 18788
rect 3694 18776 3700 18788
rect 3752 18776 3758 18828
rect 3804 18816 3832 18856
rect 4062 18844 4068 18896
rect 4120 18884 4126 18896
rect 4120 18856 9904 18884
rect 4120 18844 4126 18856
rect 7377 18819 7435 18825
rect 3804 18788 5488 18816
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18717 2835 18751
rect 2777 18711 2835 18717
rect 3421 18751 3479 18757
rect 3421 18717 3433 18751
rect 3467 18748 3479 18751
rect 4154 18748 4160 18760
rect 3467 18720 4160 18748
rect 3467 18717 3479 18720
rect 3421 18711 3479 18717
rect 4154 18708 4160 18720
rect 4212 18708 4218 18760
rect 4706 18708 4712 18760
rect 4764 18708 4770 18760
rect 4798 18708 4804 18760
rect 4856 18748 4862 18760
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 4856 18720 5365 18748
rect 4856 18708 4862 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 5258 18680 5264 18692
rect 3252 18652 5264 18680
rect 3252 18621 3280 18652
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 5460 18680 5488 18788
rect 7377 18785 7389 18819
rect 7423 18816 7435 18819
rect 7466 18816 7472 18828
rect 7423 18788 7472 18816
rect 7423 18785 7435 18788
rect 7377 18779 7435 18785
rect 7466 18776 7472 18788
rect 7524 18776 7530 18828
rect 8294 18776 8300 18828
rect 8352 18816 8358 18828
rect 8754 18816 8760 18828
rect 8352 18788 8760 18816
rect 8352 18776 8358 18788
rect 8754 18776 8760 18788
rect 8812 18776 8818 18828
rect 9398 18816 9404 18828
rect 8864 18788 9404 18816
rect 5994 18708 6000 18760
rect 6052 18708 6058 18760
rect 6454 18708 6460 18760
rect 6512 18748 6518 18760
rect 6641 18751 6699 18757
rect 6641 18748 6653 18751
rect 6512 18720 6653 18748
rect 6512 18708 6518 18720
rect 6641 18717 6653 18720
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 8386 18748 8392 18760
rect 7147 18720 8392 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 8386 18708 8392 18720
rect 8444 18708 8450 18760
rect 8570 18708 8576 18760
rect 8628 18708 8634 18760
rect 8864 18748 8892 18788
rect 9398 18776 9404 18788
rect 9456 18776 9462 18828
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 9769 18819 9827 18825
rect 9769 18816 9781 18819
rect 9548 18788 9781 18816
rect 9548 18776 9554 18788
rect 9769 18785 9781 18788
rect 9815 18785 9827 18819
rect 9876 18816 9904 18856
rect 11146 18844 11152 18896
rect 11204 18884 11210 18896
rect 12342 18884 12348 18896
rect 11204 18856 12348 18884
rect 11204 18844 11210 18856
rect 12342 18844 12348 18856
rect 12400 18844 12406 18896
rect 13464 18856 14688 18884
rect 13354 18816 13360 18828
rect 9876 18788 13360 18816
rect 9769 18779 9827 18785
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 8680 18720 8892 18748
rect 8680 18680 8708 18720
rect 9122 18708 9128 18760
rect 9180 18748 9186 18760
rect 9585 18751 9643 18757
rect 9585 18748 9597 18751
rect 9180 18720 9597 18748
rect 9180 18708 9186 18720
rect 9585 18717 9597 18720
rect 9631 18717 9643 18751
rect 11974 18748 11980 18760
rect 9585 18711 9643 18717
rect 10336 18720 11980 18748
rect 5460 18652 8708 18680
rect 8754 18640 8760 18692
rect 8812 18680 8818 18692
rect 10336 18680 10364 18720
rect 11974 18708 11980 18720
rect 12032 18708 12038 18760
rect 12158 18708 12164 18760
rect 12216 18748 12222 18760
rect 12434 18748 12440 18760
rect 12216 18720 12440 18748
rect 12216 18708 12222 18720
rect 12434 18708 12440 18720
rect 12492 18708 12498 18760
rect 13464 18757 13492 18856
rect 13633 18819 13691 18825
rect 13633 18785 13645 18819
rect 13679 18816 13691 18819
rect 13679 18788 14596 18816
rect 13679 18785 13691 18788
rect 13633 18779 13691 18785
rect 13449 18751 13507 18757
rect 13449 18717 13461 18751
rect 13495 18717 13507 18751
rect 13449 18711 13507 18717
rect 8812 18652 10364 18680
rect 10413 18683 10471 18689
rect 8812 18640 8818 18652
rect 10413 18649 10425 18683
rect 10459 18680 10471 18683
rect 12986 18680 12992 18692
rect 10459 18652 12992 18680
rect 10459 18649 10471 18652
rect 10413 18643 10471 18649
rect 12986 18640 12992 18652
rect 13044 18640 13050 18692
rect 13357 18683 13415 18689
rect 13357 18649 13369 18683
rect 13403 18680 13415 18683
rect 13722 18680 13728 18692
rect 13403 18652 13728 18680
rect 13403 18649 13415 18652
rect 13357 18643 13415 18649
rect 13722 18640 13728 18652
rect 13780 18640 13786 18692
rect 3237 18615 3295 18621
rect 3237 18581 3249 18615
rect 3283 18581 3295 18615
rect 3237 18575 3295 18581
rect 4525 18615 4583 18621
rect 4525 18581 4537 18615
rect 4571 18612 4583 18615
rect 4982 18612 4988 18624
rect 4571 18584 4988 18612
rect 4571 18581 4583 18584
rect 4525 18575 4583 18581
rect 4982 18572 4988 18584
rect 5040 18572 5046 18624
rect 5166 18572 5172 18624
rect 5224 18572 5230 18624
rect 6454 18572 6460 18624
rect 6512 18572 6518 18624
rect 6638 18572 6644 18624
rect 6696 18612 6702 18624
rect 9306 18612 9312 18624
rect 6696 18584 9312 18612
rect 6696 18572 6702 18584
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 9677 18615 9735 18621
rect 9677 18581 9689 18615
rect 9723 18612 9735 18615
rect 11698 18612 11704 18624
rect 9723 18584 11704 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 11882 18572 11888 18624
rect 11940 18572 11946 18624
rect 11974 18572 11980 18624
rect 12032 18612 12038 18624
rect 14458 18612 14464 18624
rect 12032 18584 14464 18612
rect 12032 18572 12038 18584
rect 14458 18572 14464 18584
rect 14516 18572 14522 18624
rect 14568 18612 14596 18788
rect 14660 18748 14688 18856
rect 14752 18825 14780 18924
rect 15470 18912 15476 18924
rect 15528 18952 15534 18964
rect 15746 18952 15752 18964
rect 15528 18924 15752 18952
rect 15528 18912 15534 18924
rect 15746 18912 15752 18924
rect 15804 18912 15810 18964
rect 17218 18912 17224 18964
rect 17276 18952 17282 18964
rect 17681 18955 17739 18961
rect 17681 18952 17693 18955
rect 17276 18924 17693 18952
rect 17276 18912 17282 18924
rect 17681 18921 17693 18924
rect 17727 18952 17739 18955
rect 17862 18952 17868 18964
rect 17727 18924 17868 18952
rect 17727 18921 17739 18924
rect 17681 18915 17739 18921
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 21358 18952 21364 18964
rect 20772 18924 21364 18952
rect 20772 18912 20778 18924
rect 21358 18912 21364 18924
rect 21416 18912 21422 18964
rect 22830 18912 22836 18964
rect 22888 18952 22894 18964
rect 23014 18952 23020 18964
rect 22888 18924 23020 18952
rect 22888 18912 22894 18924
rect 23014 18912 23020 18924
rect 23072 18912 23078 18964
rect 16850 18844 16856 18896
rect 16908 18884 16914 18896
rect 17770 18884 17776 18896
rect 16908 18856 17776 18884
rect 16908 18844 16914 18856
rect 17770 18844 17776 18856
rect 17828 18844 17834 18896
rect 18046 18844 18052 18896
rect 18104 18844 18110 18896
rect 18414 18844 18420 18896
rect 18472 18884 18478 18896
rect 18472 18856 18644 18884
rect 18472 18844 18478 18856
rect 14737 18819 14795 18825
rect 14737 18785 14749 18819
rect 14783 18785 14795 18819
rect 14737 18779 14795 18785
rect 14918 18776 14924 18828
rect 14976 18776 14982 18828
rect 15470 18776 15476 18828
rect 15528 18816 15534 18828
rect 16482 18816 16488 18828
rect 15528 18788 16488 18816
rect 15528 18776 15534 18788
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 17221 18819 17279 18825
rect 17221 18785 17233 18819
rect 17267 18816 17279 18819
rect 17678 18816 17684 18828
rect 17267 18788 17684 18816
rect 17267 18785 17279 18788
rect 17221 18779 17279 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 18322 18776 18328 18828
rect 18380 18816 18386 18828
rect 18380 18788 18460 18816
rect 18380 18776 18386 18788
rect 14660 18720 15516 18748
rect 14645 18683 14703 18689
rect 14645 18649 14657 18683
rect 14691 18680 14703 18683
rect 15286 18680 15292 18692
rect 14691 18652 15292 18680
rect 14691 18649 14703 18652
rect 14645 18643 14703 18649
rect 15286 18640 15292 18652
rect 15344 18640 15350 18692
rect 15194 18612 15200 18624
rect 14568 18584 15200 18612
rect 15194 18572 15200 18584
rect 15252 18572 15258 18624
rect 15488 18612 15516 18720
rect 17494 18708 17500 18760
rect 17552 18748 17558 18760
rect 18432 18748 18460 18788
rect 18506 18776 18512 18828
rect 18564 18776 18570 18828
rect 18616 18825 18644 18856
rect 22278 18844 22284 18896
rect 22336 18884 22342 18896
rect 22336 18856 23796 18884
rect 22336 18844 22342 18856
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 19116 18788 19441 18816
rect 19116 18776 19122 18788
rect 19429 18785 19441 18788
rect 19475 18785 19487 18819
rect 19429 18779 19487 18785
rect 20625 18819 20683 18825
rect 20625 18785 20637 18819
rect 20671 18816 20683 18819
rect 21910 18816 21916 18828
rect 20671 18788 21916 18816
rect 20671 18785 20683 18788
rect 20625 18779 20683 18785
rect 21910 18776 21916 18788
rect 21968 18776 21974 18828
rect 22830 18776 22836 18828
rect 22888 18816 22894 18828
rect 23768 18825 23796 18856
rect 23109 18819 23167 18825
rect 23109 18816 23121 18819
rect 22888 18788 23121 18816
rect 22888 18776 22894 18788
rect 23109 18785 23121 18788
rect 23155 18785 23167 18819
rect 23109 18779 23167 18785
rect 23753 18819 23811 18825
rect 23753 18785 23765 18819
rect 23799 18785 23811 18819
rect 23753 18779 23811 18785
rect 25222 18776 25228 18828
rect 25280 18776 25286 18828
rect 19242 18748 19248 18760
rect 17552 18720 18368 18748
rect 18432 18720 19248 18748
rect 17552 18708 17558 18720
rect 15749 18683 15807 18689
rect 15749 18649 15761 18683
rect 15795 18680 15807 18683
rect 16022 18680 16028 18692
rect 15795 18652 16028 18680
rect 15795 18649 15807 18652
rect 15749 18643 15807 18649
rect 16022 18640 16028 18652
rect 16080 18640 16086 18692
rect 16206 18640 16212 18692
rect 16264 18640 16270 18692
rect 18230 18680 18236 18692
rect 17512 18652 18236 18680
rect 17126 18612 17132 18624
rect 15488 18584 17132 18612
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 17218 18572 17224 18624
rect 17276 18612 17282 18624
rect 17512 18621 17540 18652
rect 18230 18640 18236 18652
rect 18288 18640 18294 18692
rect 18340 18680 18368 18720
rect 19242 18708 19248 18720
rect 19300 18748 19306 18760
rect 20349 18751 20407 18757
rect 20349 18748 20361 18751
rect 19300 18720 20361 18748
rect 19300 18708 19306 18720
rect 20349 18717 20361 18720
rect 20395 18717 20407 18751
rect 25041 18751 25099 18757
rect 25041 18748 25053 18751
rect 20349 18711 20407 18717
rect 22066 18720 25053 18748
rect 18506 18680 18512 18692
rect 18340 18652 18512 18680
rect 18506 18640 18512 18652
rect 18564 18640 18570 18692
rect 19518 18640 19524 18692
rect 19576 18680 19582 18692
rect 20254 18680 20260 18692
rect 19576 18652 20260 18680
rect 19576 18640 19582 18652
rect 20254 18640 20260 18652
rect 20312 18680 20318 18692
rect 20898 18680 20904 18692
rect 20312 18652 20904 18680
rect 20312 18640 20318 18652
rect 20898 18640 20904 18652
rect 20956 18640 20962 18692
rect 21082 18640 21088 18692
rect 21140 18640 21146 18692
rect 21910 18640 21916 18692
rect 21968 18680 21974 18692
rect 22066 18680 22094 18720
rect 25041 18717 25053 18720
rect 25087 18717 25099 18751
rect 25041 18711 25099 18717
rect 21968 18652 22094 18680
rect 21968 18640 21974 18652
rect 22922 18640 22928 18692
rect 22980 18640 22986 18692
rect 23014 18640 23020 18692
rect 23072 18640 23078 18692
rect 25222 18680 25228 18692
rect 24412 18652 25228 18680
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 17276 18584 17509 18612
rect 17276 18572 17282 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 17678 18572 17684 18624
rect 17736 18612 17742 18624
rect 17954 18612 17960 18624
rect 17736 18584 17960 18612
rect 17736 18572 17742 18584
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18417 18615 18475 18621
rect 18417 18581 18429 18615
rect 18463 18612 18475 18615
rect 22002 18612 22008 18624
rect 18463 18584 22008 18612
rect 18463 18581 18475 18584
rect 18417 18575 18475 18581
rect 22002 18572 22008 18584
rect 22060 18572 22066 18624
rect 22097 18615 22155 18621
rect 22097 18581 22109 18615
rect 22143 18612 22155 18615
rect 22370 18612 22376 18624
rect 22143 18584 22376 18612
rect 22143 18581 22155 18584
rect 22097 18575 22155 18581
rect 22370 18572 22376 18584
rect 22428 18572 22434 18624
rect 22557 18615 22615 18621
rect 22557 18581 22569 18615
rect 22603 18612 22615 18615
rect 24412 18612 24440 18652
rect 25222 18640 25228 18652
rect 25280 18640 25286 18692
rect 22603 18584 24440 18612
rect 22603 18581 22615 18584
rect 22557 18575 22615 18581
rect 24486 18572 24492 18624
rect 24544 18612 24550 18624
rect 24581 18615 24639 18621
rect 24581 18612 24593 18615
rect 24544 18584 24593 18612
rect 24544 18572 24550 18584
rect 24581 18581 24593 18584
rect 24627 18581 24639 18615
rect 24581 18575 24639 18581
rect 24854 18572 24860 18624
rect 24912 18612 24918 18624
rect 24949 18615 25007 18621
rect 24949 18612 24961 18615
rect 24912 18584 24961 18612
rect 24912 18572 24918 18584
rect 24949 18581 24961 18584
rect 24995 18581 25007 18615
rect 24949 18575 25007 18581
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 1578 18368 1584 18420
rect 1636 18368 1642 18420
rect 2133 18411 2191 18417
rect 2133 18377 2145 18411
rect 2179 18408 2191 18411
rect 2222 18408 2228 18420
rect 2179 18380 2228 18408
rect 2179 18377 2191 18380
rect 2133 18371 2191 18377
rect 2222 18368 2228 18380
rect 2280 18368 2286 18420
rect 3786 18368 3792 18420
rect 3844 18408 3850 18420
rect 4525 18411 4583 18417
rect 4525 18408 4537 18411
rect 3844 18380 4537 18408
rect 3844 18368 3850 18380
rect 4525 18377 4537 18380
rect 4571 18377 4583 18411
rect 4525 18371 4583 18377
rect 4890 18368 4896 18420
rect 4948 18408 4954 18420
rect 5169 18411 5227 18417
rect 5169 18408 5181 18411
rect 4948 18380 5181 18408
rect 4948 18368 4954 18380
rect 5169 18377 5181 18380
rect 5215 18377 5227 18411
rect 5169 18371 5227 18377
rect 5718 18368 5724 18420
rect 5776 18408 5782 18420
rect 5813 18411 5871 18417
rect 5813 18408 5825 18411
rect 5776 18380 5825 18408
rect 5776 18368 5782 18380
rect 5813 18377 5825 18380
rect 5859 18377 5871 18411
rect 5813 18371 5871 18377
rect 5994 18368 6000 18420
rect 6052 18408 6058 18420
rect 8297 18411 8355 18417
rect 8297 18408 8309 18411
rect 6052 18380 8309 18408
rect 6052 18368 6058 18380
rect 8297 18377 8309 18380
rect 8343 18377 8355 18411
rect 8297 18371 8355 18377
rect 8570 18368 8576 18420
rect 8628 18408 8634 18420
rect 11793 18411 11851 18417
rect 11793 18408 11805 18411
rect 8628 18380 11805 18408
rect 8628 18368 8634 18380
rect 11793 18377 11805 18380
rect 11839 18377 11851 18411
rect 11793 18371 11851 18377
rect 12066 18368 12072 18420
rect 12124 18408 12130 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 12124 18380 12173 18408
rect 12124 18368 12130 18380
rect 12161 18377 12173 18380
rect 12207 18377 12219 18411
rect 12161 18371 12219 18377
rect 14458 18368 14464 18420
rect 14516 18408 14522 18420
rect 15565 18411 15623 18417
rect 15565 18408 15577 18411
rect 14516 18380 15577 18408
rect 14516 18368 14522 18380
rect 15565 18377 15577 18380
rect 15611 18377 15623 18411
rect 15565 18371 15623 18377
rect 15657 18411 15715 18417
rect 15657 18377 15669 18411
rect 15703 18408 15715 18411
rect 15746 18408 15752 18420
rect 15703 18380 15752 18408
rect 15703 18377 15715 18380
rect 15657 18371 15715 18377
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 16482 18368 16488 18420
rect 16540 18408 16546 18420
rect 18509 18411 18567 18417
rect 18509 18408 18521 18411
rect 16540 18380 18521 18408
rect 16540 18368 16546 18380
rect 18509 18377 18521 18380
rect 18555 18377 18567 18411
rect 18509 18371 18567 18377
rect 19150 18368 19156 18420
rect 19208 18408 19214 18420
rect 19208 18380 23244 18408
rect 19208 18368 19214 18380
rect 6086 18340 6092 18352
rect 4724 18312 6092 18340
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 2777 18275 2835 18281
rect 2777 18272 2789 18275
rect 1811 18244 2789 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 2777 18241 2789 18244
rect 2823 18272 2835 18275
rect 2866 18272 2872 18284
rect 2823 18244 2872 18272
rect 2823 18241 2835 18244
rect 2777 18235 2835 18241
rect 2866 18232 2872 18244
rect 2924 18232 2930 18284
rect 2961 18275 3019 18281
rect 2961 18241 2973 18275
rect 3007 18272 3019 18275
rect 3421 18275 3479 18281
rect 3421 18272 3433 18275
rect 3007 18244 3433 18272
rect 3007 18241 3019 18244
rect 2961 18235 3019 18241
rect 3421 18241 3433 18244
rect 3467 18272 3479 18275
rect 4062 18272 4068 18284
rect 3467 18244 4068 18272
rect 3467 18241 3479 18244
rect 3421 18235 3479 18241
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 4724 18281 4752 18312
rect 6086 18300 6092 18312
rect 6144 18300 6150 18352
rect 6733 18343 6791 18349
rect 6733 18309 6745 18343
rect 6779 18340 6791 18343
rect 10502 18340 10508 18352
rect 6779 18312 7696 18340
rect 10442 18312 10508 18340
rect 6779 18309 6791 18312
rect 6733 18303 6791 18309
rect 7668 18284 7696 18312
rect 10502 18300 10508 18312
rect 10560 18340 10566 18352
rect 11057 18343 11115 18349
rect 11057 18340 11069 18343
rect 10560 18312 11069 18340
rect 10560 18300 10566 18312
rect 11057 18309 11069 18312
rect 11103 18309 11115 18343
rect 11057 18303 11115 18309
rect 11330 18300 11336 18352
rect 11388 18300 11394 18352
rect 14366 18340 14372 18352
rect 11440 18312 14372 18340
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18241 4767 18275
rect 4709 18235 4767 18241
rect 5353 18275 5411 18281
rect 5353 18241 5365 18275
rect 5399 18272 5411 18275
rect 5534 18272 5540 18284
rect 5399 18244 5540 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 5534 18232 5540 18244
rect 5592 18232 5598 18284
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 6914 18272 6920 18284
rect 6043 18244 6920 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 7098 18232 7104 18284
rect 7156 18272 7162 18284
rect 7193 18275 7251 18281
rect 7193 18272 7205 18275
rect 7156 18244 7205 18272
rect 7156 18232 7162 18244
rect 7193 18241 7205 18244
rect 7239 18241 7251 18275
rect 7193 18235 7251 18241
rect 7650 18232 7656 18284
rect 7708 18272 7714 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7708 18244 7849 18272
rect 7708 18232 7714 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 8478 18232 8484 18284
rect 8536 18232 8542 18284
rect 8938 18232 8944 18284
rect 8996 18232 9002 18284
rect 10962 18232 10968 18284
rect 11020 18272 11026 18284
rect 11440 18272 11468 18312
rect 14366 18300 14372 18312
rect 14424 18300 14430 18352
rect 14734 18300 14740 18352
rect 14792 18340 14798 18352
rect 15470 18340 15476 18352
rect 14792 18312 15476 18340
rect 14792 18300 14798 18312
rect 15470 18300 15476 18312
rect 15528 18300 15534 18352
rect 16574 18300 16580 18352
rect 16632 18340 16638 18352
rect 16632 18312 20024 18340
rect 16632 18300 16638 18312
rect 11020 18244 11468 18272
rect 11020 18232 11026 18244
rect 11974 18232 11980 18284
rect 12032 18272 12038 18284
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 12032 18244 12265 18272
rect 12032 18232 12038 18244
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 12986 18232 12992 18284
rect 13044 18272 13050 18284
rect 13354 18272 13360 18284
rect 13044 18244 13360 18272
rect 13044 18232 13050 18244
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 15102 18232 15108 18284
rect 15160 18272 15166 18284
rect 15160 18244 15884 18272
rect 15160 18232 15166 18244
rect 3789 18207 3847 18213
rect 3789 18173 3801 18207
rect 3835 18204 3847 18207
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 3835 18176 3893 18204
rect 3835 18173 3847 18176
rect 3789 18167 3847 18173
rect 3881 18173 3893 18176
rect 3927 18204 3939 18207
rect 5626 18204 5632 18216
rect 3927 18176 5632 18204
rect 3927 18173 3939 18176
rect 3881 18167 3939 18173
rect 5626 18164 5632 18176
rect 5684 18164 5690 18216
rect 6549 18207 6607 18213
rect 6549 18173 6561 18207
rect 6595 18204 6607 18207
rect 7558 18204 7564 18216
rect 6595 18176 7564 18204
rect 6595 18173 6607 18176
rect 6549 18167 6607 18173
rect 7558 18164 7564 18176
rect 7616 18164 7622 18216
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18204 9275 18207
rect 10778 18204 10784 18216
rect 9263 18176 10784 18204
rect 9263 18173 9275 18176
rect 9217 18167 9275 18173
rect 10778 18164 10784 18176
rect 10836 18164 10842 18216
rect 10888 18176 11376 18204
rect 7009 18139 7067 18145
rect 7009 18105 7021 18139
rect 7055 18136 7067 18139
rect 8846 18136 8852 18148
rect 7055 18108 8852 18136
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 8846 18096 8852 18108
rect 8904 18096 8910 18148
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18068 3295 18071
rect 4062 18068 4068 18080
rect 3283 18040 4068 18068
rect 3283 18037 3295 18040
rect 3237 18031 3295 18037
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 7650 18028 7656 18080
rect 7708 18028 7714 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 9824 18040 10701 18068
rect 9824 18028 9830 18040
rect 10689 18037 10701 18040
rect 10735 18068 10747 18071
rect 10888 18068 10916 18176
rect 10735 18040 10916 18068
rect 11348 18068 11376 18176
rect 12158 18164 12164 18216
rect 12216 18204 12222 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 12216 18176 12449 18204
rect 12216 18164 12222 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 15749 18207 15807 18213
rect 15749 18173 15761 18207
rect 15795 18173 15807 18207
rect 15749 18167 15807 18173
rect 11698 18096 11704 18148
rect 11756 18136 11762 18148
rect 15197 18139 15255 18145
rect 15197 18136 15209 18139
rect 11756 18108 15209 18136
rect 11756 18096 11762 18108
rect 15197 18105 15209 18108
rect 15243 18105 15255 18139
rect 15197 18099 15255 18105
rect 15764 18068 15792 18167
rect 15856 18136 15884 18244
rect 16758 18232 16764 18284
rect 16816 18272 16822 18284
rect 17221 18275 17279 18281
rect 17221 18272 17233 18275
rect 16816 18244 17233 18272
rect 16816 18232 16822 18244
rect 17221 18241 17233 18244
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18272 17371 18275
rect 18417 18275 18475 18281
rect 17359 18244 17632 18272
rect 17359 18241 17371 18244
rect 17313 18235 17371 18241
rect 15930 18164 15936 18216
rect 15988 18204 15994 18216
rect 16206 18204 16212 18216
rect 15988 18176 16212 18204
rect 15988 18164 15994 18176
rect 16206 18164 16212 18176
rect 16264 18204 16270 18216
rect 17497 18207 17555 18213
rect 16264 18176 17264 18204
rect 16264 18164 16270 18176
rect 17236 18148 17264 18176
rect 17497 18173 17509 18207
rect 17543 18173 17555 18207
rect 17604 18204 17632 18244
rect 18417 18241 18429 18275
rect 18463 18272 18475 18275
rect 18506 18272 18512 18284
rect 18463 18244 18512 18272
rect 18463 18241 18475 18244
rect 18417 18235 18475 18241
rect 18506 18232 18512 18244
rect 18564 18272 18570 18284
rect 19518 18272 19524 18284
rect 18564 18244 19524 18272
rect 18564 18232 18570 18244
rect 19518 18232 19524 18244
rect 19576 18232 19582 18284
rect 19613 18275 19671 18281
rect 19613 18241 19625 18275
rect 19659 18272 19671 18275
rect 19996 18272 20024 18312
rect 20254 18300 20260 18352
rect 20312 18340 20318 18352
rect 20809 18343 20867 18349
rect 20809 18340 20821 18343
rect 20312 18312 20821 18340
rect 20312 18300 20318 18312
rect 20809 18309 20821 18312
rect 20855 18309 20867 18343
rect 20809 18303 20867 18309
rect 20898 18300 20904 18352
rect 20956 18300 20962 18352
rect 23106 18340 23112 18352
rect 21008 18312 23112 18340
rect 21008 18272 21036 18312
rect 23106 18300 23112 18312
rect 23164 18300 23170 18352
rect 19659 18244 19932 18272
rect 19996 18244 21036 18272
rect 19659 18241 19671 18244
rect 19613 18235 19671 18241
rect 17678 18204 17684 18216
rect 17604 18176 17684 18204
rect 17497 18167 17555 18173
rect 16853 18139 16911 18145
rect 16853 18136 16865 18139
rect 15856 18108 16865 18136
rect 16853 18105 16865 18108
rect 16899 18105 16911 18139
rect 16853 18099 16911 18105
rect 17218 18096 17224 18148
rect 17276 18096 17282 18148
rect 11348 18040 15792 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 16206 18028 16212 18080
rect 16264 18028 16270 18080
rect 16482 18028 16488 18080
rect 16540 18068 16546 18080
rect 17512 18068 17540 18167
rect 17678 18164 17684 18176
rect 17736 18204 17742 18216
rect 17736 18176 18184 18204
rect 17736 18164 17742 18176
rect 18156 18136 18184 18176
rect 18690 18164 18696 18216
rect 18748 18164 18754 18216
rect 19702 18164 19708 18216
rect 19760 18164 19766 18216
rect 19797 18207 19855 18213
rect 19797 18173 19809 18207
rect 19843 18173 19855 18207
rect 19797 18167 19855 18173
rect 19150 18136 19156 18148
rect 18156 18108 19156 18136
rect 19150 18096 19156 18108
rect 19208 18096 19214 18148
rect 19334 18096 19340 18148
rect 19392 18136 19398 18148
rect 19812 18136 19840 18167
rect 19392 18108 19840 18136
rect 19904 18136 19932 18244
rect 21358 18232 21364 18284
rect 21416 18272 21422 18284
rect 21910 18272 21916 18284
rect 21416 18244 21916 18272
rect 21416 18232 21422 18244
rect 21910 18232 21916 18244
rect 21968 18232 21974 18284
rect 22002 18232 22008 18284
rect 22060 18232 22066 18284
rect 23216 18272 23244 18380
rect 23290 18368 23296 18420
rect 23348 18368 23354 18420
rect 24946 18368 24952 18420
rect 25004 18408 25010 18420
rect 25041 18411 25099 18417
rect 25041 18408 25053 18411
rect 25004 18380 25053 18408
rect 25004 18368 25010 18380
rect 25041 18377 25053 18380
rect 25087 18377 25099 18411
rect 25041 18371 25099 18377
rect 23750 18272 23756 18284
rect 23216 18244 23756 18272
rect 23750 18232 23756 18244
rect 23808 18232 23814 18284
rect 24949 18275 25007 18281
rect 24949 18241 24961 18275
rect 24995 18241 25007 18275
rect 24949 18235 25007 18241
rect 20993 18207 21051 18213
rect 20993 18173 21005 18207
rect 21039 18173 21051 18207
rect 20993 18167 21051 18173
rect 20714 18136 20720 18148
rect 19904 18108 20720 18136
rect 19392 18096 19398 18108
rect 20714 18096 20720 18108
rect 20772 18096 20778 18148
rect 20806 18096 20812 18148
rect 20864 18136 20870 18148
rect 21008 18136 21036 18167
rect 21082 18164 21088 18216
rect 21140 18204 21146 18216
rect 21453 18207 21511 18213
rect 21453 18204 21465 18207
rect 21140 18176 21465 18204
rect 21140 18164 21146 18176
rect 21453 18173 21465 18176
rect 21499 18173 21511 18207
rect 21453 18167 21511 18173
rect 24394 18164 24400 18216
rect 24452 18204 24458 18216
rect 24964 18204 24992 18235
rect 24452 18176 24992 18204
rect 25225 18207 25283 18213
rect 24452 18164 24458 18176
rect 25225 18173 25237 18207
rect 25271 18204 25283 18207
rect 25498 18204 25504 18216
rect 25271 18176 25504 18204
rect 25271 18173 25283 18176
rect 25225 18167 25283 18173
rect 25498 18164 25504 18176
rect 25556 18164 25562 18216
rect 20864 18108 21036 18136
rect 20864 18096 20870 18108
rect 16540 18040 17540 18068
rect 16540 18028 16546 18040
rect 17586 18028 17592 18080
rect 17644 18068 17650 18080
rect 18049 18071 18107 18077
rect 18049 18068 18061 18071
rect 17644 18040 18061 18068
rect 17644 18028 17650 18040
rect 18049 18037 18061 18040
rect 18095 18037 18107 18071
rect 18049 18031 18107 18037
rect 19245 18071 19303 18077
rect 19245 18037 19257 18071
rect 19291 18068 19303 18071
rect 19886 18068 19892 18080
rect 19291 18040 19892 18068
rect 19291 18037 19303 18040
rect 19245 18031 19303 18037
rect 19886 18028 19892 18040
rect 19944 18028 19950 18080
rect 20441 18071 20499 18077
rect 20441 18037 20453 18071
rect 20487 18068 20499 18071
rect 20990 18068 20996 18080
rect 20487 18040 20996 18068
rect 20487 18037 20499 18040
rect 20441 18031 20499 18037
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 23474 18028 23480 18080
rect 23532 18068 23538 18080
rect 24581 18071 24639 18077
rect 24581 18068 24593 18071
rect 23532 18040 24593 18068
rect 23532 18028 23538 18040
rect 24581 18037 24593 18040
rect 24627 18037 24639 18071
rect 24581 18031 24639 18037
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 3237 17867 3295 17873
rect 3237 17833 3249 17867
rect 3283 17864 3295 17867
rect 4522 17864 4528 17876
rect 3283 17836 4528 17864
rect 3283 17833 3295 17836
rect 3237 17827 3295 17833
rect 4522 17824 4528 17836
rect 4580 17824 4586 17876
rect 6362 17824 6368 17876
rect 6420 17864 6426 17876
rect 6457 17867 6515 17873
rect 6457 17864 6469 17867
rect 6420 17836 6469 17864
rect 6420 17824 6426 17836
rect 6457 17833 6469 17836
rect 6503 17833 6515 17867
rect 6457 17827 6515 17833
rect 7006 17824 7012 17876
rect 7064 17864 7070 17876
rect 7745 17867 7803 17873
rect 7745 17864 7757 17867
rect 7064 17836 7757 17864
rect 7064 17824 7070 17836
rect 7745 17833 7757 17836
rect 7791 17833 7803 17867
rect 7745 17827 7803 17833
rect 9122 17824 9128 17876
rect 9180 17864 9186 17876
rect 11146 17864 11152 17876
rect 9180 17836 11152 17864
rect 9180 17824 9186 17836
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 11517 17867 11575 17873
rect 11517 17833 11529 17867
rect 11563 17864 11575 17867
rect 12066 17864 12072 17876
rect 11563 17836 12072 17864
rect 11563 17833 11575 17836
rect 11517 17827 11575 17833
rect 12066 17824 12072 17836
rect 12124 17864 12130 17876
rect 12250 17864 12256 17876
rect 12124 17836 12256 17864
rect 12124 17824 12130 17836
rect 12250 17824 12256 17836
rect 12308 17824 12314 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13262 17864 13268 17876
rect 12492 17836 13268 17864
rect 12492 17824 12498 17836
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 13725 17867 13783 17873
rect 13725 17833 13737 17867
rect 13771 17864 13783 17867
rect 13814 17864 13820 17876
rect 13771 17836 13820 17864
rect 13771 17833 13783 17836
rect 13725 17827 13783 17833
rect 13814 17824 13820 17836
rect 13872 17864 13878 17876
rect 16482 17864 16488 17876
rect 13872 17836 16488 17864
rect 13872 17824 13878 17836
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 17126 17824 17132 17876
rect 17184 17824 17190 17876
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 20622 17864 20628 17876
rect 17276 17836 20628 17864
rect 17276 17824 17282 17836
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 20980 17867 21038 17873
rect 20980 17833 20992 17867
rect 21026 17864 21038 17867
rect 22370 17864 22376 17876
rect 21026 17836 22376 17864
rect 21026 17833 21038 17836
rect 20980 17827 21038 17833
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 22465 17867 22523 17873
rect 22465 17833 22477 17867
rect 22511 17864 22523 17867
rect 22646 17864 22652 17876
rect 22511 17836 22652 17864
rect 22511 17833 22523 17836
rect 22465 17827 22523 17833
rect 22646 17824 22652 17836
rect 22704 17824 22710 17876
rect 6638 17796 6644 17808
rect 5184 17768 6644 17796
rect 5184 17737 5212 17768
rect 6638 17756 6644 17768
rect 6696 17756 6702 17808
rect 16669 17799 16727 17805
rect 16669 17765 16681 17799
rect 16715 17796 16727 17799
rect 17310 17796 17316 17808
rect 16715 17768 17316 17796
rect 16715 17765 16727 17768
rect 16669 17759 16727 17765
rect 17310 17756 17316 17768
rect 17368 17756 17374 17808
rect 19306 17768 20392 17796
rect 5169 17731 5227 17737
rect 5169 17697 5181 17731
rect 5215 17697 5227 17731
rect 5169 17691 5227 17697
rect 5445 17731 5503 17737
rect 5445 17697 5457 17731
rect 5491 17728 5503 17731
rect 6178 17728 6184 17740
rect 5491 17700 6184 17728
rect 5491 17697 5503 17700
rect 5445 17691 5503 17697
rect 6178 17688 6184 17700
rect 6236 17688 6242 17740
rect 6546 17688 6552 17740
rect 6604 17728 6610 17740
rect 6604 17700 7972 17728
rect 6604 17688 6610 17700
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 4706 17660 4712 17672
rect 4295 17632 4712 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 5810 17620 5816 17672
rect 5868 17660 5874 17672
rect 6641 17663 6699 17669
rect 6641 17660 6653 17663
rect 5868 17632 6653 17660
rect 5868 17620 5874 17632
rect 6641 17629 6653 17632
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17660 7343 17663
rect 7558 17660 7564 17672
rect 7331 17632 7564 17660
rect 7331 17629 7343 17632
rect 7285 17623 7343 17629
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 7944 17669 7972 17700
rect 8938 17688 8944 17740
rect 8996 17728 9002 17740
rect 9769 17731 9827 17737
rect 9769 17728 9781 17731
rect 8996 17700 9781 17728
rect 8996 17688 9002 17700
rect 9769 17697 9781 17700
rect 9815 17728 9827 17731
rect 11698 17728 11704 17740
rect 9815 17700 11704 17728
rect 9815 17697 9827 17700
rect 9769 17691 9827 17697
rect 11698 17688 11704 17700
rect 11756 17728 11762 17740
rect 11882 17728 11888 17740
rect 11756 17700 11888 17728
rect 11756 17688 11762 17700
rect 11882 17688 11888 17700
rect 11940 17728 11946 17740
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11940 17700 11989 17728
rect 11940 17688 11946 17700
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 12253 17731 12311 17737
rect 12253 17697 12265 17731
rect 12299 17728 12311 17731
rect 12342 17728 12348 17740
rect 12299 17700 12348 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 12342 17688 12348 17700
rect 12400 17728 12406 17740
rect 13446 17728 13452 17740
rect 12400 17700 13452 17728
rect 12400 17688 12406 17700
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 13722 17688 13728 17740
rect 13780 17728 13786 17740
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 13780 17700 14289 17728
rect 13780 17688 13786 17700
rect 14277 17697 14289 17700
rect 14323 17697 14335 17731
rect 14277 17691 14335 17697
rect 14734 17688 14740 17740
rect 14792 17728 14798 17740
rect 14918 17728 14924 17740
rect 14792 17700 14924 17728
rect 14792 17688 14798 17700
rect 14918 17688 14924 17700
rect 14976 17688 14982 17740
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 15838 17728 15844 17740
rect 15252 17700 15844 17728
rect 15252 17688 15258 17700
rect 15838 17688 15844 17700
rect 15896 17688 15902 17740
rect 15930 17688 15936 17740
rect 15988 17728 15994 17740
rect 15988 17700 16436 17728
rect 15988 17688 15994 17700
rect 7929 17663 7987 17669
rect 7929 17629 7941 17663
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17660 8631 17663
rect 9122 17660 9128 17672
rect 8619 17632 9128 17660
rect 8619 17629 8631 17632
rect 8573 17623 8631 17629
rect 9122 17620 9128 17632
rect 9180 17620 9186 17672
rect 9309 17663 9367 17669
rect 9309 17629 9321 17663
rect 9355 17629 9367 17663
rect 16408 17660 16436 17700
rect 16574 17688 16580 17740
rect 16632 17728 16638 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 16632 17700 17693 17728
rect 16632 17688 16638 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 17589 17663 17647 17669
rect 17589 17660 17601 17663
rect 16408 17632 17601 17660
rect 9309 17623 9367 17629
rect 17589 17629 17601 17632
rect 17635 17629 17647 17663
rect 17589 17623 17647 17629
rect 4338 17552 4344 17604
rect 4396 17592 4402 17604
rect 4396 17564 9168 17592
rect 4396 17552 4402 17564
rect 4522 17484 4528 17536
rect 4580 17484 4586 17536
rect 7098 17484 7104 17536
rect 7156 17484 7162 17536
rect 8386 17484 8392 17536
rect 8444 17484 8450 17536
rect 9140 17533 9168 17564
rect 9125 17527 9183 17533
rect 9125 17493 9137 17527
rect 9171 17493 9183 17527
rect 9324 17524 9352 17623
rect 17862 17620 17868 17672
rect 17920 17660 17926 17672
rect 18785 17663 18843 17669
rect 18785 17660 18797 17663
rect 17920 17632 18797 17660
rect 17920 17620 17926 17632
rect 18785 17629 18797 17632
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 9490 17552 9496 17604
rect 9548 17592 9554 17604
rect 10042 17592 10048 17604
rect 9548 17564 10048 17592
rect 9548 17552 9554 17564
rect 10042 17552 10048 17564
rect 10100 17552 10106 17604
rect 10134 17552 10140 17604
rect 10192 17592 10198 17604
rect 10502 17592 10508 17604
rect 10192 17564 10508 17592
rect 10192 17552 10198 17564
rect 10502 17552 10508 17564
rect 10560 17552 10566 17604
rect 12986 17552 12992 17604
rect 13044 17552 13050 17604
rect 14734 17552 14740 17604
rect 14792 17592 14798 17604
rect 15654 17592 15660 17604
rect 14792 17564 15660 17592
rect 14792 17552 14798 17564
rect 15654 17552 15660 17564
rect 15712 17552 15718 17604
rect 19306 17592 19334 17768
rect 19794 17688 19800 17740
rect 19852 17728 19858 17740
rect 19889 17731 19947 17737
rect 19889 17728 19901 17731
rect 19852 17700 19901 17728
rect 19852 17688 19858 17700
rect 19889 17697 19901 17700
rect 19935 17697 19947 17731
rect 19889 17691 19947 17697
rect 20073 17731 20131 17737
rect 20073 17697 20085 17731
rect 20119 17728 20131 17731
rect 20254 17728 20260 17740
rect 20119 17700 20260 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 20254 17688 20260 17700
rect 20312 17688 20318 17740
rect 16500 17564 19334 17592
rect 11422 17524 11428 17536
rect 9324 17496 11428 17524
rect 9125 17487 9183 17493
rect 11422 17484 11428 17496
rect 11480 17484 11486 17536
rect 12250 17484 12256 17536
rect 12308 17524 12314 17536
rect 14274 17524 14280 17536
rect 12308 17496 14280 17524
rect 12308 17484 12314 17496
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 14458 17484 14464 17536
rect 14516 17524 14522 17536
rect 16500 17524 16528 17564
rect 14516 17496 16528 17524
rect 14516 17484 14522 17496
rect 17494 17484 17500 17536
rect 17552 17484 17558 17536
rect 17678 17484 17684 17536
rect 17736 17524 17742 17536
rect 18141 17527 18199 17533
rect 18141 17524 18153 17527
rect 17736 17496 18153 17524
rect 17736 17484 17742 17496
rect 18141 17493 18153 17496
rect 18187 17493 18199 17527
rect 18141 17487 18199 17493
rect 18598 17484 18604 17536
rect 18656 17484 18662 17536
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17524 19487 17527
rect 19702 17524 19708 17536
rect 19475 17496 19708 17524
rect 19475 17493 19487 17496
rect 19429 17487 19487 17493
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 19797 17527 19855 17533
rect 19797 17493 19809 17527
rect 19843 17524 19855 17527
rect 20162 17524 20168 17536
rect 19843 17496 20168 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 20162 17484 20168 17496
rect 20220 17484 20226 17536
rect 20364 17524 20392 17768
rect 22186 17756 22192 17808
rect 22244 17796 22250 17808
rect 23474 17796 23480 17808
rect 22244 17768 23480 17796
rect 22244 17756 22250 17768
rect 23474 17756 23480 17768
rect 23532 17756 23538 17808
rect 20717 17731 20775 17737
rect 20717 17697 20729 17731
rect 20763 17728 20775 17731
rect 22554 17728 22560 17740
rect 20763 17700 22560 17728
rect 20763 17697 20775 17700
rect 20717 17691 20775 17697
rect 22554 17688 22560 17700
rect 22612 17728 22618 17740
rect 23290 17728 23296 17740
rect 22612 17700 23296 17728
rect 22612 17688 22618 17700
rect 23290 17688 23296 17700
rect 23348 17688 23354 17740
rect 23842 17688 23848 17740
rect 23900 17728 23906 17740
rect 24302 17728 24308 17740
rect 23900 17700 24308 17728
rect 23900 17688 23906 17700
rect 24302 17688 24308 17700
rect 24360 17688 24366 17740
rect 23198 17620 23204 17672
rect 23256 17660 23262 17672
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 23256 17632 23673 17660
rect 23256 17620 23262 17632
rect 23661 17629 23673 17632
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 23753 17663 23811 17669
rect 23753 17629 23765 17663
rect 23799 17660 23811 17663
rect 24578 17660 24584 17672
rect 23799 17632 24584 17660
rect 23799 17629 23811 17632
rect 23753 17623 23811 17629
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 21082 17552 21088 17604
rect 21140 17592 21146 17604
rect 21450 17592 21456 17604
rect 21140 17564 21456 17592
rect 21140 17552 21146 17564
rect 21450 17552 21456 17564
rect 21508 17552 21514 17604
rect 22738 17552 22744 17604
rect 22796 17592 22802 17604
rect 22833 17595 22891 17601
rect 22833 17592 22845 17595
rect 22796 17564 22845 17592
rect 22796 17552 22802 17564
rect 22833 17561 22845 17564
rect 22879 17592 22891 17595
rect 23474 17592 23480 17604
rect 22879 17564 23480 17592
rect 22879 17561 22891 17564
rect 22833 17555 22891 17561
rect 23474 17552 23480 17564
rect 23532 17552 23538 17604
rect 24486 17552 24492 17604
rect 24544 17592 24550 17604
rect 24765 17595 24823 17601
rect 24765 17592 24777 17595
rect 24544 17564 24777 17592
rect 24544 17552 24550 17564
rect 24765 17561 24777 17564
rect 24811 17561 24823 17595
rect 24765 17555 24823 17561
rect 24949 17595 25007 17601
rect 24949 17561 24961 17595
rect 24995 17592 25007 17595
rect 25866 17592 25872 17604
rect 24995 17564 25872 17592
rect 24995 17561 25007 17564
rect 24949 17555 25007 17561
rect 25866 17552 25872 17564
rect 25924 17552 25930 17604
rect 22278 17524 22284 17536
rect 20364 17496 22284 17524
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 22922 17484 22928 17536
rect 22980 17484 22986 17536
rect 23293 17527 23351 17533
rect 23293 17493 23305 17527
rect 23339 17524 23351 17527
rect 23566 17524 23572 17536
rect 23339 17496 23572 17524
rect 23339 17493 23351 17496
rect 23293 17487 23351 17493
rect 23566 17484 23572 17496
rect 23624 17484 23630 17536
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 3881 17323 3939 17329
rect 3881 17289 3893 17323
rect 3927 17320 3939 17323
rect 3970 17320 3976 17332
rect 3927 17292 3976 17320
rect 3927 17289 3939 17292
rect 3881 17283 3939 17289
rect 3970 17280 3976 17292
rect 4028 17280 4034 17332
rect 6546 17280 6552 17332
rect 6604 17280 6610 17332
rect 7190 17280 7196 17332
rect 7248 17280 7254 17332
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 7837 17323 7895 17329
rect 7837 17320 7849 17323
rect 7432 17292 7849 17320
rect 7432 17280 7438 17292
rect 7837 17289 7849 17292
rect 7883 17289 7895 17323
rect 7837 17283 7895 17289
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 11882 17320 11888 17332
rect 8444 17292 11888 17320
rect 8444 17280 8450 17292
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 12618 17280 12624 17332
rect 12676 17320 12682 17332
rect 15841 17323 15899 17329
rect 15841 17320 15853 17323
rect 12676 17292 15853 17320
rect 12676 17280 12682 17292
rect 15841 17289 15853 17292
rect 15887 17289 15899 17323
rect 15841 17283 15899 17289
rect 15948 17292 19932 17320
rect 8294 17252 8300 17264
rect 6748 17224 8300 17252
rect 3789 17187 3847 17193
rect 3789 17153 3801 17187
rect 3835 17184 3847 17187
rect 4065 17187 4123 17193
rect 4065 17184 4077 17187
rect 3835 17156 4077 17184
rect 3835 17153 3847 17156
rect 3789 17147 3847 17153
rect 4065 17153 4077 17156
rect 4111 17184 4123 17187
rect 5534 17184 5540 17196
rect 4111 17156 5540 17184
rect 4111 17153 4123 17156
rect 4065 17147 4123 17153
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 6748 17193 6776 17224
rect 8294 17212 8300 17224
rect 8352 17212 8358 17264
rect 9493 17255 9551 17261
rect 9493 17221 9505 17255
rect 9539 17252 9551 17255
rect 9766 17252 9772 17264
rect 9539 17224 9772 17252
rect 9539 17221 9551 17224
rect 9493 17215 9551 17221
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 10134 17212 10140 17264
rect 10192 17212 10198 17264
rect 11977 17255 12035 17261
rect 11977 17221 11989 17255
rect 12023 17252 12035 17255
rect 12066 17252 12072 17264
rect 12023 17224 12072 17252
rect 12023 17221 12035 17224
rect 11977 17215 12035 17221
rect 12066 17212 12072 17224
rect 12124 17212 12130 17264
rect 13262 17212 13268 17264
rect 13320 17252 13326 17264
rect 15948 17252 15976 17292
rect 13320 17224 15976 17252
rect 13320 17212 13326 17224
rect 16390 17212 16396 17264
rect 16448 17252 16454 17264
rect 16448 17224 17448 17252
rect 16448 17212 16454 17224
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 6822 17184 6828 17196
rect 6779 17156 6828 17184
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 6822 17144 6828 17156
rect 6880 17144 6886 17196
rect 7377 17187 7435 17193
rect 7377 17153 7389 17187
rect 7423 17184 7435 17187
rect 7466 17184 7472 17196
rect 7423 17156 7472 17184
rect 7423 17153 7435 17156
rect 7377 17147 7435 17153
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17085 4583 17119
rect 4525 17079 4583 17085
rect 4801 17119 4859 17125
rect 4801 17085 4813 17119
rect 4847 17116 4859 17119
rect 7834 17116 7840 17128
rect 4847 17088 7840 17116
rect 4847 17085 4859 17088
rect 4801 17079 4859 17085
rect 4540 16980 4568 17079
rect 7834 17076 7840 17088
rect 7892 17076 7898 17128
rect 5074 17008 5080 17060
rect 5132 17048 5138 17060
rect 8036 17048 8064 17147
rect 8110 17076 8116 17128
rect 8168 17116 8174 17128
rect 8772 17116 8800 17147
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9217 17187 9275 17193
rect 9217 17184 9229 17187
rect 8996 17156 9229 17184
rect 8996 17144 9002 17156
rect 9217 17153 9229 17156
rect 9263 17153 9275 17187
rect 9217 17147 9275 17153
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 14090 17184 14096 17196
rect 13110 17170 14096 17184
rect 13096 17156 14096 17170
rect 9950 17116 9956 17128
rect 8168 17088 9956 17116
rect 8168 17076 8174 17088
rect 9950 17076 9956 17088
rect 10008 17076 10014 17128
rect 10042 17076 10048 17128
rect 10100 17116 10106 17128
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10100 17088 10977 17116
rect 10100 17076 10106 17088
rect 10965 17085 10977 17088
rect 11011 17085 11023 17119
rect 12526 17116 12532 17128
rect 10965 17079 11023 17085
rect 11256 17088 12532 17116
rect 5132 17020 8064 17048
rect 8573 17051 8631 17057
rect 5132 17008 5138 17020
rect 8573 17017 8585 17051
rect 8619 17048 8631 17051
rect 8754 17048 8760 17060
rect 8619 17020 8760 17048
rect 8619 17017 8631 17020
rect 8573 17011 8631 17017
rect 8754 17008 8760 17020
rect 8812 17008 8818 17060
rect 10042 16980 10048 16992
rect 4540 16952 10048 16980
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10594 16980 10600 16992
rect 10192 16952 10600 16980
rect 10192 16940 10198 16952
rect 10594 16940 10600 16952
rect 10652 16980 10658 16992
rect 11256 16989 11284 17088
rect 12526 17076 12532 17088
rect 12584 17116 12590 17128
rect 12986 17116 12992 17128
rect 12584 17088 12992 17116
rect 12584 17076 12590 17088
rect 12986 17076 12992 17088
rect 13044 17116 13050 17128
rect 13096 17116 13124 17156
rect 14090 17144 14096 17156
rect 14148 17184 14154 17196
rect 14461 17187 14519 17193
rect 14461 17184 14473 17187
rect 14148 17156 14473 17184
rect 14148 17144 14154 17156
rect 14461 17153 14473 17156
rect 14507 17184 14519 17187
rect 14734 17184 14740 17196
rect 14507 17156 14740 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 14734 17144 14740 17156
rect 14792 17144 14798 17196
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 13044 17088 13124 17116
rect 13044 17076 13050 17088
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13872 17088 13921 17116
rect 13872 17076 13878 17088
rect 13909 17085 13921 17088
rect 13955 17085 13967 17119
rect 13909 17079 13967 17085
rect 13446 17008 13452 17060
rect 13504 17008 13510 17060
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 14829 17051 14887 17057
rect 14829 17048 14841 17051
rect 13596 17020 14841 17048
rect 13596 17008 13602 17020
rect 14829 17017 14841 17020
rect 14875 17017 14887 17051
rect 15028 17048 15056 17147
rect 15194 17144 15200 17196
rect 15252 17184 15258 17196
rect 15252 17156 16068 17184
rect 15252 17144 15258 17156
rect 15286 17076 15292 17128
rect 15344 17116 15350 17128
rect 15930 17116 15936 17128
rect 15344 17088 15936 17116
rect 15344 17076 15350 17088
rect 15930 17076 15936 17088
rect 15988 17076 15994 17128
rect 16040 17125 16068 17156
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17221 17187 17279 17193
rect 17221 17184 17233 17187
rect 17000 17156 17233 17184
rect 17000 17144 17006 17156
rect 17221 17153 17233 17156
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17420 17125 17448 17224
rect 17678 17212 17684 17264
rect 17736 17252 17742 17264
rect 19904 17252 19932 17292
rect 20070 17280 20076 17332
rect 20128 17320 20134 17332
rect 20533 17323 20591 17329
rect 20533 17320 20545 17323
rect 20128 17292 20545 17320
rect 20128 17280 20134 17292
rect 20533 17289 20545 17292
rect 20579 17289 20591 17323
rect 20533 17283 20591 17289
rect 21082 17280 21088 17332
rect 21140 17320 21146 17332
rect 21818 17320 21824 17332
rect 21140 17292 21824 17320
rect 21140 17280 21146 17292
rect 21818 17280 21824 17292
rect 21876 17280 21882 17332
rect 22738 17320 22744 17332
rect 22296 17292 22744 17320
rect 22094 17252 22100 17264
rect 17736 17224 19090 17252
rect 19904 17224 22100 17252
rect 17736 17212 17742 17224
rect 22094 17212 22100 17224
rect 22152 17212 22158 17264
rect 18322 17144 18328 17196
rect 18380 17144 18386 17196
rect 21082 17184 21088 17196
rect 19812 17156 21088 17184
rect 16025 17119 16083 17125
rect 16025 17085 16037 17119
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 17313 17119 17371 17125
rect 17313 17085 17325 17119
rect 17359 17085 17371 17119
rect 17313 17079 17371 17085
rect 17405 17119 17463 17125
rect 17405 17085 17417 17119
rect 17451 17085 17463 17119
rect 17405 17079 17463 17085
rect 18601 17119 18659 17125
rect 18601 17085 18613 17119
rect 18647 17116 18659 17119
rect 19242 17116 19248 17128
rect 18647 17088 19248 17116
rect 18647 17085 18659 17088
rect 18601 17079 18659 17085
rect 17218 17048 17224 17060
rect 15028 17020 17224 17048
rect 14829 17011 14887 17017
rect 17218 17008 17224 17020
rect 17276 17008 17282 17060
rect 17328 17048 17356 17079
rect 19242 17076 19248 17088
rect 19300 17076 19306 17128
rect 17957 17051 18015 17057
rect 17957 17048 17969 17051
rect 17328 17020 17969 17048
rect 17957 17017 17969 17020
rect 18003 17048 18015 17051
rect 18322 17048 18328 17060
rect 18003 17020 18328 17048
rect 18003 17017 18015 17020
rect 17957 17011 18015 17017
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 19702 17008 19708 17060
rect 19760 17048 19766 17060
rect 19812 17048 19840 17156
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 21361 17187 21419 17193
rect 21361 17153 21373 17187
rect 21407 17184 21419 17187
rect 22296 17184 22324 17292
rect 22738 17280 22744 17292
rect 22796 17280 22802 17332
rect 24302 17280 24308 17332
rect 24360 17280 24366 17332
rect 22922 17212 22928 17264
rect 22980 17252 22986 17264
rect 22980 17224 23322 17252
rect 22980 17212 22986 17224
rect 21407 17156 22324 17184
rect 21407 17153 21419 17156
rect 21361 17147 21419 17153
rect 22554 17144 22560 17196
rect 22612 17144 22618 17196
rect 24854 17144 24860 17196
rect 24912 17144 24918 17196
rect 25038 17144 25044 17196
rect 25096 17144 25102 17196
rect 20070 17076 20076 17128
rect 20128 17116 20134 17128
rect 21266 17116 21272 17128
rect 20128 17088 21272 17116
rect 20128 17076 20134 17088
rect 21266 17076 21272 17088
rect 21324 17076 21330 17128
rect 21450 17076 21456 17128
rect 21508 17116 21514 17128
rect 21821 17119 21879 17125
rect 21821 17116 21833 17119
rect 21508 17088 21833 17116
rect 21508 17076 21514 17088
rect 21821 17085 21833 17088
rect 21867 17116 21879 17119
rect 22005 17119 22063 17125
rect 22005 17116 22017 17119
rect 21867 17088 22017 17116
rect 21867 17085 21879 17088
rect 21821 17079 21879 17085
rect 22005 17085 22017 17088
rect 22051 17116 22063 17119
rect 22281 17119 22339 17125
rect 22281 17116 22293 17119
rect 22051 17088 22293 17116
rect 22051 17085 22063 17088
rect 22005 17079 22063 17085
rect 22281 17085 22293 17088
rect 22327 17085 22339 17119
rect 22281 17079 22339 17085
rect 22833 17119 22891 17125
rect 22833 17085 22845 17119
rect 22879 17116 22891 17119
rect 25056 17116 25084 17144
rect 22879 17088 25084 17116
rect 22879 17085 22891 17088
rect 22833 17079 22891 17085
rect 22186 17048 22192 17060
rect 19760 17020 19840 17048
rect 20548 17020 22192 17048
rect 19760 17008 19766 17020
rect 11241 16983 11299 16989
rect 11241 16980 11253 16983
rect 10652 16952 11253 16980
rect 10652 16940 10658 16952
rect 11241 16949 11253 16952
rect 11287 16949 11299 16983
rect 11241 16943 11299 16949
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 14458 16980 14464 16992
rect 12032 16952 14464 16980
rect 12032 16940 12038 16952
rect 14458 16940 14464 16952
rect 14516 16940 14522 16992
rect 14734 16940 14740 16992
rect 14792 16980 14798 16992
rect 15473 16983 15531 16989
rect 15473 16980 15485 16983
rect 14792 16952 15485 16980
rect 14792 16940 14798 16952
rect 15473 16949 15485 16952
rect 15519 16949 15531 16983
rect 15473 16943 15531 16949
rect 16850 16940 16856 16992
rect 16908 16940 16914 16992
rect 18138 16940 18144 16992
rect 18196 16980 18202 16992
rect 20548 16980 20576 17020
rect 22186 17008 22192 17020
rect 22244 17008 22250 17060
rect 18196 16952 20576 16980
rect 18196 16940 18202 16952
rect 20622 16940 20628 16992
rect 20680 16980 20686 16992
rect 21177 16983 21235 16989
rect 21177 16980 21189 16983
rect 20680 16952 21189 16980
rect 20680 16940 20686 16952
rect 21177 16949 21189 16952
rect 21223 16949 21235 16983
rect 22296 16980 22324 17079
rect 22370 17008 22376 17060
rect 22428 17048 22434 17060
rect 22554 17048 22560 17060
rect 22428 17020 22560 17048
rect 22428 17008 22434 17020
rect 22554 17008 22560 17020
rect 22612 17008 22618 17060
rect 25041 17051 25099 17057
rect 25041 17017 25053 17051
rect 25087 17048 25099 17051
rect 25682 17048 25688 17060
rect 25087 17020 25688 17048
rect 25087 17017 25099 17020
rect 25041 17011 25099 17017
rect 25682 17008 25688 17020
rect 25740 17008 25746 17060
rect 22922 16980 22928 16992
rect 22296 16952 22928 16980
rect 21177 16943 21235 16949
rect 22922 16940 22928 16952
rect 22980 16980 22986 16992
rect 23842 16980 23848 16992
rect 22980 16952 23848 16980
rect 22980 16940 22986 16952
rect 23842 16940 23848 16952
rect 23900 16940 23906 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 6822 16736 6828 16788
rect 6880 16736 6886 16788
rect 7285 16779 7343 16785
rect 7285 16745 7297 16779
rect 7331 16776 7343 16779
rect 7466 16776 7472 16788
rect 7331 16748 7472 16776
rect 7331 16745 7343 16748
rect 7285 16739 7343 16745
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 9674 16776 9680 16788
rect 9600 16748 9680 16776
rect 7745 16711 7803 16717
rect 7745 16677 7757 16711
rect 7791 16708 7803 16711
rect 9306 16708 9312 16720
rect 7791 16680 9312 16708
rect 7791 16677 7803 16680
rect 7745 16671 7803 16677
rect 9306 16668 9312 16680
rect 9364 16668 9370 16720
rect 9493 16711 9551 16717
rect 9493 16677 9505 16711
rect 9539 16708 9551 16711
rect 9600 16708 9628 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 11238 16736 11244 16788
rect 11296 16776 11302 16788
rect 14734 16776 14740 16788
rect 11296 16748 14740 16776
rect 11296 16736 11302 16748
rect 14734 16736 14740 16748
rect 14792 16736 14798 16788
rect 16022 16736 16028 16788
rect 16080 16736 16086 16788
rect 16485 16779 16543 16785
rect 16485 16745 16497 16779
rect 16531 16776 16543 16779
rect 16666 16776 16672 16788
rect 16531 16748 16672 16776
rect 16531 16745 16543 16748
rect 16485 16739 16543 16745
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 19444 16748 21496 16776
rect 9539 16680 9628 16708
rect 9692 16680 10088 16708
rect 9539 16677 9551 16680
rect 9493 16671 9551 16677
rect 5258 16600 5264 16652
rect 5316 16600 5322 16652
rect 7469 16643 7527 16649
rect 7469 16609 7481 16643
rect 7515 16640 7527 16643
rect 8662 16640 8668 16652
rect 7515 16612 8668 16640
rect 7515 16609 7527 16612
rect 7469 16603 7527 16609
rect 4893 16575 4951 16581
rect 4893 16541 4905 16575
rect 4939 16572 4951 16575
rect 5276 16572 5304 16600
rect 7944 16581 7972 16612
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 9033 16643 9091 16649
rect 9033 16609 9045 16643
rect 9079 16640 9091 16643
rect 9582 16640 9588 16652
rect 9079 16612 9588 16640
rect 9079 16609 9091 16612
rect 9033 16603 9091 16609
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 4939 16544 5304 16572
rect 7929 16575 7987 16581
rect 4939 16541 4951 16544
rect 4893 16535 4951 16541
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 8570 16532 8576 16584
rect 8628 16568 8634 16584
rect 9692 16581 9720 16680
rect 10060 16640 10088 16680
rect 10134 16668 10140 16720
rect 10192 16708 10198 16720
rect 11974 16708 11980 16720
rect 10192 16680 11980 16708
rect 10192 16668 10198 16680
rect 11974 16668 11980 16680
rect 12032 16668 12038 16720
rect 13262 16668 13268 16720
rect 13320 16708 13326 16720
rect 13906 16708 13912 16720
rect 13320 16680 13912 16708
rect 13320 16668 13326 16680
rect 13906 16668 13912 16680
rect 13964 16668 13970 16720
rect 11330 16640 11336 16652
rect 10060 16612 11336 16640
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 11425 16643 11483 16649
rect 11425 16609 11437 16643
rect 11471 16640 11483 16643
rect 11606 16640 11612 16652
rect 11471 16612 11612 16640
rect 11471 16609 11483 16612
rect 11425 16603 11483 16609
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 12253 16643 12311 16649
rect 12253 16609 12265 16643
rect 12299 16640 12311 16643
rect 13722 16640 13728 16652
rect 12299 16612 13728 16640
rect 12299 16609 12311 16612
rect 12253 16603 12311 16609
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 14277 16643 14335 16649
rect 14277 16609 14289 16643
rect 14323 16640 14335 16643
rect 14918 16640 14924 16652
rect 14323 16612 14924 16640
rect 14323 16609 14335 16612
rect 14277 16603 14335 16609
rect 14918 16600 14924 16612
rect 14976 16600 14982 16652
rect 19444 16649 19472 16748
rect 17405 16643 17463 16649
rect 17405 16609 17417 16643
rect 17451 16640 17463 16643
rect 19429 16643 19487 16649
rect 17451 16612 19334 16640
rect 17451 16609 17463 16612
rect 17405 16603 17463 16609
rect 9677 16575 9735 16581
rect 8628 16540 8669 16568
rect 9677 16541 9689 16575
rect 9723 16541 9735 16575
rect 8628 16532 8634 16540
rect 9677 16535 9735 16541
rect 10870 16532 10876 16584
rect 10928 16572 10934 16584
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 10928 16544 11161 16572
rect 10928 16532 10934 16544
rect 11149 16541 11161 16544
rect 11195 16541 11207 16575
rect 11149 16535 11207 16541
rect 11238 16532 11244 16584
rect 11296 16532 11302 16584
rect 11698 16532 11704 16584
rect 11756 16572 11762 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11756 16544 11989 16572
rect 11756 16532 11762 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 16669 16575 16727 16581
rect 16669 16541 16681 16575
rect 16715 16541 16727 16575
rect 16669 16535 16727 16541
rect 8573 16531 8631 16532
rect 9217 16507 9275 16513
rect 9217 16473 9229 16507
rect 9263 16504 9275 16507
rect 9263 16476 9904 16504
rect 9263 16473 9275 16476
rect 9217 16467 9275 16473
rect 9876 16448 9904 16476
rect 12526 16464 12532 16516
rect 12584 16504 12590 16516
rect 14553 16507 14611 16513
rect 12584 16476 12742 16504
rect 12584 16464 12590 16476
rect 14553 16473 14565 16507
rect 14599 16504 14611 16507
rect 14826 16504 14832 16516
rect 14599 16476 14832 16504
rect 14599 16473 14611 16476
rect 14553 16467 14611 16473
rect 14826 16464 14832 16476
rect 14884 16464 14890 16516
rect 15010 16464 15016 16516
rect 15068 16464 15074 16516
rect 16684 16504 16712 16535
rect 17126 16532 17132 16584
rect 17184 16532 17190 16584
rect 17402 16504 17408 16516
rect 16684 16476 17408 16504
rect 17402 16464 17408 16476
rect 17460 16464 17466 16516
rect 17678 16464 17684 16516
rect 17736 16504 17742 16516
rect 19306 16504 19334 16612
rect 19429 16609 19441 16643
rect 19475 16609 19487 16643
rect 21468 16640 21496 16748
rect 22186 16736 22192 16788
rect 22244 16776 22250 16788
rect 23290 16776 23296 16788
rect 22244 16748 23296 16776
rect 22244 16736 22250 16748
rect 23290 16736 23296 16748
rect 23348 16736 23354 16788
rect 22278 16640 22284 16652
rect 21468 16612 22284 16640
rect 19429 16603 19487 16609
rect 22278 16600 22284 16612
rect 22336 16600 22342 16652
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16640 22615 16643
rect 22646 16640 22652 16652
rect 22603 16612 22652 16640
rect 22603 16609 22615 16612
rect 22557 16603 22615 16609
rect 22646 16600 22652 16612
rect 22704 16600 22710 16652
rect 24857 16643 24915 16649
rect 24857 16609 24869 16643
rect 24903 16640 24915 16643
rect 25590 16640 25596 16652
rect 24903 16612 25596 16640
rect 24903 16609 24915 16612
rect 24857 16603 24915 16609
rect 25590 16600 25596 16612
rect 25648 16600 25654 16652
rect 19426 16504 19432 16516
rect 17736 16476 17894 16504
rect 19306 16476 19432 16504
rect 17736 16464 17742 16476
rect 19426 16464 19432 16476
rect 19484 16464 19490 16516
rect 19702 16464 19708 16516
rect 19760 16464 19766 16516
rect 20162 16464 20168 16516
rect 20220 16464 20226 16516
rect 23842 16504 23848 16516
rect 23782 16476 23848 16504
rect 23842 16464 23848 16476
rect 23900 16464 23906 16516
rect 23934 16464 23940 16516
rect 23992 16504 23998 16516
rect 24673 16507 24731 16513
rect 24673 16504 24685 16507
rect 23992 16476 24685 16504
rect 23992 16464 23998 16476
rect 24673 16473 24685 16476
rect 24719 16473 24731 16507
rect 24673 16467 24731 16473
rect 4706 16396 4712 16448
rect 4764 16396 4770 16448
rect 8389 16439 8447 16445
rect 8389 16405 8401 16439
rect 8435 16436 8447 16439
rect 9766 16436 9772 16448
rect 8435 16408 9772 16436
rect 8435 16405 8447 16408
rect 8389 16399 8447 16405
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 9858 16396 9864 16448
rect 9916 16396 9922 16448
rect 10134 16396 10140 16448
rect 10192 16396 10198 16448
rect 10778 16396 10784 16448
rect 10836 16396 10842 16448
rect 11146 16396 11152 16448
rect 11204 16436 11210 16448
rect 11790 16436 11796 16448
rect 11204 16408 11796 16436
rect 11204 16396 11210 16408
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 12158 16436 12164 16448
rect 12032 16408 12164 16436
rect 12032 16396 12038 16408
rect 12158 16396 12164 16408
rect 12216 16436 12222 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 12216 16408 13737 16436
rect 12216 16396 12222 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 13725 16399 13783 16405
rect 17218 16396 17224 16448
rect 17276 16436 17282 16448
rect 18877 16439 18935 16445
rect 18877 16436 18889 16439
rect 17276 16408 18889 16436
rect 17276 16396 17282 16408
rect 18877 16405 18889 16408
rect 18923 16405 18935 16439
rect 18877 16399 18935 16405
rect 19242 16396 19248 16448
rect 19300 16436 19306 16448
rect 21177 16439 21235 16445
rect 21177 16436 21189 16439
rect 19300 16408 21189 16436
rect 19300 16396 19306 16408
rect 21177 16405 21189 16408
rect 21223 16436 21235 16439
rect 21266 16436 21272 16448
rect 21223 16408 21272 16436
rect 21223 16405 21235 16408
rect 21177 16399 21235 16405
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 21634 16396 21640 16448
rect 21692 16396 21698 16448
rect 23290 16396 23296 16448
rect 23348 16436 23354 16448
rect 24029 16439 24087 16445
rect 24029 16436 24041 16439
rect 23348 16408 24041 16436
rect 23348 16396 23354 16408
rect 24029 16405 24041 16408
rect 24075 16405 24087 16439
rect 24029 16399 24087 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 7834 16192 7840 16244
rect 7892 16232 7898 16244
rect 8113 16235 8171 16241
rect 8113 16232 8125 16235
rect 7892 16204 8125 16232
rect 7892 16192 7898 16204
rect 8113 16201 8125 16204
rect 8159 16201 8171 16235
rect 8113 16195 8171 16201
rect 8202 16192 8208 16244
rect 8260 16232 8266 16244
rect 8260 16204 9720 16232
rect 8260 16192 8266 16204
rect 4706 16124 4712 16176
rect 4764 16164 4770 16176
rect 9490 16164 9496 16176
rect 4764 16136 9496 16164
rect 4764 16124 4770 16136
rect 9490 16124 9496 16136
rect 9548 16124 9554 16176
rect 9692 16164 9720 16204
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 10781 16235 10839 16241
rect 10781 16232 10793 16235
rect 10192 16204 10793 16232
rect 10192 16192 10198 16204
rect 10781 16201 10793 16204
rect 10827 16201 10839 16235
rect 10781 16195 10839 16201
rect 10873 16235 10931 16241
rect 10873 16201 10885 16235
rect 10919 16232 10931 16235
rect 14369 16235 14427 16241
rect 10919 16204 13676 16232
rect 10919 16201 10931 16204
rect 10873 16195 10931 16201
rect 9692 16136 10640 16164
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 8202 16096 8208 16108
rect 7800 16068 8208 16096
rect 7800 16056 7806 16068
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 8389 16099 8447 16105
rect 8389 16065 8401 16099
rect 8435 16096 8447 16099
rect 8662 16096 8668 16108
rect 8435 16068 8668 16096
rect 8435 16065 8447 16068
rect 8389 16059 8447 16065
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 9309 16099 9367 16105
rect 9309 16065 9321 16099
rect 9355 16096 9367 16099
rect 9582 16096 9588 16108
rect 9355 16068 9588 16096
rect 9355 16065 9367 16068
rect 9309 16059 9367 16065
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 9858 16056 9864 16108
rect 9916 16096 9922 16108
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 9916 16068 9965 16096
rect 9916 16056 9922 16068
rect 9953 16065 9965 16068
rect 9999 16096 10011 16099
rect 10612 16096 10640 16136
rect 10686 16124 10692 16176
rect 10744 16164 10750 16176
rect 11882 16164 11888 16176
rect 10744 16136 11888 16164
rect 10744 16124 10750 16136
rect 11882 16124 11888 16136
rect 11940 16124 11946 16176
rect 11974 16124 11980 16176
rect 12032 16124 12038 16176
rect 12526 16124 12532 16176
rect 12584 16124 12590 16176
rect 9999 16068 10548 16096
rect 10612 16068 11652 16096
rect 9999 16065 10011 16068
rect 9953 16059 10011 16065
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 10520 16028 10548 16068
rect 10962 16028 10968 16040
rect 7340 16000 10456 16028
rect 10520 16000 10968 16028
rect 7340 15988 7346 16000
rect 6270 15920 6276 15972
rect 6328 15960 6334 15972
rect 6328 15932 9076 15960
rect 6328 15920 6334 15932
rect 8478 15852 8484 15904
rect 8536 15852 8542 15904
rect 9048 15892 9076 15932
rect 9122 15920 9128 15972
rect 9180 15920 9186 15972
rect 9769 15963 9827 15969
rect 9769 15929 9781 15963
rect 9815 15960 9827 15963
rect 10318 15960 10324 15972
rect 9815 15932 10324 15960
rect 9815 15929 9827 15932
rect 9769 15923 9827 15929
rect 10318 15920 10324 15932
rect 10376 15920 10382 15972
rect 10428 15969 10456 16000
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 10413 15963 10471 15969
rect 10413 15929 10425 15963
rect 10459 15929 10471 15963
rect 10413 15923 10471 15929
rect 10778 15892 10784 15904
rect 9048 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 11072 15892 11100 15991
rect 11624 15960 11652 16068
rect 11698 15988 11704 16040
rect 11756 15988 11762 16040
rect 12342 16028 12348 16040
rect 11808 16000 12348 16028
rect 11808 15960 11836 16000
rect 12342 15988 12348 16000
rect 12400 15988 12406 16040
rect 12710 15988 12716 16040
rect 12768 16028 12774 16040
rect 13446 16028 13452 16040
rect 12768 16000 13452 16028
rect 12768 15988 12774 16000
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 11624 15932 11836 15960
rect 13648 15960 13676 16204
rect 14369 16201 14381 16235
rect 14415 16232 14427 16235
rect 19337 16235 19395 16241
rect 19337 16232 19349 16235
rect 14415 16204 19349 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 19337 16201 19349 16204
rect 19383 16201 19395 16235
rect 19337 16195 19395 16201
rect 19426 16192 19432 16244
rect 19484 16232 19490 16244
rect 20070 16232 20076 16244
rect 19484 16204 20076 16232
rect 19484 16192 19490 16204
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 20438 16192 20444 16244
rect 20496 16232 20502 16244
rect 20993 16235 21051 16241
rect 20993 16232 21005 16235
rect 20496 16204 21005 16232
rect 20496 16192 20502 16204
rect 20993 16201 21005 16204
rect 21039 16201 21051 16235
rect 20993 16195 21051 16201
rect 23658 16192 23664 16244
rect 23716 16232 23722 16244
rect 23845 16235 23903 16241
rect 23845 16232 23857 16235
rect 23716 16204 23857 16232
rect 23716 16192 23722 16204
rect 23845 16201 23857 16204
rect 23891 16201 23903 16235
rect 23845 16195 23903 16201
rect 15746 16124 15752 16176
rect 15804 16164 15810 16176
rect 15933 16167 15991 16173
rect 15933 16164 15945 16167
rect 15804 16136 15945 16164
rect 15804 16124 15810 16136
rect 15933 16133 15945 16136
rect 15979 16133 15991 16167
rect 15933 16127 15991 16133
rect 19150 16124 19156 16176
rect 19208 16164 19214 16176
rect 19797 16167 19855 16173
rect 19797 16164 19809 16167
rect 19208 16136 19809 16164
rect 19208 16124 19214 16136
rect 19797 16133 19809 16136
rect 19843 16133 19855 16167
rect 19797 16127 19855 16133
rect 20898 16124 20904 16176
rect 20956 16124 20962 16176
rect 22373 16167 22431 16173
rect 22373 16133 22385 16167
rect 22419 16164 22431 16167
rect 24026 16164 24032 16176
rect 22419 16136 24032 16164
rect 22419 16133 22431 16136
rect 22373 16127 22431 16133
rect 24026 16124 24032 16136
rect 24084 16124 24090 16176
rect 24670 16124 24676 16176
rect 24728 16124 24734 16176
rect 13998 16056 14004 16108
rect 14056 16096 14062 16108
rect 14277 16099 14335 16105
rect 14277 16096 14289 16099
rect 14056 16068 14289 16096
rect 14056 16056 14062 16068
rect 14277 16065 14289 16068
rect 14323 16065 14335 16099
rect 14277 16059 14335 16065
rect 15841 16099 15899 16105
rect 15841 16065 15853 16099
rect 15887 16096 15899 16099
rect 16206 16096 16212 16108
rect 15887 16068 16212 16096
rect 15887 16065 15899 16068
rect 15841 16059 15899 16065
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 19058 16096 19064 16108
rect 17175 16068 19064 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 19702 16056 19708 16108
rect 19760 16056 19766 16108
rect 20162 16096 20168 16108
rect 19812 16068 20168 16096
rect 14550 15988 14556 16040
rect 14608 15988 14614 16040
rect 15194 15988 15200 16040
rect 15252 16028 15258 16040
rect 16025 16031 16083 16037
rect 16025 16028 16037 16031
rect 15252 16000 16037 16028
rect 15252 15988 15258 16000
rect 16025 15997 16037 16000
rect 16071 15997 16083 16031
rect 16025 15991 16083 15997
rect 18966 15988 18972 16040
rect 19024 16028 19030 16040
rect 19812 16028 19840 16068
rect 20162 16056 20168 16068
rect 20220 16096 20226 16108
rect 21450 16096 21456 16108
rect 20220 16068 21456 16096
rect 20220 16056 20226 16068
rect 21450 16056 21456 16068
rect 21508 16096 21514 16108
rect 21545 16099 21603 16105
rect 21545 16096 21557 16099
rect 21508 16068 21557 16096
rect 21508 16056 21514 16068
rect 21545 16065 21557 16068
rect 21591 16065 21603 16099
rect 21545 16059 21603 16065
rect 23753 16099 23811 16105
rect 23753 16065 23765 16099
rect 23799 16096 23811 16099
rect 24578 16096 24584 16108
rect 23799 16068 24584 16096
rect 23799 16065 23811 16068
rect 23753 16059 23811 16065
rect 24578 16056 24584 16068
rect 24636 16056 24642 16108
rect 19024 16000 19840 16028
rect 19889 16031 19947 16037
rect 19024 15988 19030 16000
rect 19889 15997 19901 16031
rect 19935 15997 19947 16031
rect 19889 15991 19947 15997
rect 15473 15963 15531 15969
rect 15473 15960 15485 15963
rect 13648 15932 15485 15960
rect 15473 15929 15485 15932
rect 15519 15929 15531 15963
rect 15473 15923 15531 15929
rect 17494 15920 17500 15972
rect 17552 15960 17558 15972
rect 19904 15960 19932 15991
rect 21082 15988 21088 16040
rect 21140 15988 21146 16040
rect 21726 15988 21732 16040
rect 21784 16028 21790 16040
rect 22465 16031 22523 16037
rect 22465 16028 22477 16031
rect 21784 16000 22477 16028
rect 21784 15988 21790 16000
rect 22465 15997 22477 16000
rect 22511 15997 22523 16031
rect 22465 15991 22523 15997
rect 22554 15988 22560 16040
rect 22612 15988 22618 16040
rect 23937 16031 23995 16037
rect 23937 15997 23949 16031
rect 23983 15997 23995 16031
rect 23937 15991 23995 15997
rect 17552 15932 19932 15960
rect 17552 15920 17558 15932
rect 20070 15920 20076 15972
rect 20128 15960 20134 15972
rect 22738 15960 22744 15972
rect 20128 15932 22744 15960
rect 20128 15920 20134 15932
rect 22738 15920 22744 15932
rect 22796 15960 22802 15972
rect 23017 15963 23075 15969
rect 23017 15960 23029 15963
rect 22796 15932 23029 15960
rect 22796 15920 22802 15932
rect 23017 15929 23029 15932
rect 23063 15929 23075 15963
rect 23017 15923 23075 15929
rect 23290 15920 23296 15972
rect 23348 15960 23354 15972
rect 23952 15960 23980 15991
rect 23348 15932 23980 15960
rect 24857 15963 24915 15969
rect 23348 15920 23354 15932
rect 24857 15929 24869 15963
rect 24903 15960 24915 15963
rect 25038 15960 25044 15972
rect 24903 15932 25044 15960
rect 24903 15929 24915 15932
rect 24857 15923 24915 15929
rect 25038 15920 25044 15932
rect 25096 15920 25102 15972
rect 12066 15892 12072 15904
rect 11072 15864 12072 15892
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 13906 15852 13912 15904
rect 13964 15852 13970 15904
rect 15010 15852 15016 15904
rect 15068 15892 15074 15904
rect 16298 15892 16304 15904
rect 15068 15864 16304 15892
rect 15068 15852 15074 15864
rect 16298 15852 16304 15864
rect 16356 15892 16362 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 16356 15864 16681 15892
rect 16356 15852 16362 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 17862 15852 17868 15904
rect 17920 15892 17926 15904
rect 18417 15895 18475 15901
rect 18417 15892 18429 15895
rect 17920 15864 18429 15892
rect 17920 15852 17926 15864
rect 18417 15861 18429 15864
rect 18463 15892 18475 15895
rect 18874 15892 18880 15904
rect 18463 15864 18880 15892
rect 18463 15861 18475 15864
rect 18417 15855 18475 15861
rect 18874 15852 18880 15864
rect 18932 15852 18938 15904
rect 20530 15852 20536 15904
rect 20588 15852 20594 15904
rect 22005 15895 22063 15901
rect 22005 15861 22017 15895
rect 22051 15892 22063 15895
rect 22370 15892 22376 15904
rect 22051 15864 22376 15892
rect 22051 15861 22063 15864
rect 22005 15855 22063 15861
rect 22370 15852 22376 15864
rect 22428 15852 22434 15904
rect 22554 15852 22560 15904
rect 22612 15892 22618 15904
rect 23385 15895 23443 15901
rect 23385 15892 23397 15895
rect 22612 15864 23397 15892
rect 22612 15852 22618 15864
rect 23385 15861 23397 15864
rect 23431 15861 23443 15895
rect 23385 15855 23443 15861
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 8754 15648 8760 15700
rect 8812 15648 8818 15700
rect 9861 15691 9919 15697
rect 9861 15657 9873 15691
rect 9907 15688 9919 15691
rect 9907 15660 11836 15688
rect 9907 15657 9919 15660
rect 9861 15651 9919 15657
rect 11808 15620 11836 15660
rect 11882 15648 11888 15700
rect 11940 15688 11946 15700
rect 13906 15688 13912 15700
rect 11940 15660 13912 15688
rect 11940 15648 11946 15660
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 16850 15688 16856 15700
rect 14016 15660 16856 15688
rect 14016 15620 14044 15660
rect 16850 15648 16856 15660
rect 16908 15648 16914 15700
rect 18693 15691 18751 15697
rect 18693 15688 18705 15691
rect 17052 15660 18705 15688
rect 11808 15592 13032 15620
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15552 10839 15555
rect 12710 15552 12716 15564
rect 10827 15524 12716 15552
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 12710 15512 12716 15524
rect 12768 15512 12774 15564
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15484 9459 15487
rect 9490 15484 9496 15496
rect 9447 15456 9496 15484
rect 9447 15453 9459 15456
rect 9401 15447 9459 15453
rect 9490 15444 9496 15456
rect 9548 15484 9554 15496
rect 9950 15484 9956 15496
rect 9548 15456 9956 15484
rect 9548 15444 9554 15456
rect 9950 15444 9956 15456
rect 10008 15444 10014 15496
rect 10042 15444 10048 15496
rect 10100 15444 10106 15496
rect 10505 15487 10563 15493
rect 10505 15453 10517 15487
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 10520 15416 10548 15447
rect 10686 15416 10692 15428
rect 10520 15388 10692 15416
rect 10686 15376 10692 15388
rect 10744 15376 10750 15428
rect 12526 15416 12532 15428
rect 12006 15388 12532 15416
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 13004 15416 13032 15592
rect 13188 15592 14044 15620
rect 13188 15561 13216 15592
rect 15838 15580 15844 15632
rect 15896 15620 15902 15632
rect 16025 15623 16083 15629
rect 16025 15620 16037 15623
rect 15896 15592 16037 15620
rect 15896 15580 15902 15592
rect 16025 15589 16037 15592
rect 16071 15589 16083 15623
rect 16025 15583 16083 15589
rect 16298 15580 16304 15632
rect 16356 15580 16362 15632
rect 16758 15580 16764 15632
rect 16816 15620 16822 15632
rect 17052 15620 17080 15660
rect 18693 15657 18705 15660
rect 18739 15688 18751 15691
rect 19334 15688 19340 15700
rect 18739 15660 19340 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 20530 15648 20536 15700
rect 20588 15688 20594 15700
rect 25406 15688 25412 15700
rect 20588 15660 25412 15688
rect 20588 15648 20594 15660
rect 25406 15648 25412 15660
rect 25464 15648 25470 15700
rect 16816 15592 17080 15620
rect 16816 15580 16822 15592
rect 18598 15580 18604 15632
rect 18656 15620 18662 15632
rect 18656 15592 21864 15620
rect 18656 15580 18662 15592
rect 13173 15555 13231 15561
rect 13173 15521 13185 15555
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 14182 15552 14188 15564
rect 13403 15524 14188 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 14274 15512 14280 15564
rect 14332 15552 14338 15564
rect 16945 15555 17003 15561
rect 16945 15552 16957 15555
rect 14332 15524 16957 15552
rect 14332 15512 14338 15524
rect 16945 15521 16957 15524
rect 16991 15521 17003 15555
rect 16945 15515 17003 15521
rect 17218 15512 17224 15564
rect 17276 15552 17282 15564
rect 20073 15555 20131 15561
rect 20073 15552 20085 15555
rect 17276 15524 20085 15552
rect 17276 15512 17282 15524
rect 20073 15521 20085 15524
rect 20119 15521 20131 15555
rect 20073 15515 20131 15521
rect 21174 15512 21180 15564
rect 21232 15512 21238 15564
rect 21266 15512 21272 15564
rect 21324 15512 21330 15564
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13814 15484 13820 15496
rect 13127 15456 13820 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 19978 15444 19984 15496
rect 20036 15444 20042 15496
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15484 21143 15487
rect 21836 15484 21864 15592
rect 22189 15555 22247 15561
rect 22189 15521 22201 15555
rect 22235 15552 22247 15555
rect 25774 15552 25780 15564
rect 22235 15524 25780 15552
rect 22235 15521 22247 15524
rect 22189 15515 22247 15521
rect 25774 15512 25780 15524
rect 25832 15512 25838 15564
rect 22005 15487 22063 15493
rect 22005 15484 22017 15487
rect 21131 15456 21772 15484
rect 21836 15456 22017 15484
rect 21131 15453 21143 15456
rect 21085 15447 21143 15453
rect 14458 15416 14464 15428
rect 13004 15388 14464 15416
rect 14458 15376 14464 15388
rect 14516 15376 14522 15428
rect 14553 15419 14611 15425
rect 14553 15385 14565 15419
rect 14599 15385 14611 15419
rect 14553 15379 14611 15385
rect 9217 15351 9275 15357
rect 9217 15317 9229 15351
rect 9263 15348 9275 15351
rect 11146 15348 11152 15360
rect 9263 15320 11152 15348
rect 9263 15317 9275 15320
rect 9217 15311 9275 15317
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 11606 15308 11612 15360
rect 11664 15348 11670 15360
rect 12253 15351 12311 15357
rect 12253 15348 12265 15351
rect 11664 15320 12265 15348
rect 11664 15308 11670 15320
rect 12253 15317 12265 15320
rect 12299 15317 12311 15351
rect 12253 15311 12311 15317
rect 12342 15308 12348 15360
rect 12400 15348 12406 15360
rect 12713 15351 12771 15357
rect 12713 15348 12725 15351
rect 12400 15320 12725 15348
rect 12400 15308 12406 15320
rect 12713 15317 12725 15320
rect 12759 15317 12771 15351
rect 12713 15311 12771 15317
rect 13817 15351 13875 15357
rect 13817 15317 13829 15351
rect 13863 15348 13875 15351
rect 13906 15348 13912 15360
rect 13863 15320 13912 15348
rect 13863 15317 13875 15320
rect 13817 15311 13875 15317
rect 13906 15308 13912 15320
rect 13964 15308 13970 15360
rect 14568 15348 14596 15379
rect 15010 15376 15016 15428
rect 15068 15376 15074 15428
rect 16574 15416 16580 15428
rect 15856 15388 16580 15416
rect 15856 15348 15884 15388
rect 16574 15376 16580 15388
rect 16632 15376 16638 15428
rect 16669 15419 16727 15425
rect 16669 15385 16681 15419
rect 16715 15416 16727 15419
rect 17310 15416 17316 15428
rect 16715 15388 17316 15416
rect 16715 15385 16727 15388
rect 16669 15379 16727 15385
rect 17310 15376 17316 15388
rect 17368 15376 17374 15428
rect 17678 15416 17684 15428
rect 17420 15388 17684 15416
rect 14568 15320 15884 15348
rect 17218 15308 17224 15360
rect 17276 15348 17282 15360
rect 17420 15348 17448 15388
rect 17678 15376 17684 15388
rect 17736 15376 17742 15428
rect 19889 15419 19947 15425
rect 19889 15385 19901 15419
rect 19935 15416 19947 15419
rect 21634 15416 21640 15428
rect 19935 15388 21640 15416
rect 19935 15385 19947 15388
rect 19889 15379 19947 15385
rect 21634 15376 21640 15388
rect 21692 15376 21698 15428
rect 18966 15348 18972 15360
rect 17276 15320 18972 15348
rect 17276 15308 17282 15320
rect 18966 15308 18972 15320
rect 19024 15308 19030 15360
rect 19521 15351 19579 15357
rect 19521 15317 19533 15351
rect 19567 15348 19579 15351
rect 20530 15348 20536 15360
rect 19567 15320 20536 15348
rect 19567 15317 19579 15320
rect 19521 15311 19579 15317
rect 20530 15308 20536 15320
rect 20588 15308 20594 15360
rect 20717 15351 20775 15357
rect 20717 15317 20729 15351
rect 20763 15348 20775 15351
rect 21358 15348 21364 15360
rect 20763 15320 21364 15348
rect 20763 15317 20775 15320
rect 20717 15311 20775 15317
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 21744 15348 21772 15456
rect 22005 15453 22017 15456
rect 22051 15453 22063 15487
rect 23385 15487 23443 15493
rect 23385 15484 23397 15487
rect 22005 15447 22063 15453
rect 22112 15456 23397 15484
rect 22112 15416 22140 15456
rect 23385 15453 23397 15456
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 23750 15444 23756 15496
rect 23808 15484 23814 15496
rect 24765 15487 24823 15493
rect 24765 15484 24777 15487
rect 23808 15456 24777 15484
rect 23808 15444 23814 15456
rect 24765 15453 24777 15456
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 22066 15388 22140 15416
rect 22066 15348 22094 15388
rect 22738 15376 22744 15428
rect 22796 15376 22802 15428
rect 21744 15320 22094 15348
rect 22830 15308 22836 15360
rect 22888 15308 22894 15360
rect 23474 15308 23480 15360
rect 23532 15348 23538 15360
rect 24581 15351 24639 15357
rect 24581 15348 24593 15351
rect 23532 15320 24593 15348
rect 23532 15308 23538 15320
rect 24581 15317 24593 15320
rect 24627 15317 24639 15351
rect 24581 15311 24639 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 5534 15144 5540 15156
rect 4120 15116 5540 15144
rect 4120 15104 4126 15116
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 9490 15104 9496 15156
rect 9548 15104 9554 15156
rect 9677 15147 9735 15153
rect 9677 15113 9689 15147
rect 9723 15144 9735 15147
rect 10042 15144 10048 15156
rect 9723 15116 10048 15144
rect 9723 15113 9735 15116
rect 9677 15107 9735 15113
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 10321 15147 10379 15153
rect 10321 15113 10333 15147
rect 10367 15144 10379 15147
rect 14918 15144 14924 15156
rect 10367 15116 14924 15144
rect 10367 15113 10379 15116
rect 10321 15107 10379 15113
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 18874 15144 18880 15156
rect 16132 15116 18880 15144
rect 9861 15079 9919 15085
rect 9861 15045 9873 15079
rect 9907 15076 9919 15079
rect 9907 15048 11192 15076
rect 9907 15045 9919 15048
rect 9861 15039 9919 15045
rect 11164 15020 11192 15048
rect 12526 15036 12532 15088
rect 12584 15036 12590 15088
rect 13909 15079 13967 15085
rect 13909 15045 13921 15079
rect 13955 15076 13967 15079
rect 13998 15076 14004 15088
rect 13955 15048 14004 15076
rect 13955 15045 13967 15048
rect 13909 15039 13967 15045
rect 13998 15036 14004 15048
rect 14056 15036 14062 15088
rect 14108 15048 15240 15076
rect 10502 14968 10508 15020
rect 10560 14968 10566 15020
rect 11146 14968 11152 15020
rect 11204 14968 11210 15020
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 14108 15008 14136 15048
rect 13872 14980 14136 15008
rect 14553 15011 14611 15017
rect 13872 14968 13878 14980
rect 14553 14977 14565 15011
rect 14599 15008 14611 15011
rect 15013 15011 15071 15017
rect 15013 15008 15025 15011
rect 14599 14980 15025 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 15013 14977 15025 14980
rect 15059 15008 15071 15011
rect 15102 15008 15108 15020
rect 15059 14980 15108 15008
rect 15059 14977 15071 14980
rect 15013 14971 15071 14977
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 15212 15008 15240 15048
rect 15378 15036 15384 15088
rect 15436 15076 15442 15088
rect 16132 15085 16160 15116
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 19150 15104 19156 15156
rect 19208 15144 19214 15156
rect 22462 15144 22468 15156
rect 19208 15116 22468 15144
rect 19208 15104 19214 15116
rect 22462 15104 22468 15116
rect 22520 15104 22526 15156
rect 23290 15144 23296 15156
rect 23124 15116 23296 15144
rect 15473 15079 15531 15085
rect 15473 15076 15485 15079
rect 15436 15048 15485 15076
rect 15436 15036 15442 15048
rect 15473 15045 15485 15048
rect 15519 15045 15531 15079
rect 15473 15039 15531 15045
rect 16117 15079 16175 15085
rect 16117 15045 16129 15079
rect 16163 15045 16175 15079
rect 16117 15039 16175 15045
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 17129 15079 17187 15085
rect 17129 15076 17141 15079
rect 16816 15048 17141 15076
rect 16816 15036 16822 15048
rect 17129 15045 17141 15048
rect 17175 15045 17187 15079
rect 17129 15039 17187 15045
rect 17218 15036 17224 15088
rect 17276 15076 17282 15088
rect 17276 15048 17618 15076
rect 17276 15036 17282 15048
rect 18966 15036 18972 15088
rect 19024 15076 19030 15088
rect 19024 15048 20102 15076
rect 19024 15036 19030 15048
rect 21450 15036 21456 15088
rect 21508 15036 21514 15088
rect 22094 15036 22100 15088
rect 22152 15036 22158 15088
rect 23124 15085 23152 15116
rect 23290 15104 23296 15116
rect 23348 15104 23354 15156
rect 24118 15104 24124 15156
rect 24176 15144 24182 15156
rect 24581 15147 24639 15153
rect 24581 15144 24593 15147
rect 24176 15116 24593 15144
rect 24176 15104 24182 15116
rect 24581 15113 24593 15116
rect 24627 15113 24639 15147
rect 24581 15107 24639 15113
rect 23109 15079 23167 15085
rect 23109 15045 23121 15079
rect 23155 15045 23167 15079
rect 23109 15039 23167 15045
rect 23658 15036 23664 15088
rect 23716 15036 23722 15088
rect 16482 15008 16488 15020
rect 15212 14980 16488 15008
rect 16482 14968 16488 14980
rect 16540 14968 16546 15020
rect 22186 15008 22192 15020
rect 20824 14980 22192 15008
rect 10045 14943 10103 14949
rect 10045 14909 10057 14943
rect 10091 14940 10103 14943
rect 10594 14940 10600 14952
rect 10091 14912 10600 14940
rect 10091 14909 10103 14912
rect 10045 14903 10103 14909
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 11698 14940 11704 14952
rect 10744 14912 11704 14940
rect 10744 14900 10750 14912
rect 11698 14900 11704 14912
rect 11756 14900 11762 14952
rect 11974 14900 11980 14952
rect 12032 14900 12038 14952
rect 12066 14900 12072 14952
rect 12124 14940 12130 14952
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 12124 14912 13461 14940
rect 12124 14900 12130 14912
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14940 16911 14943
rect 17126 14940 17132 14952
rect 16899 14912 17132 14940
rect 16899 14909 16911 14912
rect 16853 14903 16911 14909
rect 13630 14832 13636 14884
rect 13688 14872 13694 14884
rect 16666 14872 16672 14884
rect 13688 14844 16672 14872
rect 13688 14832 13694 14844
rect 16666 14832 16672 14844
rect 16724 14832 16730 14884
rect 10965 14807 11023 14813
rect 10965 14773 10977 14807
rect 11011 14804 11023 14807
rect 13446 14804 13452 14816
rect 11011 14776 13452 14804
rect 11011 14773 11023 14776
rect 10965 14767 11023 14773
rect 13446 14764 13452 14776
rect 13504 14764 13510 14816
rect 14826 14764 14832 14816
rect 14884 14764 14890 14816
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 16868 14804 16896 14903
rect 17126 14900 17132 14912
rect 17184 14940 17190 14952
rect 19334 14940 19340 14952
rect 17184 14912 19340 14940
rect 17184 14900 17190 14912
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14940 19671 14943
rect 19659 14912 20760 14940
rect 19659 14909 19671 14912
rect 19613 14903 19671 14909
rect 20732 14884 20760 14912
rect 18966 14832 18972 14884
rect 19024 14872 19030 14884
rect 19024 14844 19472 14872
rect 19024 14832 19030 14844
rect 16540 14776 16896 14804
rect 16540 14764 16546 14776
rect 18598 14764 18604 14816
rect 18656 14764 18662 14816
rect 19058 14764 19064 14816
rect 19116 14764 19122 14816
rect 19444 14804 19472 14844
rect 20714 14832 20720 14884
rect 20772 14832 20778 14884
rect 20824 14804 20852 14980
rect 22186 14968 22192 14980
rect 22244 14968 22250 15020
rect 21085 14943 21143 14949
rect 21085 14909 21097 14943
rect 21131 14940 21143 14943
rect 21818 14940 21824 14952
rect 21131 14912 21824 14940
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 21818 14900 21824 14912
rect 21876 14900 21882 14952
rect 22278 14900 22284 14952
rect 22336 14940 22342 14952
rect 22833 14943 22891 14949
rect 22833 14940 22845 14943
rect 22336 14912 22845 14940
rect 22336 14900 22342 14912
rect 22833 14909 22845 14912
rect 22879 14909 22891 14943
rect 25041 14943 25099 14949
rect 25041 14940 25053 14943
rect 22833 14903 22891 14909
rect 24136 14912 25053 14940
rect 21174 14832 21180 14884
rect 21232 14872 21238 14884
rect 21232 14844 22968 14872
rect 21232 14832 21238 14844
rect 19444 14776 20852 14804
rect 22189 14807 22247 14813
rect 22189 14773 22201 14807
rect 22235 14804 22247 14807
rect 22646 14804 22652 14816
rect 22235 14776 22652 14804
rect 22235 14773 22247 14776
rect 22189 14767 22247 14773
rect 22646 14764 22652 14776
rect 22704 14764 22710 14816
rect 22940 14804 22968 14844
rect 24136 14804 24164 14912
rect 25041 14909 25053 14912
rect 25087 14909 25099 14943
rect 25041 14903 25099 14909
rect 22940 14776 24164 14804
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 10413 14603 10471 14609
rect 10413 14569 10425 14603
rect 10459 14600 10471 14603
rect 10502 14600 10508 14612
rect 10459 14572 10508 14600
rect 10459 14569 10471 14572
rect 10413 14563 10471 14569
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 11146 14560 11152 14612
rect 11204 14600 11210 14612
rect 12897 14603 12955 14609
rect 11204 14572 12848 14600
rect 11204 14560 11210 14572
rect 12820 14532 12848 14572
rect 12897 14569 12909 14603
rect 12943 14600 12955 14603
rect 13630 14600 13636 14612
rect 12943 14572 13636 14600
rect 12943 14569 12955 14572
rect 12897 14563 12955 14569
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 14642 14600 14648 14612
rect 14200 14572 14648 14600
rect 13814 14532 13820 14544
rect 12820 14504 13820 14532
rect 13814 14492 13820 14504
rect 13872 14492 13878 14544
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 11606 14464 11612 14476
rect 11011 14436 11612 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 11606 14424 11612 14436
rect 11664 14424 11670 14476
rect 11974 14424 11980 14476
rect 12032 14464 12038 14476
rect 12437 14467 12495 14473
rect 12437 14464 12449 14467
rect 12032 14436 12449 14464
rect 12032 14424 12038 14436
rect 12437 14433 12449 14436
rect 12483 14433 12495 14467
rect 12437 14427 12495 14433
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 14200 14464 14228 14572
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 18966 14600 18972 14612
rect 14976 14572 18972 14600
rect 14976 14560 14982 14572
rect 18966 14560 18972 14572
rect 19024 14560 19030 14612
rect 19242 14560 19248 14612
rect 19300 14600 19306 14612
rect 19610 14600 19616 14612
rect 19300 14572 19616 14600
rect 19300 14560 19306 14572
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 20346 14560 20352 14612
rect 20404 14600 20410 14612
rect 20533 14603 20591 14609
rect 20533 14600 20545 14603
rect 20404 14572 20545 14600
rect 20404 14560 20410 14572
rect 20533 14569 20545 14572
rect 20579 14600 20591 14603
rect 21450 14600 21456 14612
rect 20579 14572 21456 14600
rect 20579 14569 20591 14572
rect 20533 14563 20591 14569
rect 21450 14560 21456 14572
rect 21508 14560 21514 14612
rect 22278 14560 22284 14612
rect 22336 14560 22342 14612
rect 22462 14560 22468 14612
rect 22520 14600 22526 14612
rect 24946 14600 24952 14612
rect 22520 14572 24952 14600
rect 22520 14560 22526 14572
rect 24946 14560 24952 14572
rect 25004 14560 25010 14612
rect 25130 14560 25136 14612
rect 25188 14600 25194 14612
rect 25409 14603 25467 14609
rect 25409 14600 25421 14603
rect 25188 14572 25421 14600
rect 25188 14560 25194 14572
rect 25409 14569 25421 14572
rect 25455 14600 25467 14603
rect 26142 14600 26148 14612
rect 25455 14572 26148 14600
rect 25455 14569 25467 14572
rect 25409 14563 25467 14569
rect 26142 14560 26148 14572
rect 26200 14560 26206 14612
rect 18233 14535 18291 14541
rect 18233 14501 18245 14535
rect 18279 14532 18291 14535
rect 18690 14532 18696 14544
rect 18279 14504 18696 14532
rect 18279 14501 18291 14504
rect 18233 14495 18291 14501
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 19429 14535 19487 14541
rect 18800 14504 19334 14532
rect 13587 14436 14228 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 12452 14328 12480 14427
rect 14274 14424 14280 14476
rect 14332 14424 14338 14476
rect 14550 14424 14556 14476
rect 14608 14424 14614 14476
rect 16482 14424 16488 14476
rect 16540 14424 16546 14476
rect 16761 14467 16819 14473
rect 16761 14433 16773 14467
rect 16807 14464 16819 14467
rect 18598 14464 18604 14476
rect 16807 14436 18604 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 18598 14424 18604 14436
rect 18656 14464 18662 14476
rect 18800 14464 18828 14504
rect 18656 14436 18828 14464
rect 19306 14464 19334 14504
rect 19429 14501 19441 14535
rect 19475 14532 19487 14535
rect 20898 14532 20904 14544
rect 19475 14504 20904 14532
rect 19475 14501 19487 14504
rect 19429 14495 19487 14501
rect 20898 14492 20904 14504
rect 20956 14492 20962 14544
rect 21468 14532 21496 14560
rect 22833 14535 22891 14541
rect 22833 14532 22845 14535
rect 21468 14504 22845 14532
rect 22833 14501 22845 14504
rect 22879 14532 22891 14535
rect 23658 14532 23664 14544
rect 22879 14504 23664 14532
rect 22879 14501 22891 14504
rect 22833 14495 22891 14501
rect 23658 14492 23664 14504
rect 23716 14532 23722 14544
rect 25225 14535 25283 14541
rect 25225 14532 25237 14535
rect 23716 14504 25237 14532
rect 23716 14492 23722 14504
rect 25225 14501 25237 14504
rect 25271 14501 25283 14535
rect 25225 14495 25283 14501
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19306 14436 19993 14464
rect 18656 14424 18662 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 23382 14424 23388 14476
rect 23440 14464 23446 14476
rect 23753 14467 23811 14473
rect 23753 14464 23765 14467
rect 23440 14436 23765 14464
rect 23440 14424 23446 14436
rect 23753 14433 23765 14436
rect 23799 14433 23811 14467
rect 23753 14427 23811 14433
rect 23937 14467 23995 14473
rect 23937 14433 23949 14467
rect 23983 14464 23995 14467
rect 24486 14464 24492 14476
rect 23983 14436 24492 14464
rect 23983 14433 23995 14436
rect 23937 14427 23995 14433
rect 24486 14424 24492 14436
rect 24544 14424 24550 14476
rect 13081 14399 13139 14405
rect 13081 14365 13093 14399
rect 13127 14396 13139 14399
rect 13906 14396 13912 14408
rect 13127 14368 13912 14396
rect 13127 14365 13139 14368
rect 13081 14359 13139 14365
rect 13906 14356 13912 14368
rect 13964 14356 13970 14408
rect 19150 14356 19156 14408
rect 19208 14372 19214 14408
rect 20809 14399 20867 14405
rect 20809 14396 20821 14399
rect 19306 14372 20821 14396
rect 19208 14368 20821 14372
rect 19208 14356 19334 14368
rect 20809 14365 20821 14368
rect 20855 14396 20867 14399
rect 22002 14396 22008 14408
rect 20855 14368 22008 14396
rect 20855 14365 20867 14368
rect 20809 14359 20867 14365
rect 22002 14356 22008 14368
rect 22060 14356 22066 14408
rect 23661 14399 23719 14405
rect 23661 14365 23673 14399
rect 23707 14396 23719 14399
rect 24854 14396 24860 14408
rect 23707 14368 24860 14396
rect 23707 14365 23719 14368
rect 23661 14359 23719 14365
rect 24854 14356 24860 14368
rect 24912 14356 24918 14408
rect 19168 14344 19334 14356
rect 12190 14300 12388 14328
rect 12452 14300 13676 14328
rect 12360 14260 12388 14300
rect 12526 14260 12532 14272
rect 12360 14232 12532 14260
rect 12526 14220 12532 14232
rect 12584 14220 12590 14272
rect 13648 14260 13676 14300
rect 15010 14288 15016 14340
rect 15068 14288 15074 14340
rect 17218 14288 17224 14340
rect 17276 14288 17282 14340
rect 19610 14288 19616 14340
rect 19668 14328 19674 14340
rect 19797 14331 19855 14337
rect 19797 14328 19809 14331
rect 19668 14300 19809 14328
rect 19668 14288 19674 14300
rect 19797 14297 19809 14300
rect 19843 14297 19855 14331
rect 19797 14291 19855 14297
rect 19886 14288 19892 14340
rect 19944 14288 19950 14340
rect 19978 14288 19984 14340
rect 20036 14328 20042 14340
rect 20036 14300 23336 14328
rect 20036 14288 20042 14300
rect 15194 14260 15200 14272
rect 13648 14232 15200 14260
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 16025 14263 16083 14269
rect 16025 14229 16037 14263
rect 16071 14260 16083 14263
rect 16574 14260 16580 14272
rect 16071 14232 16580 14260
rect 16071 14229 16083 14232
rect 16025 14223 16083 14229
rect 16574 14220 16580 14232
rect 16632 14220 16638 14272
rect 18693 14263 18751 14269
rect 18693 14229 18705 14263
rect 18739 14260 18751 14263
rect 18874 14260 18880 14272
rect 18739 14232 18880 14260
rect 18739 14229 18751 14232
rect 18693 14223 18751 14229
rect 18874 14220 18880 14232
rect 18932 14220 18938 14272
rect 19150 14220 19156 14272
rect 19208 14260 19214 14272
rect 22738 14260 22744 14272
rect 19208 14232 22744 14260
rect 19208 14220 19214 14232
rect 22738 14220 22744 14232
rect 22796 14220 22802 14272
rect 23308 14269 23336 14300
rect 24302 14288 24308 14340
rect 24360 14328 24366 14340
rect 24673 14331 24731 14337
rect 24673 14328 24685 14331
rect 24360 14300 24685 14328
rect 24360 14288 24366 14300
rect 24673 14297 24685 14300
rect 24719 14297 24731 14331
rect 24673 14291 24731 14297
rect 23293 14263 23351 14269
rect 23293 14229 23305 14263
rect 23339 14229 23351 14263
rect 23293 14223 23351 14229
rect 24118 14220 24124 14272
rect 24176 14260 24182 14272
rect 24765 14263 24823 14269
rect 24765 14260 24777 14263
rect 24176 14232 24777 14260
rect 24176 14220 24182 14232
rect 24765 14229 24777 14232
rect 24811 14229 24823 14263
rect 24765 14223 24823 14229
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 13722 14056 13728 14068
rect 11379 14028 13728 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11149 13991 11207 13997
rect 11149 13957 11161 13991
rect 11195 13988 11207 13991
rect 11514 13988 11520 14000
rect 11195 13960 11520 13988
rect 11195 13957 11207 13960
rect 11149 13951 11207 13957
rect 11514 13948 11520 13960
rect 11572 13988 11578 14000
rect 11572 13960 12020 13988
rect 11572 13948 11578 13960
rect 11992 13929 12020 13960
rect 12636 13929 12664 14028
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 14366 14056 14372 14068
rect 13872 14028 14372 14056
rect 13872 14016 13878 14028
rect 14366 14016 14372 14028
rect 14424 14016 14430 14068
rect 14642 14016 14648 14068
rect 14700 14056 14706 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 14700 14028 15485 14056
rect 14700 14016 14706 14028
rect 15473 14025 15485 14028
rect 15519 14025 15531 14059
rect 15473 14019 15531 14025
rect 16114 14016 16120 14068
rect 16172 14016 16178 14068
rect 17037 14059 17095 14065
rect 17037 14025 17049 14059
rect 17083 14056 17095 14059
rect 17126 14056 17132 14068
rect 17083 14028 17132 14056
rect 17083 14025 17095 14028
rect 17037 14019 17095 14025
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 17497 14059 17555 14065
rect 17497 14025 17509 14059
rect 17543 14056 17555 14059
rect 17586 14056 17592 14068
rect 17543 14028 17592 14056
rect 17543 14025 17555 14028
rect 17497 14019 17555 14025
rect 17586 14016 17592 14028
rect 17644 14016 17650 14068
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19392 14028 19533 14056
rect 19392 14016 19398 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20622 14056 20628 14068
rect 20404 14028 20628 14056
rect 20404 14016 20410 14028
rect 20622 14016 20628 14028
rect 20680 14016 20686 14068
rect 21085 14059 21143 14065
rect 21085 14025 21097 14059
rect 21131 14056 21143 14059
rect 21174 14056 21180 14068
rect 21131 14028 21180 14056
rect 21131 14025 21143 14028
rect 21085 14019 21143 14025
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 24026 14056 24032 14068
rect 23492 14028 24032 14056
rect 14274 13988 14280 14000
rect 13188 13960 13676 13988
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 12621 13923 12679 13929
rect 12621 13889 12633 13923
rect 12667 13889 12679 13923
rect 13188 13920 13216 13960
rect 12621 13883 12679 13889
rect 13004 13892 13216 13920
rect 13265 13923 13323 13929
rect 11882 13852 11888 13864
rect 11808 13824 11888 13852
rect 11808 13793 11836 13824
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 13004 13852 13032 13892
rect 13265 13889 13277 13923
rect 13311 13920 13323 13923
rect 13311 13892 13584 13920
rect 13311 13889 13323 13892
rect 13265 13883 13323 13889
rect 13446 13852 13452 13864
rect 12452 13824 13032 13852
rect 13096 13824 13452 13852
rect 12452 13793 12480 13824
rect 13096 13793 13124 13824
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 11793 13787 11851 13793
rect 11793 13753 11805 13787
rect 11839 13753 11851 13787
rect 11793 13747 11851 13753
rect 12437 13787 12495 13793
rect 12437 13753 12449 13787
rect 12483 13753 12495 13787
rect 12437 13747 12495 13753
rect 13081 13787 13139 13793
rect 13081 13753 13093 13787
rect 13127 13753 13139 13787
rect 13556 13784 13584 13892
rect 13648 13852 13676 13960
rect 13740 13960 14280 13988
rect 13740 13929 13768 13960
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 16316 13960 17540 13988
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13725 13883 13783 13889
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 16316 13929 16344 13960
rect 15749 13923 15807 13929
rect 15749 13920 15761 13923
rect 15160 13892 15761 13920
rect 15160 13880 15166 13892
rect 15749 13889 15761 13892
rect 15795 13889 15807 13923
rect 15749 13883 15807 13889
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13889 16359 13923
rect 16301 13883 16359 13889
rect 15470 13852 15476 13864
rect 13648 13824 15476 13852
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 15764 13852 15792 13883
rect 17402 13880 17408 13932
rect 17460 13880 17466 13932
rect 17512 13920 17540 13960
rect 17678 13948 17684 14000
rect 17736 13988 17742 14000
rect 17862 13988 17868 14000
rect 17736 13960 17868 13988
rect 17736 13948 17742 13960
rect 17862 13948 17868 13960
rect 17920 13988 17926 14000
rect 18233 13991 18291 13997
rect 18233 13988 18245 13991
rect 17920 13960 18245 13988
rect 17920 13948 17926 13960
rect 18233 13957 18245 13960
rect 18279 13988 18291 13991
rect 19058 13988 19064 14000
rect 18279 13960 19064 13988
rect 18279 13957 18291 13960
rect 18233 13951 18291 13957
rect 19058 13948 19064 13960
rect 19116 13948 19122 14000
rect 19426 13948 19432 14000
rect 19484 13988 19490 14000
rect 21910 13988 21916 14000
rect 19484 13960 21916 13988
rect 19484 13948 19490 13960
rect 21910 13948 21916 13960
rect 21968 13948 21974 14000
rect 23109 13991 23167 13997
rect 23109 13957 23121 13991
rect 23155 13988 23167 13991
rect 23492 13988 23520 14028
rect 24026 14016 24032 14028
rect 24084 14016 24090 14068
rect 23155 13960 23520 13988
rect 23155 13957 23167 13960
rect 23109 13951 23167 13957
rect 23658 13948 23664 14000
rect 23716 13948 23722 14000
rect 25130 13948 25136 14000
rect 25188 13948 25194 14000
rect 19444 13920 19472 13948
rect 17512 13892 19472 13920
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 20772 13892 21312 13920
rect 20772 13880 20778 13892
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 15764 13824 16681 13852
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 16669 13815 16727 13821
rect 17681 13855 17739 13861
rect 17681 13821 17693 13855
rect 17727 13821 17739 13855
rect 17681 13815 17739 13821
rect 13722 13784 13728 13796
rect 13556 13756 13728 13784
rect 13081 13747 13139 13753
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 17586 13744 17592 13796
rect 17644 13784 17650 13796
rect 17696 13784 17724 13815
rect 20990 13812 20996 13864
rect 21048 13852 21054 13864
rect 21284 13861 21312 13892
rect 22094 13880 22100 13932
rect 22152 13880 22158 13932
rect 22278 13880 22284 13932
rect 22336 13920 22342 13932
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 22336 13892 22845 13920
rect 22336 13880 22342 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 22833 13883 22891 13889
rect 21177 13855 21235 13861
rect 21177 13852 21189 13855
rect 21048 13824 21189 13852
rect 21048 13812 21054 13824
rect 21177 13821 21189 13824
rect 21223 13821 21235 13855
rect 21177 13815 21235 13821
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13852 21327 13855
rect 21450 13852 21456 13864
rect 21315 13824 21456 13852
rect 21315 13821 21327 13824
rect 21269 13815 21327 13821
rect 21450 13812 21456 13824
rect 21508 13812 21514 13864
rect 21818 13812 21824 13864
rect 21876 13852 21882 13864
rect 21876 13824 22324 13852
rect 21876 13812 21882 13824
rect 22296 13793 22324 13824
rect 24486 13812 24492 13864
rect 24544 13852 24550 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 24544 13824 24593 13852
rect 24544 13812 24550 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 25314 13812 25320 13864
rect 25372 13812 25378 13864
rect 17644 13756 17724 13784
rect 22281 13787 22339 13793
rect 17644 13744 17650 13756
rect 22281 13753 22293 13787
rect 22327 13753 22339 13787
rect 22281 13747 22339 13753
rect 13988 13719 14046 13725
rect 13988 13685 14000 13719
rect 14034 13716 14046 13719
rect 16022 13716 16028 13728
rect 14034 13688 16028 13716
rect 14034 13685 14046 13688
rect 13988 13679 14046 13685
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 17310 13676 17316 13728
rect 17368 13716 17374 13728
rect 18506 13716 18512 13728
rect 17368 13688 18512 13716
rect 17368 13676 17374 13688
rect 18506 13676 18512 13688
rect 18564 13676 18570 13728
rect 20714 13676 20720 13728
rect 20772 13676 20778 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 12526 13472 12532 13524
rect 12584 13512 12590 13524
rect 13722 13512 13728 13524
rect 12584 13484 13728 13512
rect 12584 13472 12590 13484
rect 13722 13472 13728 13484
rect 13780 13512 13786 13524
rect 13817 13515 13875 13521
rect 13817 13512 13829 13515
rect 13780 13484 13829 13512
rect 13780 13472 13786 13484
rect 13817 13481 13829 13484
rect 13863 13481 13875 13515
rect 13817 13475 13875 13481
rect 16022 13472 16028 13524
rect 16080 13512 16086 13524
rect 17494 13512 17500 13524
rect 16080 13484 17500 13512
rect 16080 13472 16086 13484
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 18693 13515 18751 13521
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 19702 13512 19708 13524
rect 18739 13484 19708 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 19702 13472 19708 13484
rect 19760 13472 19766 13524
rect 20622 13472 20628 13524
rect 20680 13512 20686 13524
rect 21174 13512 21180 13524
rect 20680 13484 21180 13512
rect 20680 13472 20686 13484
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 21450 13472 21456 13524
rect 21508 13472 21514 13524
rect 21726 13472 21732 13524
rect 21784 13512 21790 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 21784 13484 24593 13512
rect 21784 13472 21790 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 13446 13404 13452 13456
rect 13504 13444 13510 13456
rect 13541 13447 13599 13453
rect 13541 13444 13553 13447
rect 13504 13416 13553 13444
rect 13504 13404 13510 13416
rect 13541 13413 13553 13416
rect 13587 13444 13599 13447
rect 13587 13416 14412 13444
rect 13587 13413 13599 13416
rect 13541 13407 13599 13413
rect 12710 13376 12716 13388
rect 9600 13348 12716 13376
rect 9600 13317 9628 13348
rect 12710 13336 12716 13348
rect 12768 13376 12774 13388
rect 13354 13376 13360 13388
rect 12768 13348 13360 13376
rect 12768 13336 12774 13348
rect 13354 13336 13360 13348
rect 13412 13336 13418 13388
rect 14274 13336 14280 13388
rect 14332 13336 14338 13388
rect 14384 13376 14412 13416
rect 17862 13404 17868 13456
rect 17920 13444 17926 13456
rect 19150 13444 19156 13456
rect 17920 13416 19156 13444
rect 17920 13404 17926 13416
rect 19150 13404 19156 13416
rect 19208 13404 19214 13456
rect 19337 13447 19395 13453
rect 19337 13413 19349 13447
rect 19383 13444 19395 13447
rect 19426 13444 19432 13456
rect 19383 13416 19432 13444
rect 19383 13413 19395 13416
rect 19337 13407 19395 13413
rect 19426 13404 19432 13416
rect 19484 13404 19490 13456
rect 23658 13404 23664 13456
rect 23716 13444 23722 13456
rect 23937 13447 23995 13453
rect 23937 13444 23949 13447
rect 23716 13416 23949 13444
rect 23716 13404 23722 13416
rect 23937 13413 23949 13416
rect 23983 13444 23995 13447
rect 24121 13447 24179 13453
rect 24121 13444 24133 13447
rect 23983 13416 24133 13444
rect 23983 13413 23995 13416
rect 23937 13407 23995 13413
rect 24121 13413 24133 13416
rect 24167 13413 24179 13447
rect 24121 13407 24179 13413
rect 16390 13376 16396 13388
rect 14384 13348 16396 13376
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 18690 13376 18696 13388
rect 16807 13348 18696 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 19705 13379 19763 13385
rect 19705 13345 19717 13379
rect 19751 13376 19763 13379
rect 21910 13376 21916 13388
rect 19751 13348 21916 13376
rect 19751 13345 19763 13348
rect 19705 13339 19763 13345
rect 9585 13311 9643 13317
rect 9585 13277 9597 13311
rect 9631 13277 9643 13311
rect 11793 13311 11851 13317
rect 11793 13308 11805 13311
rect 9585 13271 9643 13277
rect 10888 13280 11805 13308
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10686 13172 10692 13184
rect 10100 13144 10692 13172
rect 10100 13132 10106 13144
rect 10686 13132 10692 13144
rect 10744 13172 10750 13184
rect 10888 13181 10916 13280
rect 11793 13277 11805 13280
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 18874 13268 18880 13320
rect 18932 13268 18938 13320
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19720 13308 19748 13339
rect 21910 13336 21916 13348
rect 21968 13376 21974 13388
rect 22278 13376 22284 13388
rect 21968 13348 22284 13376
rect 21968 13336 21974 13348
rect 22278 13336 22284 13348
rect 22336 13336 22342 13388
rect 22738 13336 22744 13388
rect 22796 13376 22802 13388
rect 22922 13376 22928 13388
rect 22796 13348 22928 13376
rect 22796 13336 22802 13348
rect 22922 13336 22928 13348
rect 22980 13336 22986 13388
rect 23750 13336 23756 13388
rect 23808 13376 23814 13388
rect 25133 13379 25191 13385
rect 25133 13376 25145 13379
rect 23808 13348 25145 13376
rect 23808 13336 23814 13348
rect 25133 13345 25145 13348
rect 25179 13345 25191 13379
rect 25133 13339 25191 13345
rect 25222 13336 25228 13388
rect 25280 13336 25286 13388
rect 19484 13280 19748 13308
rect 25041 13311 25099 13317
rect 19484 13268 19490 13280
rect 25041 13277 25053 13311
rect 25087 13308 25099 13311
rect 25240 13308 25268 13336
rect 25087 13280 25268 13308
rect 25087 13277 25099 13280
rect 25041 13271 25099 13277
rect 12066 13200 12072 13252
rect 12124 13200 12130 13252
rect 12526 13200 12532 13252
rect 12584 13200 12590 13252
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14550 13240 14556 13252
rect 14240 13212 14556 13240
rect 14240 13200 14246 13212
rect 14550 13200 14556 13212
rect 14608 13200 14614 13252
rect 15010 13240 15016 13252
rect 14936 13212 15016 13240
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10744 13144 10885 13172
rect 10744 13132 10750 13144
rect 10873 13141 10885 13144
rect 10919 13141 10931 13175
rect 10873 13135 10931 13141
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 14936 13172 14964 13212
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 17218 13200 17224 13252
rect 17276 13200 17282 13252
rect 19981 13243 20039 13249
rect 19981 13209 19993 13243
rect 20027 13209 20039 13243
rect 19981 13203 20039 13209
rect 13780 13144 14964 13172
rect 13780 13132 13786 13144
rect 16114 13132 16120 13184
rect 16172 13172 16178 13184
rect 17586 13172 17592 13184
rect 16172 13144 17592 13172
rect 16172 13132 16178 13144
rect 17586 13132 17592 13144
rect 17644 13172 17650 13184
rect 18233 13175 18291 13181
rect 18233 13172 18245 13175
rect 17644 13144 18245 13172
rect 17644 13132 17650 13144
rect 18233 13141 18245 13144
rect 18279 13141 18291 13175
rect 18233 13135 18291 13141
rect 19058 13132 19064 13184
rect 19116 13172 19122 13184
rect 19518 13172 19524 13184
rect 19116 13144 19524 13172
rect 19116 13132 19122 13144
rect 19518 13132 19524 13144
rect 19576 13132 19582 13184
rect 19996 13172 20024 13203
rect 20622 13200 20628 13252
rect 20680 13200 20686 13252
rect 22189 13243 22247 13249
rect 22189 13209 22201 13243
rect 22235 13240 22247 13243
rect 22462 13240 22468 13252
rect 22235 13212 22468 13240
rect 22235 13209 22247 13212
rect 22189 13203 22247 13209
rect 22462 13200 22468 13212
rect 22520 13200 22526 13252
rect 22738 13200 22744 13252
rect 22796 13200 22802 13252
rect 24949 13243 25007 13249
rect 24949 13209 24961 13243
rect 24995 13240 25007 13243
rect 25222 13240 25228 13252
rect 24995 13212 25228 13240
rect 24995 13209 25007 13212
rect 24949 13203 25007 13209
rect 25222 13200 25228 13212
rect 25280 13200 25286 13252
rect 20806 13172 20812 13184
rect 19996 13144 20812 13172
rect 20806 13132 20812 13144
rect 20864 13172 20870 13184
rect 23661 13175 23719 13181
rect 23661 13172 23673 13175
rect 20864 13144 23673 13172
rect 20864 13132 20870 13144
rect 23661 13141 23673 13144
rect 23707 13141 23719 13175
rect 23661 13135 23719 13141
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 12526 12928 12532 12980
rect 12584 12928 12590 12980
rect 14274 12928 14280 12980
rect 14332 12928 14338 12980
rect 15427 12971 15485 12977
rect 15427 12937 15439 12971
rect 15473 12968 15485 12971
rect 22094 12968 22100 12980
rect 15473 12940 22100 12968
rect 15473 12937 15485 12940
rect 15427 12931 15485 12937
rect 22094 12928 22100 12940
rect 22152 12928 22158 12980
rect 22462 12928 22468 12980
rect 22520 12968 22526 12980
rect 23750 12968 23756 12980
rect 22520 12940 23756 12968
rect 22520 12928 22526 12940
rect 23750 12928 23756 12940
rect 23808 12928 23814 12980
rect 24854 12928 24860 12980
rect 24912 12928 24918 12980
rect 12710 12860 12716 12912
rect 12768 12900 12774 12912
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 12768 12872 13001 12900
rect 12768 12860 12774 12872
rect 12989 12869 13001 12872
rect 13035 12869 13047 12903
rect 12989 12863 13047 12869
rect 15010 12860 15016 12912
rect 15068 12900 15074 12912
rect 16298 12900 16304 12912
rect 15068 12872 16304 12900
rect 15068 12860 15074 12872
rect 16298 12860 16304 12872
rect 16356 12900 16362 12912
rect 17218 12900 17224 12912
rect 16356 12872 17224 12900
rect 16356 12860 16362 12872
rect 17218 12860 17224 12872
rect 17276 12900 17282 12912
rect 17586 12900 17592 12912
rect 17276 12872 17592 12900
rect 17276 12860 17282 12872
rect 17586 12860 17592 12872
rect 17644 12860 17650 12912
rect 18874 12860 18880 12912
rect 18932 12900 18938 12912
rect 21542 12900 21548 12912
rect 18932 12872 21548 12900
rect 18932 12860 18938 12872
rect 21542 12860 21548 12872
rect 21600 12860 21606 12912
rect 22278 12900 22284 12912
rect 21836 12872 22284 12900
rect 15197 12835 15255 12841
rect 15197 12801 15209 12835
rect 15243 12832 15255 12835
rect 16574 12832 16580 12844
rect 15243 12804 16580 12832
rect 15243 12801 15255 12804
rect 15197 12795 15255 12801
rect 16574 12792 16580 12804
rect 16632 12792 16638 12844
rect 18414 12792 18420 12844
rect 18472 12832 18478 12844
rect 19429 12835 19487 12841
rect 19429 12832 19441 12835
rect 18472 12804 19441 12832
rect 18472 12792 18478 12804
rect 19429 12801 19441 12804
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 20625 12835 20683 12841
rect 20625 12801 20637 12835
rect 20671 12832 20683 12835
rect 21634 12832 21640 12844
rect 20671 12804 21640 12832
rect 20671 12801 20683 12804
rect 20625 12795 20683 12801
rect 21634 12792 21640 12804
rect 21692 12792 21698 12844
rect 13354 12724 13360 12776
rect 13412 12764 13418 12776
rect 14274 12764 14280 12776
rect 13412 12736 14280 12764
rect 13412 12724 13418 12736
rect 14274 12724 14280 12736
rect 14332 12764 14338 12776
rect 15470 12764 15476 12776
rect 14332 12736 15476 12764
rect 14332 12724 14338 12736
rect 15470 12724 15476 12736
rect 15528 12764 15534 12776
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 15528 12736 16865 12764
rect 15528 12724 15534 12736
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12764 17187 12767
rect 17494 12764 17500 12776
rect 17175 12736 17500 12764
rect 17175 12733 17187 12736
rect 17129 12727 17187 12733
rect 17494 12724 17500 12736
rect 17552 12764 17558 12776
rect 18322 12764 18328 12776
rect 17552 12736 18328 12764
rect 17552 12724 17558 12736
rect 18322 12724 18328 12736
rect 18380 12724 18386 12776
rect 18690 12724 18696 12776
rect 18748 12764 18754 12776
rect 19150 12764 19156 12776
rect 18748 12736 19156 12764
rect 18748 12724 18754 12736
rect 19150 12724 19156 12736
rect 19208 12724 19214 12776
rect 19518 12724 19524 12776
rect 19576 12724 19582 12776
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 18598 12656 18604 12708
rect 18656 12696 18662 12708
rect 19628 12696 19656 12727
rect 19794 12724 19800 12776
rect 19852 12764 19858 12776
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 19852 12736 20729 12764
rect 19852 12724 19858 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 20809 12767 20867 12773
rect 20809 12733 20821 12767
rect 20855 12733 20867 12767
rect 20809 12727 20867 12733
rect 18656 12668 19656 12696
rect 19707 12668 20392 12696
rect 18656 12656 18662 12668
rect 19058 12588 19064 12640
rect 19116 12588 19122 12640
rect 19150 12588 19156 12640
rect 19208 12628 19214 12640
rect 19707 12628 19735 12668
rect 19208 12600 19735 12628
rect 19208 12588 19214 12600
rect 20254 12588 20260 12640
rect 20312 12588 20318 12640
rect 20364 12628 20392 12668
rect 20622 12656 20628 12708
rect 20680 12696 20686 12708
rect 20824 12696 20852 12727
rect 21174 12724 21180 12776
rect 21232 12764 21238 12776
rect 21269 12767 21327 12773
rect 21269 12764 21281 12767
rect 21232 12736 21281 12764
rect 21232 12724 21238 12736
rect 21269 12733 21281 12736
rect 21315 12764 21327 12767
rect 21836 12764 21864 12872
rect 22278 12860 22284 12872
rect 22336 12900 22342 12912
rect 22336 12872 22770 12900
rect 22336 12860 22342 12872
rect 21910 12792 21916 12844
rect 21968 12832 21974 12844
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21968 12804 22017 12832
rect 21968 12792 21974 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 24397 12835 24455 12841
rect 24397 12801 24409 12835
rect 24443 12832 24455 12835
rect 24762 12832 24768 12844
rect 24443 12804 24768 12832
rect 24443 12801 24455 12804
rect 24397 12795 24455 12801
rect 24762 12792 24768 12804
rect 24820 12792 24826 12844
rect 21315 12736 21864 12764
rect 21315 12733 21327 12736
rect 21269 12727 21327 12733
rect 22278 12724 22284 12776
rect 22336 12764 22342 12776
rect 22738 12764 22744 12776
rect 22336 12736 22744 12764
rect 22336 12724 22342 12736
rect 22738 12724 22744 12736
rect 22796 12724 22802 12776
rect 20680 12668 20852 12696
rect 20916 12668 22094 12696
rect 20680 12656 20686 12668
rect 20916 12628 20944 12668
rect 20364 12600 20944 12628
rect 22066 12628 22094 12668
rect 24210 12656 24216 12708
rect 24268 12656 24274 12708
rect 23382 12628 23388 12640
rect 22066 12600 23388 12628
rect 23382 12588 23388 12600
rect 23440 12588 23446 12640
rect 25130 12588 25136 12640
rect 25188 12628 25194 12640
rect 25317 12631 25375 12637
rect 25317 12628 25329 12631
rect 25188 12600 25329 12628
rect 25188 12588 25194 12600
rect 25317 12597 25329 12600
rect 25363 12597 25375 12631
rect 25317 12591 25375 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 13722 12384 13728 12436
rect 13780 12384 13786 12436
rect 13906 12384 13912 12436
rect 13964 12384 13970 12436
rect 15010 12384 15016 12436
rect 15068 12424 15074 12436
rect 15381 12427 15439 12433
rect 15381 12424 15393 12427
rect 15068 12396 15393 12424
rect 15068 12384 15074 12396
rect 15381 12393 15393 12396
rect 15427 12393 15439 12427
rect 15381 12387 15439 12393
rect 16390 12384 16396 12436
rect 16448 12424 16454 12436
rect 16448 12396 17080 12424
rect 16448 12384 16454 12396
rect 17052 12356 17080 12396
rect 17494 12384 17500 12436
rect 17552 12384 17558 12436
rect 18782 12384 18788 12436
rect 18840 12384 18846 12436
rect 19886 12384 19892 12436
rect 19944 12424 19950 12436
rect 22002 12424 22008 12436
rect 19944 12396 22008 12424
rect 19944 12384 19950 12396
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 22278 12384 22284 12436
rect 22336 12424 22342 12436
rect 24029 12427 24087 12433
rect 24029 12424 24041 12427
rect 22336 12396 24041 12424
rect 22336 12384 22342 12396
rect 24029 12393 24041 12396
rect 24075 12393 24087 12427
rect 24029 12387 24087 12393
rect 24854 12384 24860 12436
rect 24912 12424 24918 12436
rect 25317 12427 25375 12433
rect 25317 12424 25329 12427
rect 24912 12396 25329 12424
rect 24912 12384 24918 12396
rect 25317 12393 25329 12396
rect 25363 12393 25375 12427
rect 25317 12387 25375 12393
rect 18800 12356 18828 12384
rect 17052 12328 18828 12356
rect 4982 12248 4988 12300
rect 5040 12288 5046 12300
rect 14277 12291 14335 12297
rect 14277 12288 14289 12291
rect 5040 12260 14289 12288
rect 5040 12248 5046 12260
rect 14277 12257 14289 12260
rect 14323 12257 14335 12291
rect 14277 12251 14335 12257
rect 15470 12248 15476 12300
rect 15528 12288 15534 12300
rect 15749 12291 15807 12297
rect 15749 12288 15761 12291
rect 15528 12260 15761 12288
rect 15528 12248 15534 12260
rect 15749 12257 15761 12260
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 17402 12248 17408 12300
rect 17460 12288 17466 12300
rect 17957 12291 18015 12297
rect 17957 12288 17969 12291
rect 17460 12260 17969 12288
rect 17460 12248 17466 12260
rect 17957 12257 17969 12260
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 18874 12248 18880 12300
rect 18932 12248 18938 12300
rect 19702 12248 19708 12300
rect 19760 12288 19766 12300
rect 20346 12288 20352 12300
rect 19760 12260 20352 12288
rect 19760 12248 19766 12260
rect 20346 12248 20352 12260
rect 20404 12248 20410 12300
rect 21358 12248 21364 12300
rect 21416 12288 21422 12300
rect 21910 12288 21916 12300
rect 21416 12260 21916 12288
rect 21416 12248 21422 12260
rect 21910 12248 21916 12260
rect 21968 12288 21974 12300
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 21968 12260 22293 12288
rect 21968 12248 21974 12260
rect 22281 12257 22293 12260
rect 22327 12257 22339 12291
rect 22281 12251 22339 12257
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12288 22615 12291
rect 24486 12288 24492 12300
rect 22603 12260 24492 12288
rect 22603 12257 22615 12260
rect 22557 12251 22615 12257
rect 24486 12248 24492 12260
rect 24544 12248 24550 12300
rect 24578 12248 24584 12300
rect 24636 12248 24642 12300
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12220 14611 12223
rect 15562 12220 15568 12232
rect 14599 12192 15568 12220
rect 14599 12189 14611 12192
rect 14553 12183 14611 12189
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 19334 12180 19340 12232
rect 19392 12220 19398 12232
rect 19429 12223 19487 12229
rect 19429 12220 19441 12223
rect 19392 12192 19441 12220
rect 19392 12180 19398 12192
rect 19429 12189 19441 12192
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 21634 12180 21640 12232
rect 21692 12180 21698 12232
rect 16025 12155 16083 12161
rect 16025 12121 16037 12155
rect 16071 12152 16083 12155
rect 16114 12152 16120 12164
rect 16071 12124 16120 12152
rect 16071 12121 16083 12124
rect 16025 12115 16083 12121
rect 16114 12112 16120 12124
rect 16172 12112 16178 12164
rect 16298 12112 16304 12164
rect 16356 12152 16362 12164
rect 16356 12124 16514 12152
rect 16356 12112 16362 12124
rect 18690 12112 18696 12164
rect 18748 12112 18754 12164
rect 19242 12152 19248 12164
rect 18800 12124 19248 12152
rect 17586 12044 17592 12096
rect 17644 12084 17650 12096
rect 18800 12084 18828 12124
rect 19242 12112 19248 12124
rect 19300 12152 19306 12164
rect 19300 12124 20194 12152
rect 19300 12112 19306 12124
rect 21542 12112 21548 12164
rect 21600 12152 21606 12164
rect 21600 12124 23046 12152
rect 21600 12112 21606 12124
rect 17644 12056 18828 12084
rect 17644 12044 17650 12056
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 19518 12084 19524 12096
rect 18932 12056 19524 12084
rect 18932 12044 18938 12056
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 19794 12044 19800 12096
rect 19852 12084 19858 12096
rect 20622 12084 20628 12096
rect 19852 12056 20628 12084
rect 19852 12044 19858 12056
rect 20622 12044 20628 12056
rect 20680 12084 20686 12096
rect 21177 12087 21235 12093
rect 21177 12084 21189 12087
rect 20680 12056 21189 12084
rect 20680 12044 20686 12056
rect 21177 12053 21189 12056
rect 21223 12053 21235 12087
rect 22940 12084 22968 12124
rect 25041 12087 25099 12093
rect 25041 12084 25053 12087
rect 22940 12056 25053 12084
rect 21177 12047 21235 12053
rect 25041 12053 25053 12056
rect 25087 12084 25099 12087
rect 25130 12084 25136 12096
rect 25087 12056 25136 12084
rect 25087 12053 25099 12056
rect 25041 12047 25099 12053
rect 25130 12044 25136 12056
rect 25188 12044 25194 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 14550 11840 14556 11892
rect 14608 11840 14614 11892
rect 15102 11840 15108 11892
rect 15160 11840 15166 11892
rect 15654 11840 15660 11892
rect 15712 11840 15718 11892
rect 19334 11880 19340 11892
rect 17144 11852 19340 11880
rect 13354 11812 13360 11824
rect 12820 11784 13360 11812
rect 12820 11753 12848 11784
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 13722 11772 13728 11824
rect 13780 11772 13786 11824
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 15289 11747 15347 11753
rect 15289 11713 15301 11747
rect 15335 11744 15347 11747
rect 15672 11744 15700 11840
rect 17144 11753 17172 11852
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 21266 11880 21272 11892
rect 19444 11852 21272 11880
rect 17494 11772 17500 11824
rect 17552 11812 17558 11824
rect 17552 11784 17894 11812
rect 17552 11772 17558 11784
rect 18874 11772 18880 11824
rect 18932 11812 18938 11824
rect 19444 11812 19472 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 25498 11880 25504 11892
rect 22066 11852 25504 11880
rect 18932 11784 19472 11812
rect 19705 11815 19763 11821
rect 18932 11772 18938 11784
rect 19705 11781 19717 11815
rect 19751 11812 19763 11815
rect 19794 11812 19800 11824
rect 19751 11784 19800 11812
rect 19751 11781 19763 11784
rect 19705 11775 19763 11781
rect 19794 11772 19800 11784
rect 19852 11772 19858 11824
rect 20990 11772 20996 11824
rect 21048 11812 21054 11824
rect 22066 11812 22094 11852
rect 25498 11840 25504 11852
rect 25556 11840 25562 11892
rect 21048 11784 22094 11812
rect 23293 11815 23351 11821
rect 21048 11772 21054 11784
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 15335 11716 15700 11744
rect 16301 11747 16359 11753
rect 15335 11713 15347 11716
rect 15289 11707 15347 11713
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 17129 11747 17187 11753
rect 16347 11716 16804 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11676 13139 11679
rect 13446 11676 13452 11688
rect 13127 11648 13452 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 14090 11568 14096 11620
rect 14148 11608 14154 11620
rect 16117 11611 16175 11617
rect 16117 11608 16129 11611
rect 14148 11580 16129 11608
rect 14148 11568 14154 11580
rect 16117 11577 16129 11580
rect 16163 11577 16175 11611
rect 16117 11571 16175 11577
rect 16776 11549 16804 11716
rect 17129 11713 17141 11747
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 19426 11704 19432 11756
rect 19484 11704 19490 11756
rect 21174 11744 21180 11756
rect 20838 11716 21180 11744
rect 21174 11704 21180 11716
rect 21232 11744 21238 11756
rect 21453 11747 21511 11753
rect 21453 11744 21465 11747
rect 21232 11716 21465 11744
rect 21232 11704 21238 11716
rect 21453 11713 21465 11716
rect 21499 11744 21511 11747
rect 21542 11744 21548 11756
rect 21499 11716 21548 11744
rect 21499 11713 21511 11716
rect 21453 11707 21511 11713
rect 21542 11704 21548 11716
rect 21600 11704 21606 11756
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11676 17463 11679
rect 18598 11676 18604 11688
rect 17451 11648 18604 11676
rect 17451 11645 17463 11648
rect 17405 11639 17463 11645
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 19334 11636 19340 11688
rect 19392 11676 19398 11688
rect 19392 11648 21772 11676
rect 19392 11636 19398 11648
rect 21082 11568 21088 11620
rect 21140 11608 21146 11620
rect 21177 11611 21235 11617
rect 21177 11608 21189 11611
rect 21140 11580 21189 11608
rect 21140 11568 21146 11580
rect 21177 11577 21189 11580
rect 21223 11608 21235 11611
rect 21634 11608 21640 11620
rect 21223 11580 21640 11608
rect 21223 11577 21235 11580
rect 21177 11571 21235 11577
rect 21634 11568 21640 11580
rect 21692 11568 21698 11620
rect 16761 11543 16819 11549
rect 16761 11509 16773 11543
rect 16807 11540 16819 11543
rect 18782 11540 18788 11552
rect 16807 11512 18788 11540
rect 16807 11509 16819 11512
rect 16761 11503 16819 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 18877 11543 18935 11549
rect 18877 11509 18889 11543
rect 18923 11540 18935 11543
rect 19702 11540 19708 11552
rect 18923 11512 19708 11540
rect 18923 11509 18935 11512
rect 18877 11503 18935 11509
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 19794 11500 19800 11552
rect 19852 11540 19858 11552
rect 20990 11540 20996 11552
rect 19852 11512 20996 11540
rect 19852 11500 19858 11512
rect 20990 11500 20996 11512
rect 21048 11500 21054 11552
rect 21744 11540 21772 11648
rect 22002 11636 22008 11688
rect 22060 11676 22066 11688
rect 22112 11676 22140 11707
rect 23934 11704 23940 11756
rect 23992 11704 23998 11756
rect 22060 11648 22140 11676
rect 22060 11636 22066 11648
rect 24762 11636 24768 11688
rect 24820 11636 24826 11688
rect 26050 11540 26056 11552
rect 21744 11512 26056 11540
rect 26050 11500 26056 11512
rect 26108 11500 26114 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 14737 11339 14795 11345
rect 14737 11305 14749 11339
rect 14783 11336 14795 11339
rect 15010 11336 15016 11348
rect 14783 11308 15016 11336
rect 14783 11305 14795 11308
rect 14737 11299 14795 11305
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 16761 11339 16819 11345
rect 15519 11308 16712 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 16114 11228 16120 11280
rect 16172 11228 16178 11280
rect 16684 11268 16712 11308
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16942 11336 16948 11348
rect 16807 11308 16948 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16942 11296 16948 11308
rect 17000 11296 17006 11348
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 17368 11308 17417 11336
rect 17368 11296 17374 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17405 11299 17463 11305
rect 18690 11296 18696 11348
rect 18748 11296 18754 11348
rect 19794 11336 19800 11348
rect 18800 11308 19800 11336
rect 18800 11268 18828 11308
rect 19794 11296 19800 11308
rect 19852 11296 19858 11348
rect 20806 11296 20812 11348
rect 20864 11336 20870 11348
rect 22005 11339 22063 11345
rect 22005 11336 22017 11339
rect 20864 11308 22017 11336
rect 20864 11296 20870 11308
rect 22005 11305 22017 11308
rect 22051 11305 22063 11339
rect 22005 11299 22063 11305
rect 16684 11240 18828 11268
rect 19242 11228 19248 11280
rect 19300 11268 19306 11280
rect 19337 11271 19395 11277
rect 19337 11268 19349 11271
rect 19300 11240 19349 11268
rect 19300 11228 19306 11240
rect 19337 11237 19349 11240
rect 19383 11268 19395 11271
rect 19429 11271 19487 11277
rect 19429 11268 19441 11271
rect 19383 11240 19441 11268
rect 19383 11237 19395 11240
rect 19337 11231 19395 11237
rect 19429 11237 19441 11240
rect 19475 11237 19487 11271
rect 19429 11231 19487 11237
rect 19610 11228 19616 11280
rect 19668 11268 19674 11280
rect 20901 11271 20959 11277
rect 20901 11268 20913 11271
rect 19668 11240 20913 11268
rect 19668 11228 19674 11240
rect 20901 11237 20913 11240
rect 20947 11268 20959 11271
rect 20990 11268 20996 11280
rect 20947 11240 20996 11268
rect 20947 11237 20959 11240
rect 20901 11231 20959 11237
rect 20990 11228 20996 11240
rect 21048 11228 21054 11280
rect 21177 11271 21235 11277
rect 21177 11237 21189 11271
rect 21223 11268 21235 11271
rect 25038 11268 25044 11280
rect 21223 11240 25044 11268
rect 21223 11237 21235 11240
rect 21177 11231 21235 11237
rect 25038 11228 25044 11240
rect 25096 11228 25102 11280
rect 17862 11200 17868 11212
rect 16960 11172 17868 11200
rect 16960 11144 16988 11172
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11200 18107 11203
rect 18414 11200 18420 11212
rect 18095 11172 18420 11200
rect 18095 11169 18107 11172
rect 18049 11163 18107 11169
rect 18414 11160 18420 11172
rect 18472 11160 18478 11212
rect 21726 11200 21732 11212
rect 19444 11172 21732 11200
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11132 15715 11135
rect 15746 11132 15752 11144
rect 15703 11104 15752 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11132 16359 11135
rect 16390 11132 16396 11144
rect 16347 11104 16396 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 16942 11092 16948 11144
rect 17000 11092 17006 11144
rect 17589 11135 17647 11141
rect 17589 11101 17601 11135
rect 17635 11101 17647 11135
rect 17589 11095 17647 11101
rect 18877 11135 18935 11141
rect 18877 11101 18889 11135
rect 18923 11132 18935 11135
rect 19444 11132 19472 11172
rect 21726 11160 21732 11172
rect 21784 11160 21790 11212
rect 23845 11203 23903 11209
rect 23845 11169 23857 11203
rect 23891 11200 23903 11203
rect 24854 11200 24860 11212
rect 23891 11172 24860 11200
rect 23891 11169 23903 11172
rect 23845 11163 23903 11169
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 20438 11132 20444 11144
rect 18923 11104 19472 11132
rect 19536 11104 20444 11132
rect 18923 11101 18935 11104
rect 18877 11095 18935 11101
rect 17604 11064 17632 11095
rect 19536 11064 19564 11104
rect 20438 11092 20444 11104
rect 20496 11092 20502 11144
rect 20898 11092 20904 11144
rect 20956 11132 20962 11144
rect 21361 11135 21419 11141
rect 21361 11132 21373 11135
rect 20956 11104 21373 11132
rect 20956 11092 20962 11104
rect 21361 11101 21373 11104
rect 21407 11101 21419 11135
rect 21361 11095 21419 11101
rect 21542 11092 21548 11144
rect 21600 11132 21606 11144
rect 21637 11135 21695 11141
rect 21637 11132 21649 11135
rect 21600 11104 21649 11132
rect 21600 11092 21606 11104
rect 21637 11101 21649 11104
rect 21683 11101 21695 11135
rect 21637 11095 21695 11101
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11132 22247 11135
rect 22370 11132 22376 11144
rect 22235 11104 22376 11132
rect 22235 11101 22247 11104
rect 22189 11095 22247 11101
rect 22370 11092 22376 11104
rect 22428 11092 22434 11144
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 24394 11092 24400 11144
rect 24452 11132 24458 11144
rect 24765 11135 24823 11141
rect 24765 11132 24777 11135
rect 24452 11104 24777 11132
rect 24452 11092 24458 11104
rect 24765 11101 24777 11104
rect 24811 11101 24823 11135
rect 24765 11095 24823 11101
rect 17604 11036 19564 11064
rect 19702 11024 19708 11076
rect 19760 11064 19766 11076
rect 19981 11067 20039 11073
rect 19981 11064 19993 11067
rect 19760 11036 19993 11064
rect 19760 11024 19766 11036
rect 19981 11033 19993 11036
rect 20027 11033 20039 11067
rect 19981 11027 20039 11033
rect 20165 11067 20223 11073
rect 20165 11033 20177 11067
rect 20211 11064 20223 11067
rect 20530 11064 20536 11076
rect 20211 11036 20536 11064
rect 20211 11033 20223 11036
rect 20165 11027 20223 11033
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 20717 11067 20775 11073
rect 20717 11033 20729 11067
rect 20763 11064 20775 11067
rect 21266 11064 21272 11076
rect 20763 11036 21272 11064
rect 20763 11033 20775 11036
rect 20717 11027 20775 11033
rect 21266 11024 21272 11036
rect 21324 11024 21330 11076
rect 21726 11024 21732 11076
rect 21784 11064 21790 11076
rect 22830 11064 22836 11076
rect 21784 11036 22836 11064
rect 21784 11024 21790 11036
rect 22830 11024 22836 11036
rect 22888 11024 22894 11076
rect 15562 10956 15568 11008
rect 15620 10996 15626 11008
rect 21910 10996 21916 11008
rect 15620 10968 21916 10996
rect 15620 10956 15626 10968
rect 21910 10956 21916 10968
rect 21968 10956 21974 11008
rect 24578 10956 24584 11008
rect 24636 10956 24642 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 15746 10752 15752 10804
rect 15804 10752 15810 10804
rect 16390 10752 16396 10804
rect 16448 10752 16454 10804
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 17037 10795 17095 10801
rect 17037 10792 17049 10795
rect 17000 10764 17049 10792
rect 17000 10752 17006 10764
rect 17037 10761 17049 10764
rect 17083 10761 17095 10795
rect 17037 10755 17095 10761
rect 17678 10752 17684 10804
rect 17736 10792 17742 10804
rect 18693 10795 18751 10801
rect 18693 10792 18705 10795
rect 17736 10764 18705 10792
rect 17736 10752 17742 10764
rect 18693 10761 18705 10764
rect 18739 10761 18751 10795
rect 22554 10792 22560 10804
rect 18693 10755 18751 10761
rect 21744 10764 22560 10792
rect 17405 10727 17463 10733
rect 17405 10693 17417 10727
rect 17451 10724 17463 10727
rect 19334 10724 19340 10736
rect 17451 10696 19340 10724
rect 17451 10693 17463 10696
rect 17405 10687 17463 10693
rect 19334 10684 19340 10696
rect 19392 10684 19398 10736
rect 21082 10724 21088 10736
rect 20088 10696 21088 10724
rect 18233 10659 18291 10665
rect 18233 10625 18245 10659
rect 18279 10656 18291 10659
rect 18322 10656 18328 10668
rect 18279 10628 18328 10656
rect 18279 10625 18291 10628
rect 18233 10619 18291 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 18874 10616 18880 10668
rect 18932 10616 18938 10668
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10656 19579 10659
rect 19978 10656 19984 10668
rect 19567 10628 19984 10656
rect 19567 10625 19579 10628
rect 19521 10619 19579 10625
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 17034 10548 17040 10600
rect 17092 10548 17098 10600
rect 20088 10588 20116 10696
rect 21082 10684 21088 10696
rect 21140 10684 21146 10736
rect 20165 10659 20223 10665
rect 20165 10625 20177 10659
rect 20211 10625 20223 10659
rect 20165 10619 20223 10625
rect 19352 10560 20116 10588
rect 20180 10588 20208 10619
rect 20714 10616 20720 10668
rect 20772 10656 20778 10668
rect 20809 10659 20867 10665
rect 20809 10656 20821 10659
rect 20772 10628 20821 10656
rect 20772 10616 20778 10628
rect 20809 10625 20821 10628
rect 20855 10625 20867 10659
rect 20809 10619 20867 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10656 21511 10659
rect 21744 10656 21772 10764
rect 22554 10752 22560 10764
rect 22612 10752 22618 10804
rect 21910 10684 21916 10736
rect 21968 10724 21974 10736
rect 23293 10727 23351 10733
rect 21968 10696 23060 10724
rect 21968 10684 21974 10696
rect 21499 10628 21772 10656
rect 21499 10625 21511 10628
rect 21453 10619 21511 10625
rect 22094 10616 22100 10668
rect 22152 10616 22158 10668
rect 23032 10656 23060 10696
rect 23293 10693 23305 10727
rect 23339 10724 23351 10727
rect 24854 10724 24860 10736
rect 23339 10696 24860 10724
rect 23339 10693 23351 10696
rect 23293 10687 23351 10693
rect 24854 10684 24860 10696
rect 24912 10684 24918 10736
rect 23937 10659 23995 10665
rect 23937 10656 23949 10659
rect 23032 10628 23949 10656
rect 23937 10625 23949 10628
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 24578 10588 24584 10600
rect 20180 10560 24584 10588
rect 17052 10520 17080 10548
rect 19352 10529 19380 10560
rect 24578 10548 24584 10560
rect 24636 10548 24642 10600
rect 24670 10548 24676 10600
rect 24728 10548 24734 10600
rect 18049 10523 18107 10529
rect 18049 10520 18061 10523
rect 17052 10492 18061 10520
rect 18049 10489 18061 10492
rect 18095 10489 18107 10523
rect 18049 10483 18107 10489
rect 19337 10523 19395 10529
rect 19337 10489 19349 10523
rect 19383 10489 19395 10523
rect 19337 10483 19395 10489
rect 19981 10523 20039 10529
rect 19981 10489 19993 10523
rect 20027 10520 20039 10523
rect 22462 10520 22468 10532
rect 20027 10492 22468 10520
rect 20027 10489 20039 10492
rect 19981 10483 20039 10489
rect 22462 10480 22468 10492
rect 22520 10480 22526 10532
rect 20625 10455 20683 10461
rect 20625 10421 20637 10455
rect 20671 10452 20683 10455
rect 21174 10452 21180 10464
rect 20671 10424 21180 10452
rect 20671 10421 20683 10424
rect 20625 10415 20683 10421
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 21266 10412 21272 10464
rect 21324 10412 21330 10464
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 17773 10251 17831 10257
rect 17773 10217 17785 10251
rect 17819 10248 17831 10251
rect 18322 10248 18328 10260
rect 17819 10220 18328 10248
rect 17819 10217 17831 10220
rect 17773 10211 17831 10217
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 19426 10208 19432 10260
rect 19484 10208 19490 10260
rect 20714 10208 20720 10260
rect 20772 10208 20778 10260
rect 21634 10257 21640 10260
rect 21624 10251 21640 10257
rect 21624 10217 21636 10251
rect 21624 10211 21640 10217
rect 21634 10208 21640 10211
rect 21692 10208 21698 10260
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 24581 10251 24639 10257
rect 24581 10248 24593 10251
rect 21876 10220 24593 10248
rect 21876 10208 21882 10220
rect 24581 10217 24593 10220
rect 24627 10217 24639 10251
rect 24581 10211 24639 10217
rect 16574 10140 16580 10192
rect 16632 10180 16638 10192
rect 16632 10152 21496 10180
rect 16632 10140 16638 10152
rect 18049 10115 18107 10121
rect 18049 10081 18061 10115
rect 18095 10112 18107 10115
rect 21266 10112 21272 10124
rect 18095 10084 21272 10112
rect 18095 10081 18107 10084
rect 18049 10075 18107 10081
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 21358 10072 21364 10124
rect 21416 10072 21422 10124
rect 21468 10112 21496 10152
rect 22830 10140 22836 10192
rect 22888 10180 22894 10192
rect 23109 10183 23167 10189
rect 23109 10180 23121 10183
rect 22888 10152 23121 10180
rect 22888 10140 22894 10152
rect 23109 10149 23121 10152
rect 23155 10180 23167 10183
rect 23155 10152 25176 10180
rect 23155 10149 23167 10152
rect 23109 10143 23167 10149
rect 23842 10112 23848 10124
rect 21468 10084 23848 10112
rect 23842 10072 23848 10084
rect 23900 10072 23906 10124
rect 25148 10121 25176 10152
rect 25133 10115 25191 10121
rect 25133 10081 25145 10115
rect 25179 10081 25191 10115
rect 25133 10075 25191 10081
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 18340 9976 18368 10007
rect 19610 10004 19616 10056
rect 19668 10004 19674 10056
rect 20714 10044 20720 10056
rect 19996 10016 20720 10044
rect 19996 9976 20024 10016
rect 20714 10004 20720 10016
rect 20772 10004 20778 10056
rect 20901 10047 20959 10053
rect 20901 10013 20913 10047
rect 20947 10044 20959 10047
rect 20947 10016 21404 10044
rect 20947 10013 20959 10016
rect 20901 10007 20959 10013
rect 18340 9948 20024 9976
rect 21376 9976 21404 10016
rect 23566 10004 23572 10056
rect 23624 10044 23630 10056
rect 24029 10047 24087 10053
rect 24029 10044 24041 10047
rect 23624 10016 24041 10044
rect 23624 10004 23630 10016
rect 24029 10013 24041 10016
rect 24075 10013 24087 10047
rect 24029 10007 24087 10013
rect 25041 10047 25099 10053
rect 25041 10013 25053 10047
rect 25087 10044 25099 10047
rect 25406 10044 25412 10056
rect 25087 10016 25412 10044
rect 25087 10013 25099 10016
rect 25041 10007 25099 10013
rect 25406 10004 25412 10016
rect 25464 10004 25470 10056
rect 21726 9976 21732 9988
rect 21376 9948 21732 9976
rect 21726 9936 21732 9948
rect 21784 9936 21790 9988
rect 21910 9936 21916 9988
rect 21968 9976 21974 9988
rect 24949 9979 25007 9985
rect 24949 9976 24961 9979
rect 21968 9948 22126 9976
rect 23216 9948 24961 9976
rect 21968 9936 21974 9948
rect 20073 9911 20131 9917
rect 20073 9877 20085 9911
rect 20119 9908 20131 9911
rect 23216 9908 23244 9948
rect 24949 9945 24961 9948
rect 24995 9945 25007 9979
rect 24949 9939 25007 9945
rect 20119 9880 23244 9908
rect 20119 9877 20131 9880
rect 20073 9871 20131 9877
rect 23842 9868 23848 9920
rect 23900 9868 23906 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 21637 9707 21695 9713
rect 21637 9673 21649 9707
rect 21683 9704 21695 9707
rect 21726 9704 21732 9716
rect 21683 9676 21732 9704
rect 21683 9673 21695 9676
rect 21637 9667 21695 9673
rect 21726 9664 21732 9676
rect 21784 9664 21790 9716
rect 19334 9636 19340 9648
rect 18892 9608 19340 9636
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 18892 9577 18920 9608
rect 19334 9596 19340 9608
rect 19392 9636 19398 9648
rect 20070 9636 20076 9648
rect 19392 9608 20076 9636
rect 19392 9596 19398 9608
rect 20070 9596 20076 9608
rect 20128 9596 20134 9648
rect 20714 9596 20720 9648
rect 20772 9636 20778 9648
rect 20772 9608 22140 9636
rect 20772 9596 20778 9608
rect 18233 9571 18291 9577
rect 18233 9568 18245 9571
rect 8536 9540 18245 9568
rect 8536 9528 8542 9540
rect 18233 9537 18245 9540
rect 18279 9537 18291 9571
rect 18233 9531 18291 9537
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9537 18935 9571
rect 18877 9531 18935 9537
rect 19521 9571 19579 9577
rect 19521 9537 19533 9571
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 20165 9571 20223 9577
rect 20165 9537 20177 9571
rect 20211 9568 20223 9571
rect 20806 9568 20812 9580
rect 20211 9540 20812 9568
rect 20211 9537 20223 9540
rect 20165 9531 20223 9537
rect 17126 9460 17132 9512
rect 17184 9500 17190 9512
rect 19536 9500 19564 9531
rect 20806 9528 20812 9540
rect 20864 9528 20870 9580
rect 20898 9528 20904 9580
rect 20956 9528 20962 9580
rect 21269 9571 21327 9577
rect 21269 9537 21281 9571
rect 21315 9568 21327 9571
rect 21542 9568 21548 9580
rect 21315 9540 21548 9568
rect 21315 9537 21327 9540
rect 21269 9531 21327 9537
rect 21542 9528 21548 9540
rect 21600 9568 21606 9580
rect 21910 9568 21916 9580
rect 21600 9540 21916 9568
rect 21600 9528 21606 9540
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 22112 9577 22140 9608
rect 23290 9596 23296 9648
rect 23348 9596 23354 9648
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22462 9528 22468 9580
rect 22520 9568 22526 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 22520 9540 23949 9568
rect 22520 9528 22526 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 21361 9503 21419 9509
rect 21361 9500 21373 9503
rect 17184 9472 18828 9500
rect 19536 9472 21373 9500
rect 17184 9460 17190 9472
rect 16206 9392 16212 9444
rect 16264 9432 16270 9444
rect 18693 9435 18751 9441
rect 18693 9432 18705 9435
rect 16264 9404 18705 9432
rect 16264 9392 16270 9404
rect 18693 9401 18705 9404
rect 18739 9401 18751 9435
rect 18693 9395 18751 9401
rect 18046 9324 18052 9376
rect 18104 9324 18110 9376
rect 18800 9364 18828 9472
rect 21361 9469 21373 9472
rect 21407 9500 21419 9503
rect 22278 9500 22284 9512
rect 21407 9472 22284 9500
rect 21407 9469 21419 9472
rect 21361 9463 21419 9469
rect 22278 9460 22284 9472
rect 22336 9460 22342 9512
rect 24762 9460 24768 9512
rect 24820 9460 24826 9512
rect 19337 9435 19395 9441
rect 19337 9401 19349 9435
rect 19383 9432 19395 9435
rect 19426 9432 19432 9444
rect 19383 9404 19432 9432
rect 19383 9401 19395 9404
rect 19337 9395 19395 9401
rect 19426 9392 19432 9404
rect 19484 9392 19490 9444
rect 20717 9435 20775 9441
rect 19536 9404 20116 9432
rect 19536 9364 19564 9404
rect 18800 9336 19564 9364
rect 19978 9324 19984 9376
rect 20036 9324 20042 9376
rect 20088 9364 20116 9404
rect 20717 9401 20729 9435
rect 20763 9432 20775 9435
rect 20763 9404 21496 9432
rect 20763 9401 20775 9404
rect 20717 9395 20775 9401
rect 20898 9364 20904 9376
rect 20088 9336 20904 9364
rect 20898 9324 20904 9336
rect 20956 9324 20962 9376
rect 21468 9364 21496 9404
rect 22462 9392 22468 9444
rect 22520 9432 22526 9444
rect 24946 9432 24952 9444
rect 22520 9404 24952 9432
rect 22520 9392 22526 9404
rect 24946 9392 24952 9404
rect 25004 9392 25010 9444
rect 24578 9364 24584 9376
rect 21468 9336 24584 9364
rect 24578 9324 24584 9336
rect 24636 9324 24642 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 11793 9163 11851 9169
rect 11793 9129 11805 9163
rect 11839 9160 11851 9163
rect 14458 9160 14464 9172
rect 11839 9132 14464 9160
rect 11839 9129 11851 9132
rect 11793 9123 11851 9129
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 18046 9120 18052 9172
rect 18104 9160 18110 9172
rect 18104 9132 22094 9160
rect 18104 9120 18110 9132
rect 19061 9095 19119 9101
rect 19061 9061 19073 9095
rect 19107 9092 19119 9095
rect 19334 9092 19340 9104
rect 19107 9064 19340 9092
rect 19107 9061 19119 9064
rect 19061 9055 19119 9061
rect 19334 9052 19340 9064
rect 19392 9052 19398 9104
rect 21269 9095 21327 9101
rect 21269 9092 21281 9095
rect 19444 9064 21281 9092
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 19444 9033 19472 9064
rect 21269 9061 21281 9064
rect 21315 9061 21327 9095
rect 22066 9092 22094 9132
rect 22278 9120 22284 9172
rect 22336 9160 22342 9172
rect 24765 9163 24823 9169
rect 24765 9160 24777 9163
rect 22336 9132 24777 9160
rect 22336 9120 22342 9132
rect 24765 9129 24777 9132
rect 24811 9129 24823 9163
rect 24765 9123 24823 9129
rect 22646 9092 22652 9104
rect 22066 9064 22652 9092
rect 21269 9055 21327 9061
rect 22646 9052 22652 9064
rect 22704 9052 22710 9104
rect 19429 9027 19487 9033
rect 19429 8993 19441 9027
rect 19475 8993 19487 9027
rect 19429 8987 19487 8993
rect 20622 8984 20628 9036
rect 20680 9024 20686 9036
rect 23845 9027 23903 9033
rect 20680 8996 22140 9024
rect 20680 8984 20686 8996
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8956 19763 8959
rect 20898 8956 20904 8968
rect 19751 8928 20904 8956
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 20898 8916 20904 8928
rect 20956 8916 20962 8968
rect 21450 8916 21456 8968
rect 21508 8916 21514 8968
rect 22112 8965 22140 8996
rect 23845 8993 23857 9027
rect 23891 9024 23903 9027
rect 24854 9024 24860 9036
rect 23891 8996 24860 9024
rect 23891 8993 23903 8996
rect 23845 8987 23903 8993
rect 24854 8984 24860 8996
rect 24912 8984 24918 9036
rect 22097 8959 22155 8965
rect 22097 8925 22109 8959
rect 22143 8925 22155 8959
rect 22097 8919 22155 8925
rect 22646 8916 22652 8968
rect 22704 8916 22710 8968
rect 6822 8848 6828 8900
rect 6880 8888 6886 8900
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 6880 8860 10333 8888
rect 6880 8848 6886 8860
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 12069 8891 12127 8897
rect 12069 8888 12081 8891
rect 11546 8860 12081 8888
rect 10321 8851 10379 8857
rect 12069 8857 12081 8860
rect 12115 8888 12127 8891
rect 12526 8888 12532 8900
rect 12115 8860 12532 8888
rect 12115 8857 12127 8860
rect 12069 8851 12127 8857
rect 12526 8848 12532 8860
rect 12584 8848 12590 8900
rect 24673 8891 24731 8897
rect 24673 8857 24685 8891
rect 24719 8857 24731 8891
rect 24673 8851 24731 8857
rect 21913 8823 21971 8829
rect 21913 8789 21925 8823
rect 21959 8820 21971 8823
rect 24688 8820 24716 8851
rect 21959 8792 24716 8820
rect 21959 8789 21971 8792
rect 21913 8783 21971 8789
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 19429 8619 19487 8625
rect 19429 8585 19441 8619
rect 19475 8616 19487 8619
rect 19886 8616 19892 8628
rect 19475 8588 19892 8616
rect 19475 8585 19487 8588
rect 19429 8579 19487 8585
rect 19886 8576 19892 8588
rect 19944 8576 19950 8628
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 21637 8619 21695 8625
rect 20036 8588 21404 8616
rect 20036 8576 20042 8588
rect 21376 8548 21404 8588
rect 21637 8585 21649 8619
rect 21683 8616 21695 8619
rect 22370 8616 22376 8628
rect 21683 8588 22376 8616
rect 21683 8585 21695 8588
rect 21637 8579 21695 8585
rect 22370 8576 22376 8588
rect 22428 8576 22434 8628
rect 20272 8520 21312 8548
rect 21376 8520 22600 8548
rect 13538 8440 13544 8492
rect 13596 8480 13602 8492
rect 20272 8489 20300 8520
rect 21284 8489 21312 8520
rect 19613 8483 19671 8489
rect 19613 8480 19625 8483
rect 13596 8452 19625 8480
rect 13596 8440 13602 8452
rect 19613 8449 19625 8452
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 20901 8483 20959 8489
rect 20901 8449 20913 8483
rect 20947 8449 20959 8483
rect 20901 8443 20959 8449
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 22002 8480 22008 8492
rect 21315 8452 22008 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 19058 8372 19064 8424
rect 19116 8412 19122 8424
rect 20916 8412 20944 8443
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 22281 8483 22339 8489
rect 22281 8449 22293 8483
rect 22327 8480 22339 8483
rect 22462 8480 22468 8492
rect 22327 8452 22468 8480
rect 22327 8449 22339 8452
rect 22281 8443 22339 8449
rect 22462 8440 22468 8452
rect 22520 8440 22526 8492
rect 22572 8480 22600 8520
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 22572 8452 23949 8480
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 24946 8480 24952 8492
rect 23937 8443 23995 8449
rect 24688 8452 24952 8480
rect 19116 8384 20944 8412
rect 23293 8415 23351 8421
rect 19116 8372 19122 8384
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 24688 8412 24716 8452
rect 24946 8440 24952 8452
rect 25004 8440 25010 8492
rect 23339 8384 24716 8412
rect 24765 8415 24823 8421
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 24765 8381 24777 8415
rect 24811 8381 24823 8415
rect 24765 8375 24823 8381
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 19300 8316 20085 8344
rect 19300 8304 19306 8316
rect 20073 8313 20085 8316
rect 20119 8313 20131 8347
rect 20073 8307 20131 8313
rect 20717 8347 20775 8353
rect 20717 8313 20729 8347
rect 20763 8344 20775 8347
rect 20763 8316 24624 8344
rect 20763 8313 20775 8316
rect 20717 8307 20775 8313
rect 24596 8276 24624 8316
rect 24670 8304 24676 8356
rect 24728 8344 24734 8356
rect 24780 8344 24808 8375
rect 24728 8316 24808 8344
rect 24728 8304 24734 8316
rect 24854 8304 24860 8356
rect 24912 8304 24918 8356
rect 24872 8276 24900 8304
rect 24596 8248 24900 8276
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 21361 8075 21419 8081
rect 21361 8041 21373 8075
rect 21407 8072 21419 8075
rect 23934 8072 23940 8084
rect 21407 8044 23940 8072
rect 21407 8041 21419 8044
rect 21361 8035 21419 8041
rect 23934 8032 23940 8044
rect 23992 8032 23998 8084
rect 15102 7964 15108 8016
rect 15160 8004 15166 8016
rect 22005 8007 22063 8013
rect 22005 8004 22017 8007
rect 15160 7976 22017 8004
rect 15160 7964 15166 7976
rect 22005 7973 22017 7976
rect 22051 7973 22063 8007
rect 22005 7967 22063 7973
rect 23474 7936 23480 7948
rect 22066 7908 23480 7936
rect 18690 7828 18696 7880
rect 18748 7868 18754 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 18748 7840 20913 7868
rect 18748 7828 18754 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7868 21603 7871
rect 22066 7868 22094 7908
rect 23474 7896 23480 7908
rect 23532 7896 23538 7948
rect 23845 7939 23903 7945
rect 23845 7905 23857 7939
rect 23891 7936 23903 7939
rect 24946 7936 24952 7948
rect 23891 7908 24952 7936
rect 23891 7905 23903 7908
rect 23845 7899 23903 7905
rect 24946 7896 24952 7908
rect 25004 7896 25010 7948
rect 21591 7840 22094 7868
rect 22189 7871 22247 7877
rect 21591 7837 21603 7840
rect 21545 7831 21603 7837
rect 22189 7837 22201 7871
rect 22235 7868 22247 7871
rect 22370 7868 22376 7880
rect 22235 7840 22376 7868
rect 22235 7837 22247 7840
rect 22189 7831 22247 7837
rect 22370 7828 22376 7840
rect 22428 7828 22434 7880
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7837 22891 7871
rect 22833 7831 22891 7837
rect 24857 7871 24915 7877
rect 24857 7837 24869 7871
rect 24903 7868 24915 7871
rect 25038 7868 25044 7880
rect 24903 7840 25044 7868
rect 24903 7837 24915 7840
rect 24857 7831 24915 7837
rect 22848 7800 22876 7831
rect 25038 7828 25044 7840
rect 25096 7828 25102 7880
rect 25866 7800 25872 7812
rect 22848 7772 25872 7800
rect 25866 7760 25872 7772
rect 25924 7760 25930 7812
rect 20714 7692 20720 7744
rect 20772 7692 20778 7744
rect 23474 7692 23480 7744
rect 23532 7732 23538 7744
rect 24673 7735 24731 7741
rect 24673 7732 24685 7735
rect 23532 7704 24685 7732
rect 23532 7692 23538 7704
rect 24673 7701 24685 7704
rect 24719 7701 24731 7735
rect 24673 7695 24731 7701
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 21269 7531 21327 7537
rect 21269 7497 21281 7531
rect 21315 7528 21327 7531
rect 22646 7528 22652 7540
rect 21315 7500 22652 7528
rect 21315 7497 21327 7500
rect 21269 7491 21327 7497
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 20714 7420 20720 7472
rect 20772 7460 20778 7472
rect 23293 7463 23351 7469
rect 20772 7432 23060 7460
rect 20772 7420 20778 7432
rect 20254 7352 20260 7404
rect 20312 7392 20318 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20312 7364 20821 7392
rect 20312 7352 20318 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 21082 7352 21088 7404
rect 21140 7392 21146 7404
rect 21453 7395 21511 7401
rect 21453 7392 21465 7395
rect 21140 7364 21465 7392
rect 21140 7352 21146 7364
rect 21453 7361 21465 7364
rect 21499 7361 21511 7395
rect 21453 7355 21511 7361
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7361 22339 7395
rect 23032 7392 23060 7432
rect 23293 7429 23305 7463
rect 23339 7460 23351 7463
rect 24854 7460 24860 7472
rect 23339 7432 24860 7460
rect 23339 7429 23351 7432
rect 23293 7423 23351 7429
rect 24854 7420 24860 7432
rect 24912 7420 24918 7472
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 23032 7364 23949 7392
rect 22281 7355 22339 7361
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 22296 7324 22324 7355
rect 25682 7324 25688 7336
rect 22296 7296 25688 7324
rect 25682 7284 25688 7296
rect 25740 7284 25746 7336
rect 20625 7259 20683 7265
rect 20625 7225 20637 7259
rect 20671 7256 20683 7259
rect 23382 7256 23388 7268
rect 20671 7228 23388 7256
rect 20671 7225 20683 7228
rect 20625 7219 20683 7225
rect 23382 7216 23388 7228
rect 23440 7216 23446 7268
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 23845 6851 23903 6857
rect 23845 6817 23857 6851
rect 23891 6848 23903 6851
rect 24854 6848 24860 6860
rect 23891 6820 24860 6848
rect 23891 6817 23903 6820
rect 23845 6811 23903 6817
rect 24854 6808 24860 6820
rect 24912 6808 24918 6860
rect 21174 6740 21180 6792
rect 21232 6780 21238 6792
rect 21545 6783 21603 6789
rect 21545 6780 21557 6783
rect 21232 6752 21557 6780
rect 21232 6740 21238 6752
rect 21545 6749 21557 6752
rect 21591 6749 21603 6783
rect 22649 6783 22707 6789
rect 22649 6780 22661 6783
rect 21545 6743 21603 6749
rect 22066 6752 22661 6780
rect 22066 6712 22094 6752
rect 22649 6749 22661 6752
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 24578 6740 24584 6792
rect 24636 6780 24642 6792
rect 24673 6783 24731 6789
rect 24673 6780 24685 6783
rect 24636 6752 24685 6780
rect 24636 6740 24642 6752
rect 24673 6749 24685 6752
rect 24719 6749 24731 6783
rect 24673 6743 24731 6749
rect 21376 6684 22094 6712
rect 24857 6715 24915 6721
rect 21376 6653 21404 6684
rect 24857 6681 24869 6715
rect 24903 6712 24915 6715
rect 25038 6712 25044 6724
rect 24903 6684 25044 6712
rect 24903 6681 24915 6684
rect 24857 6675 24915 6681
rect 25038 6672 25044 6684
rect 25096 6672 25102 6724
rect 21361 6647 21419 6653
rect 21361 6613 21373 6647
rect 21407 6613 21419 6647
rect 21361 6607 21419 6613
rect 22005 6647 22063 6653
rect 22005 6613 22017 6647
rect 22051 6644 22063 6647
rect 25222 6644 25228 6656
rect 22051 6616 25228 6644
rect 22051 6613 22063 6616
rect 22005 6607 22063 6613
rect 25222 6604 25228 6616
rect 25280 6604 25286 6656
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 23293 6375 23351 6381
rect 23293 6341 23305 6375
rect 23339 6372 23351 6375
rect 24854 6372 24860 6384
rect 23339 6344 24860 6372
rect 23339 6341 23351 6344
rect 23293 6335 23351 6341
rect 24854 6332 24860 6344
rect 24912 6332 24918 6384
rect 22278 6264 22284 6316
rect 22336 6264 22342 6316
rect 24121 6307 24179 6313
rect 24121 6273 24133 6307
rect 24167 6304 24179 6307
rect 25590 6304 25596 6316
rect 24167 6276 25596 6304
rect 24167 6273 24179 6276
rect 24121 6267 24179 6273
rect 25590 6264 25596 6276
rect 25648 6264 25654 6316
rect 24762 6196 24768 6248
rect 24820 6196 24826 6248
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 22002 5856 22008 5908
rect 22060 5856 22066 5908
rect 21361 5831 21419 5837
rect 21361 5797 21373 5831
rect 21407 5828 21419 5831
rect 23658 5828 23664 5840
rect 21407 5800 23664 5828
rect 21407 5797 21419 5800
rect 21361 5791 21419 5797
rect 23658 5788 23664 5800
rect 23716 5788 23722 5840
rect 22370 5760 22376 5772
rect 22204 5732 22376 5760
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5692 21603 5695
rect 21818 5692 21824 5704
rect 21591 5664 21824 5692
rect 21591 5661 21603 5664
rect 21545 5655 21603 5661
rect 21818 5652 21824 5664
rect 21876 5652 21882 5704
rect 22204 5701 22232 5732
rect 22370 5720 22376 5732
rect 22428 5760 22434 5772
rect 23290 5760 23296 5772
rect 22428 5732 23296 5760
rect 22428 5720 22434 5732
rect 23290 5720 23296 5732
rect 23348 5720 23354 5772
rect 24946 5720 24952 5772
rect 25004 5720 25010 5772
rect 22189 5695 22247 5701
rect 22189 5661 22201 5695
rect 22235 5661 22247 5695
rect 22189 5655 22247 5661
rect 22833 5695 22891 5701
rect 22833 5661 22845 5695
rect 22879 5692 22891 5695
rect 23474 5692 23480 5704
rect 22879 5664 23480 5692
rect 22879 5661 22891 5664
rect 22833 5655 22891 5661
rect 23474 5652 23480 5664
rect 23532 5652 23538 5704
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5692 24915 5695
rect 24964 5692 24992 5720
rect 24903 5664 24992 5692
rect 24903 5661 24915 5664
rect 24857 5655 24915 5661
rect 23845 5627 23903 5633
rect 23845 5593 23857 5627
rect 23891 5624 23903 5627
rect 24946 5624 24952 5636
rect 23891 5596 24952 5624
rect 23891 5593 23903 5596
rect 23845 5587 23903 5593
rect 24946 5584 24952 5596
rect 25004 5584 25010 5636
rect 23474 5516 23480 5568
rect 23532 5556 23538 5568
rect 24673 5559 24731 5565
rect 24673 5556 24685 5559
rect 23532 5528 24685 5556
rect 23532 5516 23538 5528
rect 24673 5525 24685 5528
rect 24719 5525 24731 5559
rect 24673 5519 24731 5525
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 20898 5244 20904 5296
rect 20956 5284 20962 5296
rect 20956 5256 23980 5284
rect 20956 5244 20962 5256
rect 22281 5219 22339 5225
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 22738 5216 22744 5228
rect 22327 5188 22744 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 22738 5176 22744 5188
rect 22796 5176 22802 5228
rect 23952 5225 23980 5256
rect 23937 5219 23995 5225
rect 23937 5185 23949 5219
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 23293 5151 23351 5157
rect 23293 5117 23305 5151
rect 23339 5117 23351 5151
rect 23293 5111 23351 5117
rect 23308 5080 23336 5111
rect 24670 5108 24676 5160
rect 24728 5108 24734 5160
rect 24946 5080 24952 5092
rect 23308 5052 24952 5080
rect 24946 5040 24952 5052
rect 25004 5040 25010 5092
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 22370 4768 22376 4820
rect 22428 4768 22434 4820
rect 22646 4564 22652 4616
rect 22704 4564 22710 4616
rect 23382 4564 23388 4616
rect 23440 4604 23446 4616
rect 24857 4607 24915 4613
rect 24857 4604 24869 4607
rect 23440 4576 24869 4604
rect 23440 4564 23446 4576
rect 24857 4573 24869 4576
rect 24903 4573 24915 4607
rect 24857 4567 24915 4573
rect 23845 4539 23903 4545
rect 23845 4505 23857 4539
rect 23891 4536 23903 4539
rect 24946 4536 24952 4548
rect 23891 4508 24952 4536
rect 23891 4505 23903 4508
rect 23845 4499 23903 4505
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 23566 4428 23572 4480
rect 23624 4468 23630 4480
rect 24673 4471 24731 4477
rect 24673 4468 24685 4471
rect 23624 4440 24685 4468
rect 23624 4428 23630 4440
rect 24673 4437 24685 4440
rect 24719 4437 24731 4471
rect 24673 4431 24731 4437
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 23952 4168 25176 4196
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 21910 4128 21916 4140
rect 20303 4100 21916 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 21910 4088 21916 4100
rect 21968 4088 21974 4140
rect 23952 4137 23980 4168
rect 22281 4131 22339 4137
rect 22281 4097 22293 4131
rect 22327 4128 22339 4131
rect 23937 4131 23995 4137
rect 22327 4100 23428 4128
rect 22327 4097 22339 4100
rect 22281 4091 22339 4097
rect 18966 4020 18972 4072
rect 19024 4060 19030 4072
rect 20162 4060 20168 4072
rect 19024 4032 20168 4060
rect 19024 4020 19030 4032
rect 20162 4020 20168 4032
rect 20220 4020 20226 4072
rect 21269 4063 21327 4069
rect 21269 4029 21281 4063
rect 21315 4060 21327 4063
rect 23293 4063 23351 4069
rect 21315 4032 22094 4060
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 22066 4004 22094 4032
rect 23293 4029 23305 4063
rect 23339 4029 23351 4063
rect 23400 4060 23428 4100
rect 23937 4097 23949 4131
rect 23983 4097 23995 4131
rect 25038 4128 25044 4140
rect 23937 4091 23995 4097
rect 24044 4100 25044 4128
rect 24044 4060 24072 4100
rect 25038 4088 25044 4100
rect 25096 4088 25102 4140
rect 25148 4128 25176 4168
rect 25774 4128 25780 4140
rect 25148 4100 25780 4128
rect 25774 4088 25780 4100
rect 25832 4088 25838 4140
rect 23400 4032 24072 4060
rect 23293 4023 23351 4029
rect 22066 3964 22100 4004
rect 22094 3952 22100 3964
rect 22152 3952 22158 4004
rect 23308 3992 23336 4023
rect 24762 4020 24768 4072
rect 24820 4020 24826 4072
rect 24946 3992 24952 4004
rect 23308 3964 24952 3992
rect 24946 3952 24952 3964
rect 25004 3952 25010 4004
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 20530 3476 20536 3528
rect 20588 3516 20594 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 20588 3488 20821 3516
rect 20588 3476 20594 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 23474 3516 23480 3528
rect 22879 3488 23480 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 23474 3476 23480 3488
rect 23532 3476 23538 3528
rect 23658 3476 23664 3528
rect 23716 3516 23722 3528
rect 24765 3519 24823 3525
rect 24765 3516 24777 3519
rect 23716 3488 24777 3516
rect 23716 3476 23722 3488
rect 24765 3485 24777 3488
rect 24811 3485 24823 3519
rect 24765 3479 24823 3485
rect 22002 3408 22008 3460
rect 22060 3408 22066 3460
rect 23845 3451 23903 3457
rect 23845 3417 23857 3451
rect 23891 3448 23903 3451
rect 25130 3448 25136 3460
rect 23891 3420 25136 3448
rect 23891 3417 23903 3420
rect 23845 3411 23903 3417
rect 25130 3408 25136 3420
rect 25188 3408 25194 3460
rect 24578 3340 24584 3392
rect 24636 3340 24642 3392
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 25314 3176 25320 3188
rect 22066 3148 25320 3176
rect 22066 3108 22094 3148
rect 25314 3136 25320 3148
rect 25372 3136 25378 3188
rect 18432 3080 22094 3108
rect 23293 3111 23351 3117
rect 18432 3049 18460 3080
rect 23293 3077 23305 3111
rect 23339 3108 23351 3111
rect 24854 3108 24860 3120
rect 23339 3080 24860 3108
rect 23339 3077 23351 3080
rect 23293 3071 23351 3077
rect 24854 3068 24860 3080
rect 24912 3068 24918 3120
rect 25133 3111 25191 3117
rect 25133 3077 25145 3111
rect 25179 3108 25191 3111
rect 25222 3108 25228 3120
rect 25179 3080 25228 3108
rect 25179 3077 25191 3080
rect 25133 3071 25191 3077
rect 25222 3068 25228 3080
rect 25280 3068 25286 3120
rect 18417 3043 18475 3049
rect 18417 3009 18429 3043
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 19610 3000 19616 3052
rect 19668 3040 19674 3052
rect 20073 3043 20131 3049
rect 20073 3040 20085 3043
rect 19668 3012 20085 3040
rect 19668 3000 19674 3012
rect 20073 3009 20085 3012
rect 20119 3009 20131 3043
rect 20073 3003 20131 3009
rect 22281 3043 22339 3049
rect 22281 3009 22293 3043
rect 22327 3040 22339 3043
rect 23566 3040 23572 3052
rect 22327 3012 23572 3040
rect 22327 3009 22339 3012
rect 22281 3003 22339 3009
rect 23566 3000 23572 3012
rect 23624 3000 23630 3052
rect 24118 3000 24124 3052
rect 24176 3000 24182 3052
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2972 19487 2975
rect 19518 2972 19524 2984
rect 19475 2944 19524 2972
rect 19475 2941 19487 2944
rect 19429 2935 19487 2941
rect 19518 2932 19524 2944
rect 19576 2932 19582 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 25038 2972 25044 2984
rect 21315 2944 25044 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 25038 2932 25044 2944
rect 25096 2932 25102 2984
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 6822 2592 6828 2644
rect 6880 2592 6886 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 22186 2632 22192 2644
rect 19576 2604 22192 2632
rect 19576 2592 19582 2604
rect 22186 2592 22192 2604
rect 22244 2592 22250 2644
rect 6914 2388 6920 2440
rect 6972 2428 6978 2440
rect 7009 2431 7067 2437
rect 7009 2428 7021 2431
rect 6972 2400 7021 2428
rect 6972 2388 6978 2400
rect 7009 2397 7021 2400
rect 7055 2428 7067 2431
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 7055 2400 7297 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2428 20315 2431
rect 22738 2428 22744 2440
rect 20303 2400 22744 2428
rect 20303 2397 20315 2400
rect 20257 2391 20315 2397
rect 22738 2388 22744 2400
rect 22796 2388 22802 2440
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2428 22891 2431
rect 24578 2428 24584 2440
rect 22879 2400 24584 2428
rect 22879 2397 22891 2400
rect 22833 2391 22891 2397
rect 24578 2388 24584 2400
rect 24636 2388 24642 2440
rect 21269 2363 21327 2369
rect 21269 2329 21281 2363
rect 21315 2360 21327 2363
rect 23382 2360 23388 2372
rect 21315 2332 23388 2360
rect 21315 2329 21327 2332
rect 21269 2323 21327 2329
rect 23382 2320 23388 2332
rect 23440 2320 23446 2372
rect 23845 2363 23903 2369
rect 23845 2329 23857 2363
rect 23891 2360 23903 2363
rect 24946 2360 24952 2372
rect 23891 2332 24952 2360
rect 23891 2329 23903 2332
rect 23845 2323 23903 2329
rect 24946 2320 24952 2332
rect 25004 2320 25010 2372
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
<< via1 >>
rect 3056 26392 3108 26444
rect 3332 26392 3384 26444
rect 5448 26324 5500 26376
rect 21272 26324 21324 26376
rect 4896 26256 4948 26308
rect 20168 26256 20220 26308
rect 6000 25032 6052 25084
rect 13728 25032 13780 25084
rect 9128 24964 9180 25016
rect 20352 24964 20404 25016
rect 1952 24896 2004 24948
rect 16028 24896 16080 24948
rect 6736 24828 6788 24880
rect 26148 24828 26200 24880
rect 14096 24692 14148 24744
rect 23388 24692 23440 24744
rect 16856 24624 16908 24676
rect 24860 24624 24912 24676
rect 4804 24556 4856 24608
rect 12624 24556 12676 24608
rect 16948 24556 17000 24608
rect 24952 24556 25004 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 6552 24395 6604 24404
rect 6552 24361 6561 24395
rect 6561 24361 6595 24395
rect 6595 24361 6604 24395
rect 6552 24352 6604 24361
rect 6644 24352 6696 24404
rect 16948 24395 17000 24404
rect 16948 24361 16957 24395
rect 16957 24361 16991 24395
rect 16991 24361 17000 24395
rect 16948 24352 17000 24361
rect 4988 24284 5040 24336
rect 6184 24216 6236 24268
rect 3884 24148 3936 24200
rect 4160 24191 4212 24200
rect 4160 24157 4169 24191
rect 4169 24157 4203 24191
rect 4203 24157 4212 24191
rect 4160 24148 4212 24157
rect 6644 24148 6696 24200
rect 7012 24148 7064 24200
rect 9128 24327 9180 24336
rect 9128 24293 9137 24327
rect 9137 24293 9171 24327
rect 9171 24293 9180 24327
rect 9128 24284 9180 24293
rect 11704 24327 11756 24336
rect 11704 24293 11713 24327
rect 11713 24293 11747 24327
rect 11747 24293 11756 24327
rect 11704 24284 11756 24293
rect 12348 24284 12400 24336
rect 9680 24216 9732 24268
rect 11244 24216 11296 24268
rect 16396 24284 16448 24336
rect 8668 24080 8720 24132
rect 9496 24148 9548 24200
rect 12440 24191 12492 24200
rect 12440 24157 12449 24191
rect 12449 24157 12483 24191
rect 12483 24157 12492 24191
rect 12440 24148 12492 24157
rect 16028 24259 16080 24268
rect 16028 24225 16037 24259
rect 16037 24225 16071 24259
rect 16071 24225 16080 24259
rect 16028 24216 16080 24225
rect 19156 24352 19208 24404
rect 22008 24352 22060 24404
rect 18052 24284 18104 24336
rect 17960 24216 18012 24268
rect 18236 24284 18288 24336
rect 21732 24284 21784 24336
rect 18788 24259 18840 24268
rect 18788 24225 18797 24259
rect 18797 24225 18831 24259
rect 18831 24225 18840 24259
rect 18788 24216 18840 24225
rect 24308 24352 24360 24404
rect 24400 24395 24452 24404
rect 24400 24361 24409 24395
rect 24409 24361 24443 24395
rect 24443 24361 24452 24395
rect 24400 24352 24452 24361
rect 15108 24148 15160 24200
rect 23204 24216 23256 24268
rect 12808 24080 12860 24132
rect 14556 24080 14608 24132
rect 6460 24012 6512 24064
rect 10232 24012 10284 24064
rect 15016 24080 15068 24132
rect 20812 24148 20864 24200
rect 22284 24191 22336 24200
rect 22284 24157 22293 24191
rect 22293 24157 22327 24191
rect 22327 24157 22336 24191
rect 22284 24148 22336 24157
rect 24400 24148 24452 24200
rect 20904 24080 20956 24132
rect 22652 24080 22704 24132
rect 23940 24080 23992 24132
rect 16948 24012 17000 24064
rect 17408 24055 17460 24064
rect 17408 24021 17417 24055
rect 17417 24021 17451 24055
rect 17451 24021 17460 24055
rect 17408 24012 17460 24021
rect 17684 24012 17736 24064
rect 19248 24012 19300 24064
rect 19800 24012 19852 24064
rect 23204 24012 23256 24064
rect 23572 24012 23624 24064
rect 24492 24012 24544 24064
rect 25412 24055 25464 24064
rect 25412 24021 25421 24055
rect 25421 24021 25455 24055
rect 25455 24021 25464 24055
rect 25412 24012 25464 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 1308 23672 1360 23724
rect 5172 23740 5224 23792
rect 7564 23740 7616 23792
rect 10140 23740 10192 23792
rect 10876 23783 10928 23792
rect 10876 23749 10885 23783
rect 10885 23749 10919 23783
rect 10919 23749 10928 23783
rect 10876 23740 10928 23749
rect 13728 23808 13780 23860
rect 15016 23808 15068 23860
rect 15384 23808 15436 23860
rect 17684 23808 17736 23860
rect 17316 23740 17368 23792
rect 4804 23715 4856 23724
rect 4804 23681 4813 23715
rect 4813 23681 4847 23715
rect 4847 23681 4856 23715
rect 4804 23672 4856 23681
rect 5448 23672 5500 23724
rect 6644 23604 6696 23656
rect 6736 23604 6788 23656
rect 6920 23604 6972 23656
rect 7104 23536 7156 23588
rect 7840 23604 7892 23656
rect 16120 23672 16172 23724
rect 17132 23672 17184 23724
rect 17868 23672 17920 23724
rect 11980 23604 12032 23656
rect 12808 23536 12860 23588
rect 14740 23647 14792 23656
rect 14740 23613 14749 23647
rect 14749 23613 14783 23647
rect 14783 23613 14792 23647
rect 14740 23604 14792 23613
rect 14924 23604 14976 23656
rect 20812 23740 20864 23792
rect 23572 23808 23624 23860
rect 24308 23851 24360 23860
rect 24308 23817 24317 23851
rect 24317 23817 24351 23851
rect 24351 23817 24360 23851
rect 24308 23808 24360 23817
rect 23940 23740 23992 23792
rect 24584 23740 24636 23792
rect 24768 23783 24820 23792
rect 24768 23749 24777 23783
rect 24777 23749 24811 23783
rect 24811 23749 24820 23783
rect 24768 23740 24820 23749
rect 18052 23715 18104 23724
rect 18052 23681 18061 23715
rect 18061 23681 18095 23715
rect 18095 23681 18104 23715
rect 18052 23672 18104 23681
rect 22008 23672 22060 23724
rect 18788 23604 18840 23656
rect 20720 23604 20772 23656
rect 20904 23647 20956 23656
rect 20904 23613 20913 23647
rect 20913 23613 20947 23647
rect 20947 23613 20956 23647
rect 20904 23604 20956 23613
rect 22284 23647 22336 23656
rect 22284 23613 22293 23647
rect 22293 23613 22327 23647
rect 22327 23613 22336 23647
rect 22284 23604 22336 23613
rect 22560 23647 22612 23656
rect 17776 23536 17828 23588
rect 7012 23468 7064 23520
rect 13636 23468 13688 23520
rect 15844 23468 15896 23520
rect 16856 23511 16908 23520
rect 16856 23477 16865 23511
rect 16865 23477 16899 23511
rect 16899 23477 16908 23511
rect 16856 23468 16908 23477
rect 16948 23468 17000 23520
rect 20260 23536 20312 23588
rect 21732 23536 21784 23588
rect 22560 23613 22569 23647
rect 22569 23613 22603 23647
rect 22603 23613 22612 23647
rect 22560 23604 22612 23613
rect 22652 23604 22704 23656
rect 25504 23604 25556 23656
rect 19800 23511 19852 23520
rect 19800 23477 19809 23511
rect 19809 23477 19843 23511
rect 19843 23477 19852 23511
rect 19800 23468 19852 23477
rect 21640 23468 21692 23520
rect 24584 23511 24636 23520
rect 24584 23477 24593 23511
rect 24593 23477 24627 23511
rect 24627 23477 24636 23511
rect 24584 23468 24636 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 6644 23264 6696 23316
rect 7380 23264 7432 23316
rect 11796 23264 11848 23316
rect 7288 23196 7340 23248
rect 7472 23196 7524 23248
rect 2780 23128 2832 23180
rect 8392 23128 8444 23180
rect 9220 23128 9272 23180
rect 5908 23060 5960 23112
rect 9312 23060 9364 23112
rect 4344 22992 4396 23044
rect 6276 22992 6328 23044
rect 4712 22967 4764 22976
rect 4712 22933 4721 22967
rect 4721 22933 4755 22967
rect 4755 22933 4764 22967
rect 4712 22924 4764 22933
rect 6460 22992 6512 23044
rect 12532 23196 12584 23248
rect 13452 23196 13504 23248
rect 13636 23264 13688 23316
rect 14832 23264 14884 23316
rect 16304 23264 16356 23316
rect 17960 23264 18012 23316
rect 24492 23264 24544 23316
rect 16948 23196 17000 23248
rect 19340 23196 19392 23248
rect 20720 23196 20772 23248
rect 23388 23196 23440 23248
rect 10508 23171 10560 23180
rect 10508 23137 10517 23171
rect 10517 23137 10551 23171
rect 10551 23137 10560 23171
rect 10508 23128 10560 23137
rect 11612 23128 11664 23180
rect 7656 22924 7708 22976
rect 11796 23060 11848 23112
rect 13912 23128 13964 23180
rect 17132 23128 17184 23180
rect 17408 23128 17460 23180
rect 17868 23171 17920 23180
rect 17868 23137 17877 23171
rect 17877 23137 17911 23171
rect 17911 23137 17920 23171
rect 17868 23128 17920 23137
rect 18420 23128 18472 23180
rect 18696 23128 18748 23180
rect 20996 23128 21048 23180
rect 22284 23128 22336 23180
rect 23296 23128 23348 23180
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 14280 23060 14332 23112
rect 17960 23060 18012 23112
rect 18052 23060 18104 23112
rect 19340 23060 19392 23112
rect 20812 23060 20864 23112
rect 21272 23060 21324 23112
rect 23204 23060 23256 23112
rect 13452 22992 13504 23044
rect 13544 22967 13596 22976
rect 13544 22933 13553 22967
rect 13553 22933 13587 22967
rect 13587 22933 13596 22967
rect 13544 22924 13596 22933
rect 14372 23035 14424 23044
rect 14372 23001 14381 23035
rect 14381 23001 14415 23035
rect 14415 23001 14424 23035
rect 14372 22992 14424 23001
rect 15844 22992 15896 23044
rect 17132 22992 17184 23044
rect 17408 22992 17460 23044
rect 18512 23035 18564 23044
rect 18512 23001 18521 23035
rect 18521 23001 18555 23035
rect 18555 23001 18564 23035
rect 18512 22992 18564 23001
rect 18604 22992 18656 23044
rect 19708 23035 19760 23044
rect 19708 23001 19717 23035
rect 19717 23001 19751 23035
rect 19751 23001 19760 23035
rect 19708 22992 19760 23001
rect 22008 22992 22060 23044
rect 23664 22992 23716 23044
rect 14648 22924 14700 22976
rect 16672 22924 16724 22976
rect 16856 22924 16908 22976
rect 17868 22924 17920 22976
rect 19800 22924 19852 22976
rect 22560 22924 22612 22976
rect 24032 22924 24084 22976
rect 24768 22924 24820 22976
rect 25964 22924 26016 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 2780 22720 2832 22772
rect 4712 22720 4764 22772
rect 12624 22720 12676 22772
rect 4252 22652 4304 22704
rect 5724 22695 5776 22704
rect 5724 22661 5733 22695
rect 5733 22661 5767 22695
rect 5767 22661 5776 22695
rect 5724 22652 5776 22661
rect 7380 22652 7432 22704
rect 8760 22695 8812 22704
rect 8760 22661 8769 22695
rect 8769 22661 8803 22695
rect 8803 22661 8812 22695
rect 8760 22652 8812 22661
rect 10416 22652 10468 22704
rect 11612 22652 11664 22704
rect 13544 22652 13596 22704
rect 14648 22720 14700 22772
rect 14740 22720 14792 22772
rect 15844 22720 15896 22772
rect 18420 22720 18472 22772
rect 1308 22584 1360 22636
rect 3792 22584 3844 22636
rect 6644 22627 6696 22636
rect 6644 22593 6653 22627
rect 6653 22593 6687 22627
rect 6687 22593 6696 22627
rect 6644 22584 6696 22593
rect 5356 22516 5408 22568
rect 9036 22516 9088 22568
rect 12256 22559 12308 22568
rect 12256 22525 12265 22559
rect 12265 22525 12299 22559
rect 12299 22525 12308 22559
rect 12256 22516 12308 22525
rect 12992 22627 13044 22636
rect 12992 22593 13001 22627
rect 13001 22593 13035 22627
rect 13035 22593 13044 22627
rect 12992 22584 13044 22593
rect 13636 22627 13688 22636
rect 13636 22593 13645 22627
rect 13645 22593 13679 22627
rect 13679 22593 13688 22627
rect 13636 22584 13688 22593
rect 15752 22584 15804 22636
rect 16028 22584 16080 22636
rect 16580 22584 16632 22636
rect 4068 22380 4120 22432
rect 4160 22380 4212 22432
rect 11336 22448 11388 22500
rect 11888 22448 11940 22500
rect 12992 22448 13044 22500
rect 11152 22423 11204 22432
rect 11152 22389 11161 22423
rect 11161 22389 11195 22423
rect 11195 22389 11204 22423
rect 11152 22380 11204 22389
rect 11244 22380 11296 22432
rect 13636 22380 13688 22432
rect 14280 22380 14332 22432
rect 16488 22448 16540 22500
rect 17776 22516 17828 22568
rect 19248 22720 19300 22772
rect 20536 22720 20588 22772
rect 19708 22652 19760 22704
rect 20444 22652 20496 22704
rect 19800 22584 19852 22636
rect 20168 22584 20220 22636
rect 16580 22380 16632 22432
rect 16672 22380 16724 22432
rect 19432 22448 19484 22500
rect 19892 22516 19944 22568
rect 21272 22763 21324 22772
rect 21272 22729 21281 22763
rect 21281 22729 21315 22763
rect 21315 22729 21324 22763
rect 21272 22720 21324 22729
rect 23664 22720 23716 22772
rect 24584 22720 24636 22772
rect 23572 22695 23624 22704
rect 23572 22661 23581 22695
rect 23581 22661 23615 22695
rect 23615 22661 23624 22695
rect 23572 22652 23624 22661
rect 22192 22516 22244 22568
rect 22284 22559 22336 22568
rect 22284 22525 22293 22559
rect 22293 22525 22327 22559
rect 22327 22525 22336 22559
rect 22284 22516 22336 22525
rect 23296 22627 23348 22636
rect 23296 22593 23305 22627
rect 23305 22593 23339 22627
rect 23339 22593 23348 22627
rect 23296 22584 23348 22593
rect 25044 22516 25096 22568
rect 23204 22448 23256 22500
rect 20812 22380 20864 22432
rect 21364 22380 21416 22432
rect 22744 22380 22796 22432
rect 25136 22380 25188 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 7656 22176 7708 22228
rect 12072 22176 12124 22228
rect 12164 22176 12216 22228
rect 12532 22176 12584 22228
rect 14648 22176 14700 22228
rect 2412 22108 2464 22160
rect 2780 22108 2832 22160
rect 2872 22083 2924 22092
rect 2872 22049 2881 22083
rect 2881 22049 2915 22083
rect 2915 22049 2924 22083
rect 2872 22040 2924 22049
rect 6092 22083 6144 22092
rect 6092 22049 6101 22083
rect 6101 22049 6135 22083
rect 6135 22049 6144 22083
rect 6092 22040 6144 22049
rect 8300 22083 8352 22092
rect 8300 22049 8309 22083
rect 8309 22049 8343 22083
rect 8343 22049 8352 22083
rect 8300 22040 8352 22049
rect 9036 22040 9088 22092
rect 11060 22040 11112 22092
rect 11336 22040 11388 22092
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 4620 21972 4672 22024
rect 6368 21972 6420 22024
rect 7380 22015 7432 22024
rect 7380 21981 7389 22015
rect 7389 21981 7423 22015
rect 7423 21981 7432 22015
rect 7380 21972 7432 21981
rect 12256 22040 12308 22092
rect 12624 22040 12676 22092
rect 13636 22040 13688 22092
rect 17040 22176 17092 22228
rect 18420 22176 18472 22228
rect 22836 22176 22888 22228
rect 23204 22176 23256 22228
rect 23480 22176 23532 22228
rect 25320 22176 25372 22228
rect 15660 22108 15712 22160
rect 16488 22108 16540 22160
rect 17776 22108 17828 22160
rect 17868 22108 17920 22160
rect 19892 22108 19944 22160
rect 17040 22083 17092 22092
rect 17040 22049 17049 22083
rect 17049 22049 17083 22083
rect 17083 22049 17092 22083
rect 17040 22040 17092 22049
rect 4896 21904 4948 21956
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 10048 21879 10100 21888
rect 10048 21845 10057 21879
rect 10057 21845 10091 21879
rect 10091 21845 10100 21879
rect 10048 21836 10100 21845
rect 14280 22015 14332 22024
rect 14280 21981 14289 22015
rect 14289 21981 14323 22015
rect 14323 21981 14332 22015
rect 14280 21972 14332 21981
rect 15936 21972 15988 22024
rect 18052 22040 18104 22092
rect 20720 22040 20772 22092
rect 23480 22083 23532 22092
rect 10968 21947 11020 21956
rect 10968 21913 10977 21947
rect 10977 21913 11011 21947
rect 11011 21913 11020 21947
rect 10968 21904 11020 21913
rect 11428 21904 11480 21956
rect 13544 21947 13596 21956
rect 13544 21913 13553 21947
rect 13553 21913 13587 21947
rect 13587 21913 13596 21947
rect 13544 21904 13596 21913
rect 15844 21904 15896 21956
rect 19340 21972 19392 22024
rect 22100 21972 22152 22024
rect 22468 21972 22520 22024
rect 22744 22015 22796 22024
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 23204 22015 23256 22024
rect 23204 21981 23213 22015
rect 23213 21981 23247 22015
rect 23247 21981 23256 22015
rect 23204 21972 23256 21981
rect 18604 21904 18656 21956
rect 18696 21947 18748 21956
rect 18696 21913 18705 21947
rect 18705 21913 18739 21947
rect 18739 21913 18748 21947
rect 18696 21904 18748 21913
rect 19432 21904 19484 21956
rect 19524 21947 19576 21956
rect 19524 21913 19533 21947
rect 19533 21913 19567 21947
rect 19567 21913 19576 21947
rect 19524 21904 19576 21913
rect 21180 21904 21232 21956
rect 23480 22049 23489 22083
rect 23489 22049 23523 22083
rect 23523 22049 23532 22083
rect 23480 22040 23532 22049
rect 24860 22040 24912 22092
rect 25136 22083 25188 22092
rect 25136 22049 25145 22083
rect 25145 22049 25179 22083
rect 25179 22049 25188 22083
rect 25136 22040 25188 22049
rect 11980 21836 12032 21888
rect 12256 21836 12308 21888
rect 16212 21836 16264 21888
rect 16672 21836 16724 21888
rect 16856 21879 16908 21888
rect 16856 21845 16865 21879
rect 16865 21845 16899 21879
rect 16899 21845 16908 21879
rect 16856 21836 16908 21845
rect 17040 21836 17092 21888
rect 17500 21836 17552 21888
rect 17684 21879 17736 21888
rect 17684 21845 17693 21879
rect 17693 21845 17727 21879
rect 17727 21845 17736 21879
rect 17684 21836 17736 21845
rect 17868 21836 17920 21888
rect 18236 21836 18288 21888
rect 18880 21879 18932 21888
rect 18880 21845 18889 21879
rect 18889 21845 18923 21879
rect 18923 21845 18932 21879
rect 18880 21836 18932 21845
rect 18972 21836 19024 21888
rect 20260 21836 20312 21888
rect 22008 21836 22060 21888
rect 24216 21836 24268 21888
rect 24584 21879 24636 21888
rect 24584 21845 24593 21879
rect 24593 21845 24627 21879
rect 24627 21845 24636 21879
rect 24584 21836 24636 21845
rect 24676 21836 24728 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 2228 21632 2280 21684
rect 9404 21632 9456 21684
rect 10048 21632 10100 21684
rect 13176 21632 13228 21684
rect 13360 21632 13412 21684
rect 17684 21632 17736 21684
rect 3424 21564 3476 21616
rect 4160 21496 4212 21548
rect 8484 21564 8536 21616
rect 16488 21564 16540 21616
rect 6736 21539 6788 21548
rect 6736 21505 6745 21539
rect 6745 21505 6779 21539
rect 6779 21505 6788 21539
rect 6736 21496 6788 21505
rect 7380 21539 7432 21548
rect 7380 21505 7389 21539
rect 7389 21505 7423 21539
rect 7423 21505 7432 21539
rect 7380 21496 7432 21505
rect 9036 21539 9088 21548
rect 9036 21505 9045 21539
rect 9045 21505 9079 21539
rect 9079 21505 9088 21539
rect 9036 21496 9088 21505
rect 10416 21496 10468 21548
rect 11428 21496 11480 21548
rect 12256 21496 12308 21548
rect 3516 21471 3568 21480
rect 3516 21437 3525 21471
rect 3525 21437 3559 21471
rect 3559 21437 3568 21471
rect 3516 21428 3568 21437
rect 5080 21471 5132 21480
rect 5080 21437 5089 21471
rect 5089 21437 5123 21471
rect 5123 21437 5132 21471
rect 5080 21428 5132 21437
rect 7288 21428 7340 21480
rect 9312 21471 9364 21480
rect 9312 21437 9321 21471
rect 9321 21437 9355 21471
rect 9355 21437 9364 21471
rect 9312 21428 9364 21437
rect 9404 21428 9456 21480
rect 10692 21428 10744 21480
rect 12624 21428 12676 21480
rect 13452 21428 13504 21480
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 15200 21496 15252 21548
rect 15936 21496 15988 21548
rect 15108 21428 15160 21480
rect 15476 21471 15528 21480
rect 15476 21437 15485 21471
rect 15485 21437 15519 21471
rect 15519 21437 15528 21471
rect 15476 21428 15528 21437
rect 15660 21471 15712 21480
rect 15660 21437 15669 21471
rect 15669 21437 15703 21471
rect 15703 21437 15712 21471
rect 15660 21428 15712 21437
rect 16304 21428 16356 21480
rect 19156 21564 19208 21616
rect 21088 21632 21140 21684
rect 17408 21539 17460 21548
rect 17408 21505 17417 21539
rect 17417 21505 17451 21539
rect 17451 21505 17460 21539
rect 17408 21496 17460 21505
rect 18880 21496 18932 21548
rect 19248 21496 19300 21548
rect 16948 21428 17000 21480
rect 6552 21335 6604 21344
rect 6552 21301 6561 21335
rect 6561 21301 6595 21335
rect 6595 21301 6604 21335
rect 6552 21292 6604 21301
rect 14464 21360 14516 21412
rect 17132 21360 17184 21412
rect 17316 21360 17368 21412
rect 10692 21292 10744 21344
rect 10784 21335 10836 21344
rect 10784 21301 10793 21335
rect 10793 21301 10827 21335
rect 10827 21301 10836 21335
rect 10784 21292 10836 21301
rect 10876 21292 10928 21344
rect 12808 21292 12860 21344
rect 16028 21292 16080 21344
rect 19708 21428 19760 21480
rect 20260 21496 20312 21548
rect 22744 21564 22796 21616
rect 21916 21496 21968 21548
rect 22192 21496 22244 21548
rect 23664 21564 23716 21616
rect 25228 21564 25280 21616
rect 21272 21428 21324 21480
rect 21456 21428 21508 21480
rect 23296 21496 23348 21548
rect 25136 21428 25188 21480
rect 18328 21360 18380 21412
rect 19340 21292 19392 21344
rect 19984 21292 20036 21344
rect 23756 21292 23808 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 3976 21088 4028 21140
rect 9220 21088 9272 21140
rect 10416 21088 10468 21140
rect 3424 21020 3476 21072
rect 2780 20995 2832 21004
rect 2780 20961 2789 20995
rect 2789 20961 2823 20995
rect 2823 20961 2832 20995
rect 2780 20952 2832 20961
rect 4252 20952 4304 21004
rect 7012 20952 7064 21004
rect 8484 21020 8536 21072
rect 10048 21020 10100 21072
rect 10508 20952 10560 21004
rect 10784 21020 10836 21072
rect 12440 21020 12492 21072
rect 13636 21088 13688 21140
rect 14464 21131 14516 21140
rect 14464 21097 14473 21131
rect 14473 21097 14507 21131
rect 14507 21097 14516 21131
rect 14464 21088 14516 21097
rect 11060 20952 11112 21004
rect 14740 20952 14792 21004
rect 17960 21088 18012 21140
rect 18512 21088 18564 21140
rect 18696 21088 18748 21140
rect 20444 21088 20496 21140
rect 21916 21088 21968 21140
rect 22652 21088 22704 21140
rect 22744 21088 22796 21140
rect 2228 20927 2280 20936
rect 2228 20893 2237 20927
rect 2237 20893 2271 20927
rect 2271 20893 2280 20927
rect 2228 20884 2280 20893
rect 5724 20884 5776 20936
rect 6276 20884 6328 20936
rect 6920 20927 6972 20936
rect 6920 20893 6929 20927
rect 6929 20893 6963 20927
rect 6963 20893 6972 20927
rect 6920 20884 6972 20893
rect 9312 20884 9364 20936
rect 12440 20884 12492 20936
rect 12992 20884 13044 20936
rect 6736 20816 6788 20868
rect 10968 20816 11020 20868
rect 11152 20816 11204 20868
rect 11428 20816 11480 20868
rect 13268 20816 13320 20868
rect 15476 20884 15528 20936
rect 14004 20816 14056 20868
rect 15844 20859 15896 20868
rect 15844 20825 15853 20859
rect 15853 20825 15887 20859
rect 15887 20825 15896 20859
rect 15844 20816 15896 20825
rect 15936 20816 15988 20868
rect 16488 20884 16540 20936
rect 17408 21020 17460 21072
rect 17684 21020 17736 21072
rect 22008 21020 22060 21072
rect 18328 20995 18380 21004
rect 18328 20961 18337 20995
rect 18337 20961 18371 20995
rect 18371 20961 18380 20995
rect 18328 20952 18380 20961
rect 18696 20952 18748 21004
rect 20904 20952 20956 21004
rect 21824 20952 21876 21004
rect 21916 20952 21968 21004
rect 25044 20952 25096 21004
rect 17684 20884 17736 20936
rect 5816 20791 5868 20800
rect 5816 20757 5825 20791
rect 5825 20757 5859 20791
rect 5859 20757 5868 20791
rect 5816 20748 5868 20757
rect 9312 20791 9364 20800
rect 9312 20757 9321 20791
rect 9321 20757 9355 20791
rect 9355 20757 9364 20791
rect 9312 20748 9364 20757
rect 10324 20791 10376 20800
rect 10324 20757 10333 20791
rect 10333 20757 10367 20791
rect 10367 20757 10376 20791
rect 10324 20748 10376 20757
rect 10416 20791 10468 20800
rect 10416 20757 10425 20791
rect 10425 20757 10459 20791
rect 10459 20757 10468 20791
rect 10416 20748 10468 20757
rect 10508 20748 10560 20800
rect 10876 20748 10928 20800
rect 13636 20748 13688 20800
rect 14096 20748 14148 20800
rect 15476 20748 15528 20800
rect 17040 20859 17092 20868
rect 17040 20825 17049 20859
rect 17049 20825 17083 20859
rect 17083 20825 17092 20859
rect 17040 20816 17092 20825
rect 19064 20816 19116 20868
rect 17408 20748 17460 20800
rect 17592 20748 17644 20800
rect 19340 20884 19392 20936
rect 23480 20884 23532 20936
rect 20260 20816 20312 20868
rect 20996 20816 21048 20868
rect 22652 20859 22704 20868
rect 22652 20825 22661 20859
rect 22661 20825 22695 20859
rect 22695 20825 22704 20859
rect 22652 20816 22704 20825
rect 23388 20816 23440 20868
rect 23664 20816 23716 20868
rect 23848 20816 23900 20868
rect 25228 20816 25280 20868
rect 21088 20748 21140 20800
rect 21640 20791 21692 20800
rect 21640 20757 21649 20791
rect 21649 20757 21683 20791
rect 21683 20757 21692 20791
rect 21640 20748 21692 20757
rect 22836 20791 22888 20800
rect 22836 20757 22845 20791
rect 22845 20757 22879 20791
rect 22879 20757 22888 20791
rect 22836 20748 22888 20757
rect 24584 20791 24636 20800
rect 24584 20757 24593 20791
rect 24593 20757 24627 20791
rect 24627 20757 24636 20791
rect 24584 20748 24636 20757
rect 24860 20748 24912 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 4988 20544 5040 20596
rect 5172 20587 5224 20596
rect 5172 20553 5181 20587
rect 5181 20553 5215 20587
rect 5215 20553 5224 20587
rect 5172 20544 5224 20553
rect 10324 20544 10376 20596
rect 10968 20544 11020 20596
rect 12440 20587 12492 20596
rect 12440 20553 12449 20587
rect 12449 20553 12483 20587
rect 12483 20553 12492 20587
rect 12440 20544 12492 20553
rect 12532 20587 12584 20596
rect 12532 20553 12541 20587
rect 12541 20553 12575 20587
rect 12575 20553 12584 20587
rect 12532 20544 12584 20553
rect 12716 20544 12768 20596
rect 17592 20544 17644 20596
rect 18696 20587 18748 20596
rect 18696 20553 18705 20587
rect 18705 20553 18739 20587
rect 18739 20553 18748 20587
rect 18696 20544 18748 20553
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 4712 20476 4764 20528
rect 5264 20476 5316 20528
rect 11428 20476 11480 20528
rect 12164 20476 12216 20528
rect 13544 20476 13596 20528
rect 18512 20476 18564 20528
rect 19156 20476 19208 20528
rect 20260 20544 20312 20596
rect 20812 20544 20864 20596
rect 23664 20544 23716 20596
rect 22192 20476 22244 20528
rect 22560 20476 22612 20528
rect 22744 20476 22796 20528
rect 23756 20519 23808 20528
rect 23756 20485 23765 20519
rect 23765 20485 23799 20519
rect 23799 20485 23808 20519
rect 23756 20476 23808 20485
rect 25228 20476 25280 20528
rect 5540 20408 5592 20460
rect 7196 20408 7248 20460
rect 7288 20451 7340 20460
rect 7288 20417 7297 20451
rect 7297 20417 7331 20451
rect 7331 20417 7340 20451
rect 7288 20408 7340 20417
rect 3332 20383 3384 20392
rect 3332 20349 3341 20383
rect 3341 20349 3375 20383
rect 3375 20349 3384 20383
rect 3332 20340 3384 20349
rect 9036 20451 9088 20460
rect 9036 20417 9045 20451
rect 9045 20417 9079 20451
rect 9079 20417 9088 20451
rect 9036 20408 9088 20417
rect 12808 20408 12860 20460
rect 8852 20272 8904 20324
rect 4068 20204 4120 20256
rect 4160 20204 4212 20256
rect 6092 20204 6144 20256
rect 8392 20247 8444 20256
rect 8392 20213 8401 20247
rect 8401 20213 8435 20247
rect 8435 20213 8444 20247
rect 8392 20204 8444 20213
rect 10048 20340 10100 20392
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 12440 20272 12492 20324
rect 15844 20451 15896 20460
rect 15844 20417 15853 20451
rect 15853 20417 15887 20451
rect 15887 20417 15896 20451
rect 15844 20408 15896 20417
rect 16488 20408 16540 20460
rect 23296 20408 23348 20460
rect 17684 20340 17736 20392
rect 19248 20383 19300 20392
rect 19248 20349 19257 20383
rect 19257 20349 19291 20383
rect 19291 20349 19300 20383
rect 19248 20340 19300 20349
rect 19892 20340 19944 20392
rect 21456 20340 21508 20392
rect 22376 20340 22428 20392
rect 22560 20383 22612 20392
rect 22560 20349 22569 20383
rect 22569 20349 22603 20383
rect 22603 20349 22612 20383
rect 22560 20340 22612 20349
rect 22652 20383 22704 20392
rect 22652 20349 22661 20383
rect 22661 20349 22695 20383
rect 22695 20349 22704 20383
rect 22652 20340 22704 20349
rect 16212 20272 16264 20324
rect 21548 20272 21600 20324
rect 22284 20272 22336 20324
rect 13820 20204 13872 20256
rect 14280 20204 14332 20256
rect 15108 20204 15160 20256
rect 15936 20247 15988 20256
rect 15936 20213 15945 20247
rect 15945 20213 15979 20247
rect 15979 20213 15988 20247
rect 15936 20204 15988 20213
rect 16028 20204 16080 20256
rect 16396 20204 16448 20256
rect 20812 20204 20864 20256
rect 21180 20204 21232 20256
rect 21824 20204 21876 20256
rect 23848 20340 23900 20392
rect 25228 20247 25280 20256
rect 25228 20213 25237 20247
rect 25237 20213 25271 20247
rect 25271 20213 25280 20247
rect 25228 20204 25280 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 1584 20000 1636 20052
rect 3976 20000 4028 20052
rect 6736 20000 6788 20052
rect 7196 20000 7248 20052
rect 5080 19932 5132 19984
rect 15292 20000 15344 20052
rect 16948 20000 17000 20052
rect 17592 20000 17644 20052
rect 19156 20000 19208 20052
rect 20260 20000 20312 20052
rect 21088 20000 21140 20052
rect 21916 20000 21968 20052
rect 24676 20000 24728 20052
rect 2044 19864 2096 19916
rect 2320 19796 2372 19848
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 5172 19839 5224 19848
rect 5172 19805 5181 19839
rect 5181 19805 5215 19839
rect 5215 19805 5224 19839
rect 5172 19796 5224 19805
rect 6736 19796 6788 19848
rect 9496 19796 9548 19848
rect 13452 19932 13504 19984
rect 13544 19932 13596 19984
rect 14096 19932 14148 19984
rect 14556 19932 14608 19984
rect 16396 19932 16448 19984
rect 18512 19932 18564 19984
rect 10968 19907 11020 19916
rect 10968 19873 10977 19907
rect 10977 19873 11011 19907
rect 11011 19873 11020 19907
rect 10968 19864 11020 19873
rect 11060 19864 11112 19916
rect 11244 19796 11296 19848
rect 11612 19839 11664 19848
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 7840 19728 7892 19780
rect 4528 19703 4580 19712
rect 4528 19669 4537 19703
rect 4537 19669 4571 19703
rect 4571 19669 4580 19703
rect 4528 19660 4580 19669
rect 5540 19660 5592 19712
rect 6644 19660 6696 19712
rect 8300 19660 8352 19712
rect 9128 19703 9180 19712
rect 9128 19669 9137 19703
rect 9137 19669 9171 19703
rect 9171 19669 9180 19703
rect 9128 19660 9180 19669
rect 10876 19660 10928 19712
rect 12164 19728 12216 19780
rect 13912 19796 13964 19848
rect 14188 19796 14240 19848
rect 13452 19728 13504 19780
rect 16948 19796 17000 19848
rect 18972 19932 19024 19984
rect 23572 19932 23624 19984
rect 18696 19864 18748 19916
rect 23296 19864 23348 19916
rect 24124 19864 24176 19916
rect 22928 19796 22980 19848
rect 15200 19728 15252 19780
rect 16212 19771 16264 19780
rect 16212 19737 16221 19771
rect 16221 19737 16255 19771
rect 16255 19737 16264 19771
rect 16212 19728 16264 19737
rect 16396 19728 16448 19780
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 16304 19703 16356 19712
rect 16304 19669 16313 19703
rect 16313 19669 16347 19703
rect 16347 19669 16356 19703
rect 16304 19660 16356 19669
rect 16580 19660 16632 19712
rect 20076 19728 20128 19780
rect 21364 19771 21416 19780
rect 21364 19737 21373 19771
rect 21373 19737 21407 19771
rect 21407 19737 21416 19771
rect 21364 19728 21416 19737
rect 21824 19728 21876 19780
rect 26056 19728 26108 19780
rect 19616 19660 19668 19712
rect 20812 19660 20864 19712
rect 23020 19660 23072 19712
rect 23112 19703 23164 19712
rect 23112 19669 23121 19703
rect 23121 19669 23155 19703
rect 23155 19669 23164 19703
rect 23112 19660 23164 19669
rect 23388 19660 23440 19712
rect 23480 19660 23532 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 5172 19456 5224 19508
rect 9220 19456 9272 19508
rect 3608 19320 3660 19372
rect 8208 19388 8260 19440
rect 10784 19456 10836 19508
rect 12164 19456 12216 19508
rect 5448 19320 5500 19372
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 1676 19252 1728 19304
rect 4528 19295 4580 19304
rect 4528 19261 4537 19295
rect 4537 19261 4571 19295
rect 4571 19261 4580 19295
rect 4528 19252 4580 19261
rect 6460 19295 6512 19304
rect 6460 19261 6469 19295
rect 6469 19261 6503 19295
rect 6503 19261 6512 19295
rect 6460 19252 6512 19261
rect 7564 19320 7616 19372
rect 7840 19320 7892 19372
rect 8300 19320 8352 19372
rect 7104 19252 7156 19304
rect 6920 19184 6972 19236
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 9036 19363 9088 19372
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 11612 19320 11664 19372
rect 13820 19456 13872 19508
rect 13912 19456 13964 19508
rect 14464 19499 14516 19508
rect 14464 19465 14473 19499
rect 14473 19465 14507 19499
rect 14507 19465 14516 19499
rect 14464 19456 14516 19465
rect 14832 19456 14884 19508
rect 16396 19456 16448 19508
rect 13544 19388 13596 19440
rect 14280 19388 14332 19440
rect 18696 19456 18748 19508
rect 14924 19320 14976 19372
rect 19892 19388 19944 19440
rect 20996 19388 21048 19440
rect 9404 19252 9456 19304
rect 11980 19252 12032 19304
rect 12072 19295 12124 19304
rect 12072 19261 12081 19295
rect 12081 19261 12115 19295
rect 12115 19261 12124 19295
rect 12072 19252 12124 19261
rect 15108 19252 15160 19304
rect 16028 19252 16080 19304
rect 16488 19320 16540 19372
rect 18328 19320 18380 19372
rect 19156 19320 19208 19372
rect 19708 19363 19760 19372
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 17316 19295 17368 19304
rect 17316 19261 17325 19295
rect 17325 19261 17359 19295
rect 17359 19261 17368 19295
rect 17316 19252 17368 19261
rect 2872 19116 2924 19168
rect 12164 19184 12216 19236
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 10968 19116 11020 19168
rect 11152 19116 11204 19168
rect 12256 19116 12308 19168
rect 13452 19116 13504 19168
rect 16304 19116 16356 19168
rect 16396 19116 16448 19168
rect 19708 19184 19760 19236
rect 19892 19295 19944 19304
rect 19892 19261 19901 19295
rect 19901 19261 19935 19295
rect 19935 19261 19944 19295
rect 19892 19252 19944 19261
rect 21824 19456 21876 19508
rect 22192 19456 22244 19508
rect 22468 19499 22520 19508
rect 22468 19465 22477 19499
rect 22477 19465 22511 19499
rect 22511 19465 22520 19499
rect 22468 19456 22520 19465
rect 23940 19456 23992 19508
rect 25044 19499 25096 19508
rect 25044 19465 25053 19499
rect 25053 19465 25087 19499
rect 25087 19465 25096 19499
rect 25044 19456 25096 19465
rect 21364 19388 21416 19440
rect 23848 19388 23900 19440
rect 22284 19320 22336 19372
rect 21548 19252 21600 19304
rect 22928 19320 22980 19372
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23296 19320 23348 19329
rect 21824 19184 21876 19236
rect 25228 19252 25280 19304
rect 25320 19295 25372 19304
rect 25320 19261 25329 19295
rect 25329 19261 25363 19295
rect 25363 19261 25372 19295
rect 25320 19252 25372 19261
rect 19156 19116 19208 19168
rect 21088 19116 21140 19168
rect 21732 19116 21784 19168
rect 23388 19116 23440 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 3700 18912 3752 18964
rect 4804 18912 4856 18964
rect 5908 18912 5960 18964
rect 8208 18912 8260 18964
rect 8852 18912 8904 18964
rect 9772 18912 9824 18964
rect 10324 18912 10376 18964
rect 11244 18912 11296 18964
rect 14280 18955 14332 18964
rect 14280 18921 14289 18955
rect 14289 18921 14323 18955
rect 14323 18921 14332 18955
rect 14280 18912 14332 18921
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 3700 18776 3752 18828
rect 4068 18844 4120 18896
rect 4160 18708 4212 18760
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 4804 18708 4856 18760
rect 5264 18640 5316 18692
rect 7472 18776 7524 18828
rect 8300 18776 8352 18828
rect 8760 18776 8812 18828
rect 6000 18751 6052 18760
rect 6000 18717 6009 18751
rect 6009 18717 6043 18751
rect 6043 18717 6052 18751
rect 6000 18708 6052 18717
rect 6460 18708 6512 18760
rect 8392 18708 8444 18760
rect 8576 18751 8628 18760
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 8576 18708 8628 18717
rect 9404 18776 9456 18828
rect 9496 18776 9548 18828
rect 11152 18844 11204 18896
rect 12348 18844 12400 18896
rect 13360 18776 13412 18828
rect 9128 18708 9180 18760
rect 8760 18640 8812 18692
rect 11980 18708 12032 18760
rect 12164 18708 12216 18760
rect 12440 18708 12492 18760
rect 12992 18640 13044 18692
rect 13728 18640 13780 18692
rect 4988 18572 5040 18624
rect 5172 18615 5224 18624
rect 5172 18581 5181 18615
rect 5181 18581 5215 18615
rect 5215 18581 5224 18615
rect 5172 18572 5224 18581
rect 6460 18615 6512 18624
rect 6460 18581 6469 18615
rect 6469 18581 6503 18615
rect 6503 18581 6512 18615
rect 6460 18572 6512 18581
rect 6644 18572 6696 18624
rect 9312 18572 9364 18624
rect 11704 18572 11756 18624
rect 11888 18615 11940 18624
rect 11888 18581 11897 18615
rect 11897 18581 11931 18615
rect 11931 18581 11940 18615
rect 11888 18572 11940 18581
rect 11980 18572 12032 18624
rect 14464 18572 14516 18624
rect 15476 18912 15528 18964
rect 15752 18912 15804 18964
rect 17224 18912 17276 18964
rect 17868 18912 17920 18964
rect 20720 18912 20772 18964
rect 21364 18912 21416 18964
rect 22836 18912 22888 18964
rect 23020 18912 23072 18964
rect 16856 18844 16908 18896
rect 17776 18844 17828 18896
rect 18052 18887 18104 18896
rect 18052 18853 18061 18887
rect 18061 18853 18095 18887
rect 18095 18853 18104 18887
rect 18052 18844 18104 18853
rect 18420 18844 18472 18896
rect 14924 18819 14976 18828
rect 14924 18785 14933 18819
rect 14933 18785 14967 18819
rect 14967 18785 14976 18819
rect 14924 18776 14976 18785
rect 15476 18819 15528 18828
rect 15476 18785 15485 18819
rect 15485 18785 15519 18819
rect 15519 18785 15528 18819
rect 15476 18776 15528 18785
rect 16488 18776 16540 18828
rect 17684 18776 17736 18828
rect 18328 18776 18380 18828
rect 15292 18640 15344 18692
rect 15200 18572 15252 18624
rect 17500 18708 17552 18760
rect 18512 18819 18564 18828
rect 18512 18785 18521 18819
rect 18521 18785 18555 18819
rect 18555 18785 18564 18819
rect 18512 18776 18564 18785
rect 22284 18844 22336 18896
rect 19064 18776 19116 18828
rect 21916 18776 21968 18828
rect 22836 18776 22888 18828
rect 25228 18819 25280 18828
rect 25228 18785 25237 18819
rect 25237 18785 25271 18819
rect 25271 18785 25280 18819
rect 25228 18776 25280 18785
rect 16028 18640 16080 18692
rect 16212 18640 16264 18692
rect 17132 18572 17184 18624
rect 17224 18572 17276 18624
rect 18236 18640 18288 18692
rect 19248 18708 19300 18760
rect 18512 18640 18564 18692
rect 19524 18640 19576 18692
rect 20260 18640 20312 18692
rect 20904 18640 20956 18692
rect 21088 18640 21140 18692
rect 21916 18640 21968 18692
rect 22928 18683 22980 18692
rect 22928 18649 22937 18683
rect 22937 18649 22971 18683
rect 22971 18649 22980 18683
rect 22928 18640 22980 18649
rect 23020 18683 23072 18692
rect 23020 18649 23029 18683
rect 23029 18649 23063 18683
rect 23063 18649 23072 18683
rect 23020 18640 23072 18649
rect 17684 18572 17736 18624
rect 17960 18572 18012 18624
rect 22008 18572 22060 18624
rect 22376 18572 22428 18624
rect 25228 18640 25280 18692
rect 24492 18572 24544 18624
rect 24860 18572 24912 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 2228 18411 2280 18420
rect 2228 18377 2237 18411
rect 2237 18377 2271 18411
rect 2271 18377 2280 18411
rect 2228 18368 2280 18377
rect 3792 18368 3844 18420
rect 4896 18368 4948 18420
rect 5724 18368 5776 18420
rect 6000 18368 6052 18420
rect 8576 18368 8628 18420
rect 12072 18368 12124 18420
rect 14464 18368 14516 18420
rect 15752 18368 15804 18420
rect 16488 18368 16540 18420
rect 19156 18368 19208 18420
rect 2872 18232 2924 18284
rect 4068 18232 4120 18284
rect 6092 18300 6144 18352
rect 10508 18300 10560 18352
rect 11336 18343 11388 18352
rect 11336 18309 11345 18343
rect 11345 18309 11379 18343
rect 11379 18309 11388 18343
rect 11336 18300 11388 18309
rect 5540 18232 5592 18284
rect 6920 18232 6972 18284
rect 7104 18232 7156 18284
rect 7656 18232 7708 18284
rect 8484 18275 8536 18284
rect 8484 18241 8493 18275
rect 8493 18241 8527 18275
rect 8527 18241 8536 18275
rect 8484 18232 8536 18241
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 10968 18232 11020 18284
rect 14372 18300 14424 18352
rect 14740 18343 14792 18352
rect 14740 18309 14749 18343
rect 14749 18309 14783 18343
rect 14783 18309 14792 18343
rect 14740 18300 14792 18309
rect 15476 18300 15528 18352
rect 16580 18300 16632 18352
rect 11980 18232 12032 18284
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 13360 18232 13412 18284
rect 15108 18232 15160 18284
rect 5632 18164 5684 18216
rect 7564 18164 7616 18216
rect 10784 18164 10836 18216
rect 8852 18096 8904 18148
rect 4068 18028 4120 18080
rect 7656 18071 7708 18080
rect 7656 18037 7665 18071
rect 7665 18037 7699 18071
rect 7699 18037 7708 18071
rect 7656 18028 7708 18037
rect 9772 18028 9824 18080
rect 12164 18164 12216 18216
rect 11704 18096 11756 18148
rect 16764 18232 16816 18284
rect 15936 18164 15988 18216
rect 16212 18164 16264 18216
rect 18512 18232 18564 18284
rect 19524 18232 19576 18284
rect 20260 18300 20312 18352
rect 20904 18343 20956 18352
rect 20904 18309 20913 18343
rect 20913 18309 20947 18343
rect 20947 18309 20956 18343
rect 20904 18300 20956 18309
rect 23112 18300 23164 18352
rect 17224 18096 17276 18148
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 16212 18028 16264 18037
rect 16488 18028 16540 18080
rect 17684 18164 17736 18216
rect 18696 18207 18748 18216
rect 18696 18173 18705 18207
rect 18705 18173 18739 18207
rect 18739 18173 18748 18207
rect 18696 18164 18748 18173
rect 19708 18207 19760 18216
rect 19708 18173 19717 18207
rect 19717 18173 19751 18207
rect 19751 18173 19760 18207
rect 19708 18164 19760 18173
rect 19156 18096 19208 18148
rect 19340 18096 19392 18148
rect 21364 18232 21416 18284
rect 21916 18232 21968 18284
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 23296 18411 23348 18420
rect 23296 18377 23305 18411
rect 23305 18377 23339 18411
rect 23339 18377 23348 18411
rect 23296 18368 23348 18377
rect 24952 18368 25004 18420
rect 23756 18232 23808 18284
rect 20720 18096 20772 18148
rect 20812 18096 20864 18148
rect 21088 18164 21140 18216
rect 24400 18207 24452 18216
rect 24400 18173 24409 18207
rect 24409 18173 24443 18207
rect 24443 18173 24452 18207
rect 24400 18164 24452 18173
rect 25504 18164 25556 18216
rect 17592 18028 17644 18080
rect 19892 18028 19944 18080
rect 20996 18028 21048 18080
rect 23480 18028 23532 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 4528 17824 4580 17876
rect 6368 17824 6420 17876
rect 7012 17824 7064 17876
rect 9128 17824 9180 17876
rect 11152 17824 11204 17876
rect 12072 17824 12124 17876
rect 12256 17824 12308 17876
rect 12440 17824 12492 17876
rect 13268 17824 13320 17876
rect 13820 17824 13872 17876
rect 16488 17824 16540 17876
rect 17132 17867 17184 17876
rect 17132 17833 17141 17867
rect 17141 17833 17175 17867
rect 17175 17833 17184 17867
rect 17132 17824 17184 17833
rect 17224 17824 17276 17876
rect 20628 17824 20680 17876
rect 22376 17824 22428 17876
rect 22652 17824 22704 17876
rect 6644 17756 6696 17808
rect 17316 17756 17368 17808
rect 6184 17688 6236 17740
rect 6552 17688 6604 17740
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 5816 17620 5868 17672
rect 7564 17620 7616 17672
rect 8944 17688 8996 17740
rect 11704 17688 11756 17740
rect 11888 17688 11940 17740
rect 12348 17688 12400 17740
rect 13452 17688 13504 17740
rect 13728 17688 13780 17740
rect 14740 17688 14792 17740
rect 14924 17731 14976 17740
rect 14924 17697 14933 17731
rect 14933 17697 14967 17731
rect 14967 17697 14976 17731
rect 14924 17688 14976 17697
rect 15200 17731 15252 17740
rect 15200 17697 15209 17731
rect 15209 17697 15243 17731
rect 15243 17697 15252 17731
rect 15200 17688 15252 17697
rect 15844 17688 15896 17740
rect 15936 17688 15988 17740
rect 9128 17620 9180 17672
rect 16580 17688 16632 17740
rect 4344 17552 4396 17604
rect 4528 17527 4580 17536
rect 4528 17493 4537 17527
rect 4537 17493 4571 17527
rect 4571 17493 4580 17527
rect 4528 17484 4580 17493
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7104 17484 7156 17493
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 17868 17620 17920 17672
rect 9496 17552 9548 17604
rect 10048 17595 10100 17604
rect 10048 17561 10057 17595
rect 10057 17561 10091 17595
rect 10091 17561 10100 17595
rect 10048 17552 10100 17561
rect 10140 17552 10192 17604
rect 10508 17552 10560 17604
rect 12992 17552 13044 17604
rect 14740 17552 14792 17604
rect 15660 17552 15712 17604
rect 19800 17688 19852 17740
rect 20260 17688 20312 17740
rect 11428 17484 11480 17536
rect 12256 17484 12308 17536
rect 14280 17484 14332 17536
rect 14464 17484 14516 17536
rect 17500 17527 17552 17536
rect 17500 17493 17509 17527
rect 17509 17493 17543 17527
rect 17543 17493 17552 17527
rect 17500 17484 17552 17493
rect 17684 17484 17736 17536
rect 18604 17527 18656 17536
rect 18604 17493 18613 17527
rect 18613 17493 18647 17527
rect 18647 17493 18656 17527
rect 18604 17484 18656 17493
rect 19708 17484 19760 17536
rect 20168 17484 20220 17536
rect 22192 17756 22244 17808
rect 23480 17756 23532 17808
rect 22560 17688 22612 17740
rect 23296 17688 23348 17740
rect 23848 17731 23900 17740
rect 23848 17697 23857 17731
rect 23857 17697 23891 17731
rect 23891 17697 23900 17731
rect 23848 17688 23900 17697
rect 24308 17688 24360 17740
rect 23204 17620 23256 17672
rect 24584 17620 24636 17672
rect 21088 17552 21140 17604
rect 21456 17552 21508 17604
rect 22744 17552 22796 17604
rect 23480 17552 23532 17604
rect 24492 17595 24544 17604
rect 24492 17561 24501 17595
rect 24501 17561 24535 17595
rect 24535 17561 24544 17595
rect 24492 17552 24544 17561
rect 25872 17552 25924 17604
rect 22284 17484 22336 17536
rect 22928 17527 22980 17536
rect 22928 17493 22937 17527
rect 22937 17493 22971 17527
rect 22971 17493 22980 17527
rect 22928 17484 22980 17493
rect 23572 17484 23624 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 3976 17280 4028 17332
rect 6552 17323 6604 17332
rect 6552 17289 6561 17323
rect 6561 17289 6595 17323
rect 6595 17289 6604 17323
rect 6552 17280 6604 17289
rect 7196 17323 7248 17332
rect 7196 17289 7205 17323
rect 7205 17289 7239 17323
rect 7239 17289 7248 17323
rect 7196 17280 7248 17289
rect 7380 17280 7432 17332
rect 8392 17280 8444 17332
rect 11888 17280 11940 17332
rect 12624 17280 12676 17332
rect 5540 17144 5592 17196
rect 8300 17212 8352 17264
rect 9772 17212 9824 17264
rect 10140 17212 10192 17264
rect 12072 17212 12124 17264
rect 13268 17212 13320 17264
rect 16396 17212 16448 17264
rect 6828 17144 6880 17196
rect 7472 17144 7524 17196
rect 7840 17076 7892 17128
rect 5080 17008 5132 17060
rect 8116 17076 8168 17128
rect 8944 17144 8996 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 9956 17076 10008 17128
rect 10048 17076 10100 17128
rect 8760 17008 8812 17060
rect 10048 16940 10100 16992
rect 10140 16940 10192 16992
rect 10600 16940 10652 16992
rect 12532 17076 12584 17128
rect 12992 17076 13044 17128
rect 14096 17144 14148 17196
rect 14740 17144 14792 17196
rect 13820 17076 13872 17128
rect 13452 17051 13504 17060
rect 13452 17017 13461 17051
rect 13461 17017 13495 17051
rect 13495 17017 13504 17051
rect 13452 17008 13504 17017
rect 13544 17008 13596 17060
rect 15200 17144 15252 17196
rect 15292 17076 15344 17128
rect 15936 17119 15988 17128
rect 15936 17085 15945 17119
rect 15945 17085 15979 17119
rect 15979 17085 15988 17119
rect 15936 17076 15988 17085
rect 16948 17144 17000 17196
rect 17684 17212 17736 17264
rect 20076 17280 20128 17332
rect 21088 17280 21140 17332
rect 21824 17280 21876 17332
rect 22100 17212 22152 17264
rect 18328 17187 18380 17196
rect 18328 17153 18337 17187
rect 18337 17153 18371 17187
rect 18371 17153 18380 17187
rect 18328 17144 18380 17153
rect 17224 17008 17276 17060
rect 19248 17076 19300 17128
rect 18328 17008 18380 17060
rect 19708 17008 19760 17060
rect 21088 17144 21140 17196
rect 22744 17280 22796 17332
rect 24308 17323 24360 17332
rect 24308 17289 24317 17323
rect 24317 17289 24351 17323
rect 24351 17289 24360 17323
rect 24308 17280 24360 17289
rect 22928 17212 22980 17264
rect 22560 17187 22612 17196
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 24860 17187 24912 17196
rect 24860 17153 24869 17187
rect 24869 17153 24903 17187
rect 24903 17153 24912 17187
rect 24860 17144 24912 17153
rect 25044 17144 25096 17196
rect 20076 17119 20128 17128
rect 20076 17085 20085 17119
rect 20085 17085 20119 17119
rect 20119 17085 20128 17119
rect 20076 17076 20128 17085
rect 21272 17076 21324 17128
rect 21456 17076 21508 17128
rect 11980 16940 12032 16992
rect 14464 16940 14516 16992
rect 14740 16940 14792 16992
rect 16856 16983 16908 16992
rect 16856 16949 16865 16983
rect 16865 16949 16899 16983
rect 16899 16949 16908 16983
rect 16856 16940 16908 16949
rect 18144 16940 18196 16992
rect 22192 17008 22244 17060
rect 20628 16940 20680 16992
rect 22376 17008 22428 17060
rect 22560 17008 22612 17060
rect 25688 17008 25740 17060
rect 22928 16940 22980 16992
rect 23848 16940 23900 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 6828 16779 6880 16788
rect 6828 16745 6837 16779
rect 6837 16745 6871 16779
rect 6871 16745 6880 16779
rect 6828 16736 6880 16745
rect 7472 16736 7524 16788
rect 9312 16668 9364 16720
rect 9680 16736 9732 16788
rect 11244 16736 11296 16788
rect 14740 16736 14792 16788
rect 16028 16779 16080 16788
rect 16028 16745 16037 16779
rect 16037 16745 16071 16779
rect 16071 16745 16080 16779
rect 16028 16736 16080 16745
rect 16672 16736 16724 16788
rect 5264 16643 5316 16652
rect 5264 16609 5273 16643
rect 5273 16609 5307 16643
rect 5307 16609 5316 16643
rect 5264 16600 5316 16609
rect 8668 16600 8720 16652
rect 9588 16600 9640 16652
rect 8576 16571 8628 16584
rect 8576 16537 8585 16571
rect 8585 16537 8619 16571
rect 8619 16537 8628 16571
rect 10140 16668 10192 16720
rect 11980 16668 12032 16720
rect 13268 16668 13320 16720
rect 13912 16668 13964 16720
rect 11336 16600 11388 16652
rect 11612 16600 11664 16652
rect 13728 16600 13780 16652
rect 14924 16600 14976 16652
rect 8576 16532 8628 16537
rect 10876 16532 10928 16584
rect 11244 16575 11296 16584
rect 11244 16541 11253 16575
rect 11253 16541 11287 16575
rect 11287 16541 11296 16575
rect 11244 16532 11296 16541
rect 11704 16532 11756 16584
rect 12532 16464 12584 16516
rect 14832 16464 14884 16516
rect 15016 16464 15068 16516
rect 17132 16575 17184 16584
rect 17132 16541 17141 16575
rect 17141 16541 17175 16575
rect 17175 16541 17184 16575
rect 17132 16532 17184 16541
rect 17408 16464 17460 16516
rect 17684 16464 17736 16516
rect 22192 16736 22244 16788
rect 23296 16736 23348 16788
rect 22284 16643 22336 16652
rect 22284 16609 22293 16643
rect 22293 16609 22327 16643
rect 22327 16609 22336 16643
rect 22284 16600 22336 16609
rect 22652 16600 22704 16652
rect 25596 16600 25648 16652
rect 19432 16464 19484 16516
rect 19708 16507 19760 16516
rect 19708 16473 19717 16507
rect 19717 16473 19751 16507
rect 19751 16473 19760 16507
rect 19708 16464 19760 16473
rect 20168 16464 20220 16516
rect 23848 16464 23900 16516
rect 23940 16464 23992 16516
rect 4712 16439 4764 16448
rect 4712 16405 4721 16439
rect 4721 16405 4755 16439
rect 4755 16405 4764 16439
rect 4712 16396 4764 16405
rect 9772 16396 9824 16448
rect 9864 16396 9916 16448
rect 10140 16439 10192 16448
rect 10140 16405 10149 16439
rect 10149 16405 10183 16439
rect 10183 16405 10192 16439
rect 10140 16396 10192 16405
rect 10784 16439 10836 16448
rect 10784 16405 10793 16439
rect 10793 16405 10827 16439
rect 10827 16405 10836 16439
rect 10784 16396 10836 16405
rect 11152 16396 11204 16448
rect 11796 16396 11848 16448
rect 11980 16396 12032 16448
rect 12164 16396 12216 16448
rect 17224 16396 17276 16448
rect 19248 16396 19300 16448
rect 21272 16396 21324 16448
rect 21640 16439 21692 16448
rect 21640 16405 21649 16439
rect 21649 16405 21683 16439
rect 21683 16405 21692 16439
rect 21640 16396 21692 16405
rect 23296 16396 23348 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 7840 16192 7892 16244
rect 8208 16192 8260 16244
rect 4712 16124 4764 16176
rect 9496 16124 9548 16176
rect 10140 16192 10192 16244
rect 7748 16056 7800 16108
rect 8208 16056 8260 16108
rect 8668 16099 8720 16108
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 9588 16056 9640 16108
rect 9864 16056 9916 16108
rect 10692 16124 10744 16176
rect 11888 16124 11940 16176
rect 11980 16167 12032 16176
rect 11980 16133 11989 16167
rect 11989 16133 12023 16167
rect 12023 16133 12032 16167
rect 11980 16124 12032 16133
rect 12532 16124 12584 16176
rect 7288 15988 7340 16040
rect 6276 15920 6328 15972
rect 8484 15895 8536 15904
rect 8484 15861 8493 15895
rect 8493 15861 8527 15895
rect 8527 15861 8536 15895
rect 8484 15852 8536 15861
rect 9128 15963 9180 15972
rect 9128 15929 9137 15963
rect 9137 15929 9171 15963
rect 9171 15929 9180 15963
rect 9128 15920 9180 15929
rect 10324 15920 10376 15972
rect 10968 15988 11020 16040
rect 10784 15852 10836 15904
rect 11704 16031 11756 16040
rect 11704 15997 11713 16031
rect 11713 15997 11747 16031
rect 11747 15997 11756 16031
rect 11704 15988 11756 15997
rect 12348 15988 12400 16040
rect 12716 15988 12768 16040
rect 13452 16031 13504 16040
rect 13452 15997 13461 16031
rect 13461 15997 13495 16031
rect 13495 15997 13504 16031
rect 13452 15988 13504 15997
rect 19432 16192 19484 16244
rect 20076 16192 20128 16244
rect 20444 16192 20496 16244
rect 23664 16192 23716 16244
rect 15752 16124 15804 16176
rect 19156 16124 19208 16176
rect 20904 16167 20956 16176
rect 20904 16133 20913 16167
rect 20913 16133 20947 16167
rect 20947 16133 20956 16167
rect 20904 16124 20956 16133
rect 24032 16124 24084 16176
rect 24676 16167 24728 16176
rect 24676 16133 24685 16167
rect 24685 16133 24719 16167
rect 24719 16133 24728 16167
rect 24676 16124 24728 16133
rect 14004 16056 14056 16108
rect 16212 16056 16264 16108
rect 19064 16056 19116 16108
rect 19708 16099 19760 16108
rect 19708 16065 19717 16099
rect 19717 16065 19751 16099
rect 19751 16065 19760 16099
rect 19708 16056 19760 16065
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 15200 15988 15252 16040
rect 18972 15988 19024 16040
rect 20168 16056 20220 16108
rect 21456 16056 21508 16108
rect 24584 16056 24636 16108
rect 17500 15920 17552 15972
rect 21088 16031 21140 16040
rect 21088 15997 21097 16031
rect 21097 15997 21131 16031
rect 21131 15997 21140 16031
rect 21088 15988 21140 15997
rect 21732 15988 21784 16040
rect 22560 16031 22612 16040
rect 22560 15997 22569 16031
rect 22569 15997 22603 16031
rect 22603 15997 22612 16031
rect 22560 15988 22612 15997
rect 20076 15920 20128 15972
rect 22744 15920 22796 15972
rect 23296 15920 23348 15972
rect 25044 15920 25096 15972
rect 12072 15852 12124 15904
rect 13912 15895 13964 15904
rect 13912 15861 13921 15895
rect 13921 15861 13955 15895
rect 13955 15861 13964 15895
rect 13912 15852 13964 15861
rect 15016 15895 15068 15904
rect 15016 15861 15025 15895
rect 15025 15861 15059 15895
rect 15059 15861 15068 15895
rect 15016 15852 15068 15861
rect 16304 15852 16356 15904
rect 17868 15852 17920 15904
rect 18880 15852 18932 15904
rect 20536 15895 20588 15904
rect 20536 15861 20545 15895
rect 20545 15861 20579 15895
rect 20579 15861 20588 15895
rect 20536 15852 20588 15861
rect 22376 15852 22428 15904
rect 22560 15852 22612 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 8760 15691 8812 15700
rect 8760 15657 8769 15691
rect 8769 15657 8803 15691
rect 8803 15657 8812 15691
rect 8760 15648 8812 15657
rect 11888 15648 11940 15700
rect 13912 15648 13964 15700
rect 16856 15648 16908 15700
rect 12716 15512 12768 15564
rect 9496 15444 9548 15496
rect 9956 15444 10008 15496
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 10692 15376 10744 15428
rect 12532 15376 12584 15428
rect 15844 15580 15896 15632
rect 16304 15623 16356 15632
rect 16304 15589 16313 15623
rect 16313 15589 16347 15623
rect 16347 15589 16356 15623
rect 16304 15580 16356 15589
rect 16764 15580 16816 15632
rect 19340 15648 19392 15700
rect 20536 15648 20588 15700
rect 25412 15648 25464 15700
rect 18604 15580 18656 15632
rect 14188 15512 14240 15564
rect 14280 15555 14332 15564
rect 14280 15521 14289 15555
rect 14289 15521 14323 15555
rect 14323 15521 14332 15555
rect 14280 15512 14332 15521
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 21180 15555 21232 15564
rect 21180 15521 21189 15555
rect 21189 15521 21223 15555
rect 21223 15521 21232 15555
rect 21180 15512 21232 15521
rect 21272 15555 21324 15564
rect 21272 15521 21281 15555
rect 21281 15521 21315 15555
rect 21315 15521 21324 15555
rect 21272 15512 21324 15521
rect 13820 15444 13872 15496
rect 19984 15487 20036 15496
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 25780 15512 25832 15564
rect 14464 15376 14516 15428
rect 11152 15308 11204 15360
rect 11612 15308 11664 15360
rect 12348 15308 12400 15360
rect 13912 15308 13964 15360
rect 15016 15376 15068 15428
rect 16580 15376 16632 15428
rect 17316 15376 17368 15428
rect 17224 15308 17276 15360
rect 17684 15376 17736 15428
rect 21640 15376 21692 15428
rect 18972 15351 19024 15360
rect 18972 15317 18981 15351
rect 18981 15317 19015 15351
rect 19015 15317 19024 15351
rect 18972 15308 19024 15317
rect 20536 15308 20588 15360
rect 21364 15308 21416 15360
rect 23756 15444 23808 15496
rect 22744 15419 22796 15428
rect 22744 15385 22753 15419
rect 22753 15385 22787 15419
rect 22787 15385 22796 15419
rect 22744 15376 22796 15385
rect 22836 15351 22888 15360
rect 22836 15317 22845 15351
rect 22845 15317 22879 15351
rect 22879 15317 22888 15351
rect 22836 15308 22888 15317
rect 23480 15308 23532 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 4068 15104 4120 15156
rect 5540 15104 5592 15156
rect 9496 15147 9548 15156
rect 9496 15113 9505 15147
rect 9505 15113 9539 15147
rect 9539 15113 9548 15147
rect 9496 15104 9548 15113
rect 10048 15104 10100 15156
rect 14924 15104 14976 15156
rect 12532 15036 12584 15088
rect 14004 15036 14056 15088
rect 10508 15011 10560 15020
rect 10508 14977 10517 15011
rect 10517 14977 10551 15011
rect 10551 14977 10560 15011
rect 10508 14968 10560 14977
rect 11152 15011 11204 15020
rect 11152 14977 11161 15011
rect 11161 14977 11195 15011
rect 11195 14977 11204 15011
rect 11152 14968 11204 14977
rect 13820 14968 13872 15020
rect 15108 14968 15160 15020
rect 15384 15036 15436 15088
rect 18880 15104 18932 15156
rect 19156 15104 19208 15156
rect 22468 15104 22520 15156
rect 16764 15036 16816 15088
rect 17224 15036 17276 15088
rect 18972 15036 19024 15088
rect 21456 15079 21508 15088
rect 21456 15045 21465 15079
rect 21465 15045 21499 15079
rect 21499 15045 21508 15079
rect 21456 15036 21508 15045
rect 22100 15079 22152 15088
rect 22100 15045 22109 15079
rect 22109 15045 22143 15079
rect 22143 15045 22152 15079
rect 22100 15036 22152 15045
rect 23296 15104 23348 15156
rect 24124 15104 24176 15156
rect 23664 15036 23716 15088
rect 16488 14968 16540 15020
rect 10600 14900 10652 14952
rect 10692 14900 10744 14952
rect 11704 14943 11756 14952
rect 11704 14909 11713 14943
rect 11713 14909 11747 14943
rect 11747 14909 11756 14943
rect 11704 14900 11756 14909
rect 11980 14943 12032 14952
rect 11980 14909 11989 14943
rect 11989 14909 12023 14943
rect 12023 14909 12032 14943
rect 11980 14900 12032 14909
rect 12072 14900 12124 14952
rect 13636 14832 13688 14884
rect 16672 14832 16724 14884
rect 13452 14764 13504 14816
rect 14832 14807 14884 14816
rect 14832 14773 14841 14807
rect 14841 14773 14875 14807
rect 14875 14773 14884 14807
rect 14832 14764 14884 14773
rect 16488 14764 16540 14816
rect 17132 14900 17184 14952
rect 19340 14943 19392 14952
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 18972 14832 19024 14884
rect 18604 14807 18656 14816
rect 18604 14773 18613 14807
rect 18613 14773 18647 14807
rect 18647 14773 18656 14807
rect 18604 14764 18656 14773
rect 19064 14807 19116 14816
rect 19064 14773 19073 14807
rect 19073 14773 19107 14807
rect 19107 14773 19116 14807
rect 19064 14764 19116 14773
rect 20720 14832 20772 14884
rect 22192 14968 22244 15020
rect 21824 14900 21876 14952
rect 22284 14900 22336 14952
rect 21180 14832 21232 14884
rect 22652 14764 22704 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 10508 14560 10560 14612
rect 11152 14560 11204 14612
rect 13636 14560 13688 14612
rect 13820 14492 13872 14544
rect 11612 14424 11664 14476
rect 11980 14424 12032 14476
rect 14648 14560 14700 14612
rect 14924 14560 14976 14612
rect 18972 14560 19024 14612
rect 19248 14560 19300 14612
rect 19616 14560 19668 14612
rect 20352 14560 20404 14612
rect 21456 14560 21508 14612
rect 22284 14603 22336 14612
rect 22284 14569 22293 14603
rect 22293 14569 22327 14603
rect 22327 14569 22336 14603
rect 22284 14560 22336 14569
rect 22468 14560 22520 14612
rect 24952 14560 25004 14612
rect 25136 14560 25188 14612
rect 26148 14560 26200 14612
rect 18696 14492 18748 14544
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 14280 14467 14332 14476
rect 14280 14433 14289 14467
rect 14289 14433 14323 14467
rect 14323 14433 14332 14467
rect 14280 14424 14332 14433
rect 14556 14467 14608 14476
rect 14556 14433 14565 14467
rect 14565 14433 14599 14467
rect 14599 14433 14608 14467
rect 14556 14424 14608 14433
rect 16488 14467 16540 14476
rect 16488 14433 16497 14467
rect 16497 14433 16531 14467
rect 16531 14433 16540 14467
rect 16488 14424 16540 14433
rect 18604 14424 18656 14476
rect 20904 14492 20956 14544
rect 23664 14492 23716 14544
rect 23388 14424 23440 14476
rect 24492 14424 24544 14476
rect 13912 14356 13964 14408
rect 19156 14356 19208 14408
rect 22008 14356 22060 14408
rect 24860 14356 24912 14408
rect 12532 14220 12584 14272
rect 15016 14288 15068 14340
rect 17224 14288 17276 14340
rect 19616 14288 19668 14340
rect 19892 14331 19944 14340
rect 19892 14297 19901 14331
rect 19901 14297 19935 14331
rect 19935 14297 19944 14331
rect 19892 14288 19944 14297
rect 19984 14288 20036 14340
rect 15200 14220 15252 14272
rect 16580 14220 16632 14272
rect 18880 14220 18932 14272
rect 19156 14220 19208 14272
rect 22744 14220 22796 14272
rect 24308 14288 24360 14340
rect 24124 14220 24176 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 11520 13948 11572 14000
rect 13728 14016 13780 14068
rect 13820 14016 13872 14068
rect 14372 14016 14424 14068
rect 14648 14016 14700 14068
rect 16120 14059 16172 14068
rect 16120 14025 16129 14059
rect 16129 14025 16163 14059
rect 16163 14025 16172 14059
rect 16120 14016 16172 14025
rect 17132 14016 17184 14068
rect 17592 14016 17644 14068
rect 19340 14016 19392 14068
rect 20352 14059 20404 14068
rect 20352 14025 20361 14059
rect 20361 14025 20395 14059
rect 20395 14025 20404 14059
rect 20352 14016 20404 14025
rect 20628 14016 20680 14068
rect 21180 14016 21232 14068
rect 11888 13812 11940 13864
rect 13452 13812 13504 13864
rect 14280 13948 14332 14000
rect 15108 13880 15160 13932
rect 15476 13812 15528 13864
rect 17408 13923 17460 13932
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 17684 13948 17736 14000
rect 17868 13948 17920 14000
rect 19064 13948 19116 14000
rect 19432 13948 19484 14000
rect 21916 13948 21968 14000
rect 24032 14016 24084 14068
rect 23664 13948 23716 14000
rect 25136 13991 25188 14000
rect 25136 13957 25145 13991
rect 25145 13957 25179 13991
rect 25179 13957 25188 13991
rect 25136 13948 25188 13957
rect 20720 13880 20772 13932
rect 13728 13744 13780 13796
rect 17592 13744 17644 13796
rect 20996 13812 21048 13864
rect 22100 13923 22152 13932
rect 22100 13889 22109 13923
rect 22109 13889 22143 13923
rect 22143 13889 22152 13923
rect 22100 13880 22152 13889
rect 22284 13880 22336 13932
rect 21456 13812 21508 13864
rect 21824 13812 21876 13864
rect 24492 13812 24544 13864
rect 25320 13855 25372 13864
rect 25320 13821 25329 13855
rect 25329 13821 25363 13855
rect 25363 13821 25372 13855
rect 25320 13812 25372 13821
rect 16028 13676 16080 13728
rect 17316 13676 17368 13728
rect 18512 13676 18564 13728
rect 20720 13719 20772 13728
rect 20720 13685 20729 13719
rect 20729 13685 20763 13719
rect 20763 13685 20772 13719
rect 20720 13676 20772 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 12532 13472 12584 13524
rect 13728 13472 13780 13524
rect 16028 13515 16080 13524
rect 16028 13481 16037 13515
rect 16037 13481 16071 13515
rect 16071 13481 16080 13515
rect 16028 13472 16080 13481
rect 17500 13472 17552 13524
rect 19708 13472 19760 13524
rect 20628 13472 20680 13524
rect 21180 13472 21232 13524
rect 21456 13515 21508 13524
rect 21456 13481 21465 13515
rect 21465 13481 21499 13515
rect 21499 13481 21508 13515
rect 21456 13472 21508 13481
rect 21732 13472 21784 13524
rect 13452 13404 13504 13456
rect 12716 13336 12768 13388
rect 13360 13336 13412 13388
rect 14280 13379 14332 13388
rect 14280 13345 14289 13379
rect 14289 13345 14323 13379
rect 14323 13345 14332 13379
rect 14280 13336 14332 13345
rect 17868 13404 17920 13456
rect 19156 13404 19208 13456
rect 19432 13404 19484 13456
rect 23664 13404 23716 13456
rect 16396 13336 16448 13388
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 18696 13336 18748 13388
rect 21916 13379 21968 13388
rect 10048 13132 10100 13184
rect 10692 13132 10744 13184
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 19432 13268 19484 13320
rect 21916 13345 21925 13379
rect 21925 13345 21959 13379
rect 21959 13345 21968 13379
rect 21916 13336 21968 13345
rect 22284 13336 22336 13388
rect 22744 13336 22796 13388
rect 22928 13336 22980 13388
rect 23756 13336 23808 13388
rect 25228 13336 25280 13388
rect 12072 13243 12124 13252
rect 12072 13209 12081 13243
rect 12081 13209 12115 13243
rect 12115 13209 12124 13243
rect 12072 13200 12124 13209
rect 12532 13200 12584 13252
rect 14188 13200 14240 13252
rect 14556 13243 14608 13252
rect 14556 13209 14565 13243
rect 14565 13209 14599 13243
rect 14599 13209 14608 13243
rect 14556 13200 14608 13209
rect 13728 13132 13780 13184
rect 15016 13200 15068 13252
rect 17224 13200 17276 13252
rect 16120 13132 16172 13184
rect 17592 13132 17644 13184
rect 19064 13132 19116 13184
rect 19524 13132 19576 13184
rect 20628 13200 20680 13252
rect 22468 13200 22520 13252
rect 22744 13200 22796 13252
rect 25228 13200 25280 13252
rect 20812 13132 20864 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 12532 12971 12584 12980
rect 12532 12937 12541 12971
rect 12541 12937 12575 12971
rect 12575 12937 12584 12971
rect 12532 12928 12584 12937
rect 14280 12971 14332 12980
rect 14280 12937 14289 12971
rect 14289 12937 14323 12971
rect 14323 12937 14332 12971
rect 14280 12928 14332 12937
rect 22100 12928 22152 12980
rect 22468 12928 22520 12980
rect 23756 12971 23808 12980
rect 23756 12937 23765 12971
rect 23765 12937 23799 12971
rect 23799 12937 23808 12971
rect 23756 12928 23808 12937
rect 24860 12971 24912 12980
rect 24860 12937 24869 12971
rect 24869 12937 24903 12971
rect 24903 12937 24912 12971
rect 24860 12928 24912 12937
rect 12716 12860 12768 12912
rect 15016 12860 15068 12912
rect 16304 12903 16356 12912
rect 16304 12869 16313 12903
rect 16313 12869 16347 12903
rect 16347 12869 16356 12903
rect 16304 12860 16356 12869
rect 17224 12860 17276 12912
rect 17592 12860 17644 12912
rect 18880 12860 18932 12912
rect 21548 12903 21600 12912
rect 21548 12869 21557 12903
rect 21557 12869 21591 12903
rect 21591 12869 21600 12903
rect 21548 12860 21600 12869
rect 16580 12792 16632 12844
rect 18420 12792 18472 12844
rect 21640 12792 21692 12844
rect 13360 12724 13412 12776
rect 14280 12724 14332 12776
rect 15476 12724 15528 12776
rect 17500 12724 17552 12776
rect 18328 12724 18380 12776
rect 18696 12724 18748 12776
rect 19156 12724 19208 12776
rect 19524 12767 19576 12776
rect 19524 12733 19533 12767
rect 19533 12733 19567 12767
rect 19567 12733 19576 12767
rect 19524 12724 19576 12733
rect 18604 12699 18656 12708
rect 18604 12665 18613 12699
rect 18613 12665 18647 12699
rect 18647 12665 18656 12699
rect 19800 12724 19852 12776
rect 18604 12656 18656 12665
rect 19064 12631 19116 12640
rect 19064 12597 19073 12631
rect 19073 12597 19107 12631
rect 19107 12597 19116 12631
rect 19064 12588 19116 12597
rect 19156 12588 19208 12640
rect 20260 12631 20312 12640
rect 20260 12597 20269 12631
rect 20269 12597 20303 12631
rect 20303 12597 20312 12631
rect 20260 12588 20312 12597
rect 20628 12656 20680 12708
rect 21180 12724 21232 12776
rect 22284 12860 22336 12912
rect 21916 12792 21968 12844
rect 24768 12792 24820 12844
rect 22284 12767 22336 12776
rect 22284 12733 22293 12767
rect 22293 12733 22327 12767
rect 22327 12733 22336 12767
rect 22284 12724 22336 12733
rect 22744 12724 22796 12776
rect 24216 12699 24268 12708
rect 24216 12665 24225 12699
rect 24225 12665 24259 12699
rect 24259 12665 24268 12699
rect 24216 12656 24268 12665
rect 23388 12588 23440 12640
rect 25136 12588 25188 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 13728 12427 13780 12436
rect 13728 12393 13737 12427
rect 13737 12393 13771 12427
rect 13771 12393 13780 12427
rect 13728 12384 13780 12393
rect 13912 12427 13964 12436
rect 13912 12393 13921 12427
rect 13921 12393 13955 12427
rect 13955 12393 13964 12427
rect 13912 12384 13964 12393
rect 15016 12384 15068 12436
rect 16396 12384 16448 12436
rect 17500 12427 17552 12436
rect 17500 12393 17509 12427
rect 17509 12393 17543 12427
rect 17543 12393 17552 12427
rect 17500 12384 17552 12393
rect 18788 12384 18840 12436
rect 19892 12384 19944 12436
rect 22008 12384 22060 12436
rect 22284 12384 22336 12436
rect 24860 12384 24912 12436
rect 4988 12248 5040 12300
rect 15476 12248 15528 12300
rect 17408 12248 17460 12300
rect 18880 12291 18932 12300
rect 18880 12257 18889 12291
rect 18889 12257 18923 12291
rect 18923 12257 18932 12291
rect 18880 12248 18932 12257
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 20352 12248 20404 12300
rect 21364 12248 21416 12300
rect 21916 12248 21968 12300
rect 24492 12248 24544 12300
rect 24584 12291 24636 12300
rect 24584 12257 24593 12291
rect 24593 12257 24627 12291
rect 24627 12257 24636 12291
rect 24584 12248 24636 12257
rect 15568 12180 15620 12232
rect 19340 12180 19392 12232
rect 21640 12223 21692 12232
rect 21640 12189 21649 12223
rect 21649 12189 21683 12223
rect 21683 12189 21692 12223
rect 21640 12180 21692 12189
rect 16120 12112 16172 12164
rect 16304 12112 16356 12164
rect 18696 12155 18748 12164
rect 18696 12121 18705 12155
rect 18705 12121 18739 12155
rect 18739 12121 18748 12155
rect 18696 12112 18748 12121
rect 17592 12044 17644 12096
rect 19248 12112 19300 12164
rect 21548 12112 21600 12164
rect 18880 12044 18932 12096
rect 19524 12044 19576 12096
rect 19800 12044 19852 12096
rect 20628 12044 20680 12096
rect 25136 12044 25188 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 15108 11883 15160 11892
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 15660 11883 15712 11892
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 13360 11772 13412 11824
rect 13728 11772 13780 11824
rect 19340 11840 19392 11892
rect 17500 11772 17552 11824
rect 18880 11772 18932 11824
rect 21272 11840 21324 11892
rect 19800 11772 19852 11824
rect 20996 11772 21048 11824
rect 25504 11840 25556 11892
rect 24860 11772 24912 11824
rect 13452 11636 13504 11688
rect 14096 11568 14148 11620
rect 19432 11747 19484 11756
rect 19432 11713 19441 11747
rect 19441 11713 19475 11747
rect 19475 11713 19484 11747
rect 19432 11704 19484 11713
rect 21180 11704 21232 11756
rect 21548 11704 21600 11756
rect 18604 11636 18656 11688
rect 19340 11636 19392 11688
rect 21088 11568 21140 11620
rect 21640 11568 21692 11620
rect 18788 11500 18840 11552
rect 19708 11500 19760 11552
rect 19800 11500 19852 11552
rect 20996 11500 21048 11552
rect 22008 11636 22060 11688
rect 23940 11747 23992 11756
rect 23940 11713 23949 11747
rect 23949 11713 23983 11747
rect 23983 11713 23992 11747
rect 23940 11704 23992 11713
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 26056 11500 26108 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 15016 11296 15068 11348
rect 16120 11271 16172 11280
rect 16120 11237 16129 11271
rect 16129 11237 16163 11271
rect 16163 11237 16172 11271
rect 16120 11228 16172 11237
rect 16948 11296 17000 11348
rect 17316 11296 17368 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 19800 11296 19852 11348
rect 20812 11296 20864 11348
rect 19248 11228 19300 11280
rect 19616 11228 19668 11280
rect 20996 11228 21048 11280
rect 25044 11228 25096 11280
rect 17868 11160 17920 11212
rect 18420 11160 18472 11212
rect 15752 11092 15804 11144
rect 16396 11092 16448 11144
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 21732 11160 21784 11212
rect 24860 11160 24912 11212
rect 20444 11135 20496 11144
rect 20444 11101 20453 11135
rect 20453 11101 20487 11135
rect 20487 11101 20496 11135
rect 20444 11092 20496 11101
rect 20904 11092 20956 11144
rect 21548 11092 21600 11144
rect 22376 11092 22428 11144
rect 22652 11135 22704 11144
rect 22652 11101 22661 11135
rect 22661 11101 22695 11135
rect 22695 11101 22704 11135
rect 22652 11092 22704 11101
rect 24400 11092 24452 11144
rect 19708 11067 19760 11076
rect 19708 11033 19717 11067
rect 19717 11033 19751 11067
rect 19751 11033 19760 11067
rect 19708 11024 19760 11033
rect 20536 11024 20588 11076
rect 21272 11024 21324 11076
rect 21732 11024 21784 11076
rect 22836 11024 22888 11076
rect 15568 10956 15620 11008
rect 21916 10956 21968 11008
rect 24584 10999 24636 11008
rect 24584 10965 24593 10999
rect 24593 10965 24627 10999
rect 24627 10965 24636 10999
rect 24584 10956 24636 10965
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 15752 10795 15804 10804
rect 15752 10761 15761 10795
rect 15761 10761 15795 10795
rect 15795 10761 15804 10795
rect 15752 10752 15804 10761
rect 16396 10795 16448 10804
rect 16396 10761 16405 10795
rect 16405 10761 16439 10795
rect 16439 10761 16448 10795
rect 16396 10752 16448 10761
rect 16948 10752 17000 10804
rect 17684 10752 17736 10804
rect 19340 10684 19392 10736
rect 18328 10616 18380 10668
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 19984 10616 20036 10668
rect 17040 10548 17092 10600
rect 21088 10684 21140 10736
rect 20720 10616 20772 10668
rect 22560 10752 22612 10804
rect 21916 10684 21968 10736
rect 22100 10659 22152 10668
rect 22100 10625 22109 10659
rect 22109 10625 22143 10659
rect 22143 10625 22152 10659
rect 22100 10616 22152 10625
rect 24860 10684 24912 10736
rect 24584 10548 24636 10600
rect 24676 10591 24728 10600
rect 24676 10557 24685 10591
rect 24685 10557 24719 10591
rect 24719 10557 24728 10591
rect 24676 10548 24728 10557
rect 22468 10480 22520 10532
rect 21180 10412 21232 10464
rect 21272 10455 21324 10464
rect 21272 10421 21281 10455
rect 21281 10421 21315 10455
rect 21315 10421 21324 10455
rect 21272 10412 21324 10421
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 18328 10208 18380 10260
rect 19432 10251 19484 10260
rect 19432 10217 19441 10251
rect 19441 10217 19475 10251
rect 19475 10217 19484 10251
rect 19432 10208 19484 10217
rect 20720 10251 20772 10260
rect 20720 10217 20729 10251
rect 20729 10217 20763 10251
rect 20763 10217 20772 10251
rect 20720 10208 20772 10217
rect 21640 10251 21692 10260
rect 21640 10217 21670 10251
rect 21670 10217 21692 10251
rect 21640 10208 21692 10217
rect 21824 10208 21876 10260
rect 16580 10140 16632 10192
rect 21272 10072 21324 10124
rect 21364 10115 21416 10124
rect 21364 10081 21373 10115
rect 21373 10081 21407 10115
rect 21407 10081 21416 10115
rect 21364 10072 21416 10081
rect 22836 10140 22888 10192
rect 23848 10072 23900 10124
rect 19616 10047 19668 10056
rect 19616 10013 19625 10047
rect 19625 10013 19659 10047
rect 19659 10013 19668 10047
rect 19616 10004 19668 10013
rect 20720 10004 20772 10056
rect 23572 10004 23624 10056
rect 25412 10004 25464 10056
rect 21732 9936 21784 9988
rect 21916 9936 21968 9988
rect 23848 9911 23900 9920
rect 23848 9877 23857 9911
rect 23857 9877 23891 9911
rect 23891 9877 23900 9911
rect 23848 9868 23900 9877
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 21732 9664 21784 9716
rect 8484 9528 8536 9580
rect 19340 9596 19392 9648
rect 20076 9596 20128 9648
rect 20720 9596 20772 9648
rect 17132 9460 17184 9512
rect 20812 9528 20864 9580
rect 20904 9571 20956 9580
rect 20904 9537 20913 9571
rect 20913 9537 20947 9571
rect 20947 9537 20956 9571
rect 20904 9528 20956 9537
rect 21548 9528 21600 9580
rect 21916 9528 21968 9580
rect 23296 9639 23348 9648
rect 23296 9605 23305 9639
rect 23305 9605 23339 9639
rect 23339 9605 23348 9639
rect 23296 9596 23348 9605
rect 22468 9528 22520 9580
rect 16212 9392 16264 9444
rect 18052 9367 18104 9376
rect 18052 9333 18061 9367
rect 18061 9333 18095 9367
rect 18095 9333 18104 9367
rect 18052 9324 18104 9333
rect 22284 9460 22336 9512
rect 24768 9503 24820 9512
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 19432 9392 19484 9444
rect 19984 9367 20036 9376
rect 19984 9333 19993 9367
rect 19993 9333 20027 9367
rect 20027 9333 20036 9367
rect 19984 9324 20036 9333
rect 20904 9324 20956 9376
rect 22468 9392 22520 9444
rect 24952 9392 25004 9444
rect 24584 9324 24636 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 14464 9120 14516 9172
rect 18052 9120 18104 9172
rect 19340 9052 19392 9104
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 22284 9120 22336 9172
rect 22652 9052 22704 9104
rect 20628 8984 20680 9036
rect 20904 8916 20956 8968
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 24860 8984 24912 9036
rect 22652 8959 22704 8968
rect 22652 8925 22661 8959
rect 22661 8925 22695 8959
rect 22695 8925 22704 8959
rect 22652 8916 22704 8925
rect 6828 8848 6880 8900
rect 12532 8848 12584 8900
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 19892 8576 19944 8628
rect 19984 8576 20036 8628
rect 22376 8576 22428 8628
rect 13544 8440 13596 8492
rect 19064 8372 19116 8424
rect 22008 8440 22060 8492
rect 22468 8440 22520 8492
rect 24952 8440 25004 8492
rect 19248 8304 19300 8356
rect 24676 8304 24728 8356
rect 24860 8304 24912 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 23940 8032 23992 8084
rect 15108 7964 15160 8016
rect 18696 7828 18748 7880
rect 23480 7896 23532 7948
rect 24952 7896 25004 7948
rect 22376 7828 22428 7880
rect 25044 7828 25096 7880
rect 25872 7760 25924 7812
rect 20720 7735 20772 7744
rect 20720 7701 20729 7735
rect 20729 7701 20763 7735
rect 20763 7701 20772 7735
rect 20720 7692 20772 7701
rect 23480 7692 23532 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 22652 7488 22704 7540
rect 20720 7420 20772 7472
rect 20260 7352 20312 7404
rect 21088 7352 21140 7404
rect 24860 7420 24912 7472
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 25688 7284 25740 7336
rect 23388 7216 23440 7268
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 24860 6808 24912 6860
rect 21180 6740 21232 6792
rect 24584 6740 24636 6792
rect 25044 6672 25096 6724
rect 25228 6604 25280 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 24860 6332 24912 6384
rect 22284 6307 22336 6316
rect 22284 6273 22293 6307
rect 22293 6273 22327 6307
rect 22327 6273 22336 6307
rect 22284 6264 22336 6273
rect 25596 6264 25648 6316
rect 24768 6239 24820 6248
rect 24768 6205 24777 6239
rect 24777 6205 24811 6239
rect 24811 6205 24820 6239
rect 24768 6196 24820 6205
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 22008 5899 22060 5908
rect 22008 5865 22017 5899
rect 22017 5865 22051 5899
rect 22051 5865 22060 5899
rect 22008 5856 22060 5865
rect 23664 5788 23716 5840
rect 21824 5652 21876 5704
rect 22376 5720 22428 5772
rect 23296 5720 23348 5772
rect 24952 5720 25004 5772
rect 23480 5652 23532 5704
rect 24952 5584 25004 5636
rect 23480 5516 23532 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 20904 5244 20956 5296
rect 22744 5176 22796 5228
rect 24676 5151 24728 5160
rect 24676 5117 24685 5151
rect 24685 5117 24719 5151
rect 24719 5117 24728 5151
rect 24676 5108 24728 5117
rect 24952 5040 25004 5092
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 22376 4811 22428 4820
rect 22376 4777 22385 4811
rect 22385 4777 22419 4811
rect 22419 4777 22428 4811
rect 22376 4768 22428 4777
rect 22652 4607 22704 4616
rect 22652 4573 22661 4607
rect 22661 4573 22695 4607
rect 22695 4573 22704 4607
rect 22652 4564 22704 4573
rect 23388 4564 23440 4616
rect 24952 4496 25004 4548
rect 23572 4428 23624 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 21916 4088 21968 4140
rect 18972 4020 19024 4072
rect 20168 4020 20220 4072
rect 25044 4088 25096 4140
rect 25780 4088 25832 4140
rect 22100 3952 22152 4004
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 24952 3952 25004 4004
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 20536 3476 20588 3528
rect 23480 3476 23532 3528
rect 23664 3476 23716 3528
rect 22008 3451 22060 3460
rect 22008 3417 22017 3451
rect 22017 3417 22051 3451
rect 22051 3417 22060 3451
rect 22008 3408 22060 3417
rect 25136 3408 25188 3460
rect 24584 3383 24636 3392
rect 24584 3349 24593 3383
rect 24593 3349 24627 3383
rect 24627 3349 24636 3383
rect 24584 3340 24636 3349
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 25320 3136 25372 3188
rect 24860 3068 24912 3120
rect 25228 3068 25280 3120
rect 19616 3000 19668 3052
rect 23572 3000 23624 3052
rect 24124 3043 24176 3052
rect 24124 3009 24133 3043
rect 24133 3009 24167 3043
rect 24167 3009 24176 3043
rect 24124 3000 24176 3009
rect 19524 2932 19576 2984
rect 25044 2932 25096 2984
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 6828 2635 6880 2644
rect 6828 2601 6837 2635
rect 6837 2601 6871 2635
rect 6871 2601 6880 2635
rect 6828 2592 6880 2601
rect 19524 2592 19576 2644
rect 22192 2592 22244 2644
rect 6920 2388 6972 2440
rect 22744 2388 22796 2440
rect 24584 2388 24636 2440
rect 23388 2320 23440 2372
rect 24952 2320 25004 2372
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
<< metal2 >>
rect 1674 26200 1730 27000
rect 2042 26200 2098 27000
rect 2134 26208 2190 26217
rect 1306 23760 1362 23769
rect 1306 23695 1308 23704
rect 1360 23695 1362 23704
rect 1308 23666 1360 23672
rect 1306 22672 1362 22681
rect 1306 22607 1308 22616
rect 1360 22607 1362 22616
rect 1308 22578 1360 22584
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 20058 1624 20198
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1688 19310 1716 26200
rect 1952 24948 2004 24954
rect 1952 24890 2004 24896
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1964 18970 1992 24890
rect 2056 19922 2084 26200
rect 2410 26200 2466 27000
rect 2778 26466 2834 27000
rect 2778 26450 3096 26466
rect 2778 26444 3108 26450
rect 2778 26438 3056 26444
rect 2778 26200 2834 26438
rect 3056 26386 3108 26392
rect 3146 26330 3202 27000
rect 3332 26444 3384 26450
rect 3332 26386 3384 26392
rect 2884 26302 3202 26330
rect 2134 26143 2190 26152
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1582 18864 1638 18873
rect 1582 18799 1638 18808
rect 1596 18426 1624 18799
rect 2148 18766 2176 26143
rect 2424 22166 2452 26200
rect 2778 24848 2834 24857
rect 2778 24783 2834 24792
rect 2792 23186 2820 24783
rect 2780 23180 2832 23186
rect 2780 23122 2832 23128
rect 2792 22778 2820 23122
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2412 22160 2464 22166
rect 2412 22102 2464 22108
rect 2780 22160 2832 22166
rect 2780 22102 2832 22108
rect 2228 21684 2280 21690
rect 2228 21626 2280 21632
rect 2240 20942 2268 21626
rect 2792 21010 2820 22102
rect 2884 22098 2912 26302
rect 3146 26200 3202 26302
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2780 21004 2832 21010
rect 2780 20946 2832 20952
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 3344 20398 3372 26386
rect 3514 26200 3570 27000
rect 3882 26330 3938 27000
rect 3882 26302 4108 26330
rect 3882 26200 3938 26302
rect 3422 25936 3478 25945
rect 3422 25871 3478 25880
rect 3436 21622 3464 25871
rect 3424 21616 3476 21622
rect 3424 21558 3476 21564
rect 3528 21486 3556 26200
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3792 22636 3844 22642
rect 3792 22578 3844 22584
rect 3698 22128 3754 22137
rect 3698 22063 3754 22072
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3606 21448 3662 21457
rect 3606 21383 3662 21392
rect 3424 21072 3476 21078
rect 3424 21014 3476 21020
rect 3332 20392 3384 20398
rect 3332 20334 3384 20340
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2226 19952 2282 19961
rect 2226 19887 2282 19896
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2240 18426 2268 19887
rect 2320 19848 2372 19854
rect 2320 19790 2372 19796
rect 2332 19417 2360 19790
rect 2318 19408 2374 19417
rect 2318 19343 2374 19352
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2884 18290 2912 19110
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3436 17678 3464 21014
rect 3620 19378 3648 21383
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3712 18970 3740 22063
rect 3700 18964 3752 18970
rect 3700 18906 3752 18912
rect 3712 18834 3740 18906
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 3804 18426 3832 22578
rect 3896 19514 3924 24142
rect 4080 22522 4108 26302
rect 4250 26200 4306 27000
rect 4618 26330 4674 27000
rect 4356 26302 4674 26330
rect 4986 26330 5042 27000
rect 5354 26330 5410 27000
rect 4158 24304 4214 24313
rect 4158 24239 4214 24248
rect 4172 24206 4200 24239
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4264 22710 4292 26200
rect 4356 23050 4384 26302
rect 4618 26200 4674 26302
rect 4896 26308 4948 26314
rect 4896 26250 4948 26256
rect 4986 26302 5120 26330
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4816 23730 4844 24550
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4344 23044 4396 23050
rect 4344 22986 4396 22992
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4724 22778 4752 22918
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4252 22704 4304 22710
rect 4252 22646 4304 22652
rect 4080 22494 4292 22522
rect 4068 22432 4120 22438
rect 4068 22374 4120 22380
rect 4160 22432 4212 22438
rect 4160 22374 4212 22380
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3988 21146 4016 21966
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 4080 20913 4108 22374
rect 4172 21554 4200 22374
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4264 21010 4292 22494
rect 4908 22094 4936 26250
rect 4986 26200 5042 26302
rect 4988 24336 5040 24342
rect 4988 24278 5040 24284
rect 4816 22066 4936 22094
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4252 21004 4304 21010
rect 4252 20946 4304 20952
rect 4066 20904 4122 20913
rect 4066 20839 4122 20848
rect 4080 20318 4384 20346
rect 4080 20262 4108 20318
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3988 17338 4016 19994
rect 4068 18896 4120 18902
rect 4068 18838 4120 18844
rect 4080 18290 4108 18838
rect 4172 18766 4200 20198
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 4080 15162 4108 18022
rect 4356 17610 4384 20318
rect 4526 19816 4582 19825
rect 4526 19751 4582 19760
rect 4540 19718 4568 19751
rect 4528 19712 4580 19718
rect 4528 19654 4580 19660
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4540 17882 4568 19246
rect 4528 17876 4580 17882
rect 4528 17818 4580 17824
rect 4344 17604 4396 17610
rect 4344 17546 4396 17552
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 4540 12889 4568 17478
rect 4632 14521 4660 21966
rect 4712 20528 4764 20534
rect 4712 20470 4764 20476
rect 4724 19854 4752 20470
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4710 19272 4766 19281
rect 4710 19207 4766 19216
rect 4724 18766 4752 19207
rect 4816 18970 4844 22066
rect 4896 21956 4948 21962
rect 4896 21898 4948 21904
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4816 18766 4844 18906
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4908 18426 4936 21898
rect 5000 20602 5028 24278
rect 5092 21486 5120 26302
rect 5184 26302 5410 26330
rect 5448 26376 5500 26382
rect 5448 26318 5500 26324
rect 5184 23798 5212 26302
rect 5354 26200 5410 26302
rect 5262 24984 5318 24993
rect 5262 24919 5318 24928
rect 5172 23792 5224 23798
rect 5172 23734 5224 23740
rect 5276 23576 5304 24919
rect 5460 23882 5488 26318
rect 5722 26200 5778 27000
rect 6090 26200 6146 27000
rect 6458 26330 6514 27000
rect 6196 26302 6514 26330
rect 5184 23548 5304 23576
rect 5368 23854 5488 23882
rect 5080 21480 5132 21486
rect 5080 21422 5132 21428
rect 5184 20602 5212 23548
rect 5368 23474 5396 23854
rect 5448 23724 5500 23730
rect 5448 23666 5500 23672
rect 5276 23446 5396 23474
rect 4988 20596 5040 20602
rect 4988 20538 5040 20544
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 5276 20534 5304 23446
rect 5356 22568 5408 22574
rect 5356 22510 5408 22516
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 4988 18624 5040 18630
rect 4988 18566 5040 18572
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4710 17776 4766 17785
rect 4710 17711 4766 17720
rect 4724 17678 4752 17711
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4724 16182 4752 16390
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4618 14512 4674 14521
rect 4618 14447 4674 14456
rect 4526 12880 4582 12889
rect 4526 12815 4582 12824
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 5000 12306 5028 18566
rect 5092 17066 5120 19926
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5184 19514 5212 19790
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5170 18728 5226 18737
rect 5368 18714 5396 22510
rect 5460 19378 5488 23666
rect 5736 22710 5764 26200
rect 6000 25084 6052 25090
rect 6000 25026 6052 25032
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 5724 22704 5776 22710
rect 5724 22646 5776 22652
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5552 20369 5580 20402
rect 5538 20360 5594 20369
rect 5538 20295 5594 20304
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5276 18698 5396 18714
rect 5170 18663 5226 18672
rect 5264 18692 5396 18698
rect 5184 18630 5212 18663
rect 5316 18686 5396 18692
rect 5264 18634 5316 18640
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5552 18290 5580 19654
rect 5736 18426 5764 20878
rect 5816 20800 5868 20806
rect 5816 20742 5868 20748
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5632 18216 5684 18222
rect 5630 18184 5632 18193
rect 5684 18184 5686 18193
rect 5630 18119 5686 18128
rect 5828 17678 5856 20742
rect 5920 18970 5948 23054
rect 6012 19378 6040 25026
rect 6104 22098 6132 26200
rect 6196 24274 6224 26302
rect 6458 26200 6514 26302
rect 6826 26200 6882 27000
rect 7194 26200 7250 27000
rect 7562 26200 7618 27000
rect 7930 26330 7986 27000
rect 7668 26302 7986 26330
rect 6550 25120 6606 25129
rect 6550 25055 6606 25064
rect 6366 24712 6422 24721
rect 6366 24647 6422 24656
rect 6184 24268 6236 24274
rect 6184 24210 6236 24216
rect 6182 23624 6238 23633
rect 6182 23559 6238 23568
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 5908 18964 5960 18970
rect 5908 18906 5960 18912
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6012 18426 6040 18702
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6104 18358 6132 20198
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 6196 17746 6224 23559
rect 6276 23044 6328 23050
rect 6276 22986 6328 22992
rect 6288 22273 6316 22986
rect 6380 22930 6408 24647
rect 6564 24410 6592 25055
rect 6736 24880 6788 24886
rect 6736 24822 6788 24828
rect 6552 24404 6604 24410
rect 6552 24346 6604 24352
rect 6644 24404 6696 24410
rect 6644 24346 6696 24352
rect 6656 24206 6684 24346
rect 6644 24200 6696 24206
rect 6644 24142 6696 24148
rect 6460 24064 6512 24070
rect 6460 24006 6512 24012
rect 6472 23050 6500 24006
rect 6748 23662 6776 24822
rect 6644 23656 6696 23662
rect 6644 23598 6696 23604
rect 6736 23656 6788 23662
rect 6736 23598 6788 23604
rect 6656 23322 6684 23598
rect 6644 23316 6696 23322
rect 6644 23258 6696 23264
rect 6460 23044 6512 23050
rect 6460 22986 6512 22992
rect 6380 22902 6500 22930
rect 6274 22264 6330 22273
rect 6274 22199 6330 22208
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5538 17232 5594 17241
rect 5538 17167 5540 17176
rect 5592 17167 5594 17176
rect 5540 17138 5592 17144
rect 5080 17060 5132 17066
rect 5080 17002 5132 17008
rect 5262 16688 5318 16697
rect 5262 16623 5264 16632
rect 5316 16623 5318 16632
rect 5264 16594 5316 16600
rect 6288 15978 6316 20878
rect 6380 17882 6408 21966
rect 6472 19310 6500 22902
rect 6644 22636 6696 22642
rect 6644 22578 6696 22584
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6472 18766 6500 19246
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 6472 17921 6500 18566
rect 6458 17912 6514 17921
rect 6368 17876 6420 17882
rect 6458 17847 6514 17856
rect 6368 17818 6420 17824
rect 6564 17746 6592 21286
rect 6656 19718 6684 22578
rect 6840 22094 6868 26200
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 6920 23656 6972 23662
rect 6918 23624 6920 23633
rect 6972 23624 6974 23633
rect 6918 23559 6974 23568
rect 7024 23526 7052 24142
rect 7102 23624 7158 23633
rect 7102 23559 7104 23568
rect 7156 23559 7158 23568
rect 7104 23530 7156 23536
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 7102 22672 7158 22681
rect 7102 22607 7158 22616
rect 6840 22066 7052 22094
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6748 20874 6776 21490
rect 7024 21010 7052 22066
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 6920 20936 6972 20942
rect 6920 20878 6972 20884
rect 6736 20868 6788 20874
rect 6736 20810 6788 20816
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6748 19854 6776 19994
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6644 19712 6696 19718
rect 6644 19654 6696 19660
rect 6932 19394 6960 20878
rect 6932 19366 7052 19394
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 6644 18624 6696 18630
rect 6644 18566 6696 18572
rect 6656 17814 6684 18566
rect 6932 18290 6960 19178
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 7024 17882 7052 19366
rect 7116 19310 7144 22607
rect 7208 21468 7236 26200
rect 7576 23798 7604 26200
rect 7564 23792 7616 23798
rect 7564 23734 7616 23740
rect 7380 23316 7432 23322
rect 7380 23258 7432 23264
rect 7288 23248 7340 23254
rect 7288 23190 7340 23196
rect 7300 21593 7328 23190
rect 7392 22710 7420 23258
rect 7472 23248 7524 23254
rect 7472 23190 7524 23196
rect 7562 23216 7618 23225
rect 7380 22704 7432 22710
rect 7380 22646 7432 22652
rect 7380 22024 7432 22030
rect 7378 21992 7380 22001
rect 7432 21992 7434 22001
rect 7378 21927 7434 21936
rect 7286 21584 7342 21593
rect 7286 21519 7342 21528
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7288 21480 7340 21486
rect 7208 21440 7288 21468
rect 7288 21422 7340 21428
rect 7196 20460 7248 20466
rect 7196 20402 7248 20408
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7208 20058 7236 20402
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7116 18290 7144 19246
rect 7104 18284 7156 18290
rect 7104 18226 7156 18232
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 6644 17808 6696 17814
rect 6644 17750 6696 17756
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 7194 17640 7250 17649
rect 7194 17575 7250 17584
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5552 12209 5580 15098
rect 6564 13977 6592 17274
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6840 16794 6868 17138
rect 7116 17105 7144 17478
rect 7208 17338 7236 17575
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7102 17096 7158 17105
rect 7102 17031 7158 17040
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 7300 16046 7328 20402
rect 7392 17338 7420 21490
rect 7484 18834 7512 23190
rect 7562 23151 7618 23160
rect 7576 19378 7604 23151
rect 7668 22982 7696 26302
rect 7930 26200 7986 26302
rect 8298 26200 8354 27000
rect 8666 26200 8722 27000
rect 9034 26330 9090 27000
rect 8772 26302 9090 26330
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7562 19000 7618 19009
rect 7562 18935 7618 18944
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7576 18222 7604 18935
rect 7668 18290 7696 22170
rect 7852 19786 7880 23598
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 8312 22098 8340 26200
rect 8680 24138 8708 26200
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8392 23180 8444 23186
rect 8392 23122 8444 23128
rect 8404 23089 8432 23122
rect 8390 23080 8446 23089
rect 8390 23015 8446 23024
rect 8666 22808 8722 22817
rect 8666 22743 8722 22752
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8482 21720 8538 21729
rect 8482 21655 8538 21664
rect 8496 21622 8524 21655
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 8484 21072 8536 21078
rect 8484 21014 8536 21020
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7746 19136 7802 19145
rect 7746 19071 7802 19080
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7470 18048 7526 18057
rect 7470 17983 7526 17992
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7484 17202 7512 17983
rect 7576 17678 7604 18158
rect 7656 18080 7708 18086
rect 7760 18057 7788 19071
rect 7656 18022 7708 18028
rect 7746 18048 7802 18057
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7484 16794 7512 17138
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7668 15065 7696 18022
rect 7746 17983 7802 17992
rect 7852 17864 7880 19314
rect 8220 18970 8248 19382
rect 8312 19378 8340 19654
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7760 17836 7880 17864
rect 7760 16114 7788 17836
rect 7838 17776 7894 17785
rect 7838 17711 7894 17720
rect 7852 17134 7880 17711
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8312 17270 8340 18770
rect 8404 18766 8432 20198
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8496 18290 8524 21014
rect 8574 19408 8630 19417
rect 8574 19343 8576 19352
rect 8628 19343 8630 19352
rect 8576 19314 8628 19320
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8588 18426 8616 18702
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8404 17338 8432 17478
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 8128 16504 8156 17070
rect 8680 16658 8708 22743
rect 8772 22710 8800 26302
rect 9034 26200 9090 26302
rect 9402 26200 9458 27000
rect 9770 26330 9826 27000
rect 9692 26302 9826 26330
rect 9128 25016 9180 25022
rect 9128 24958 9180 24964
rect 9140 24342 9168 24958
rect 9128 24336 9180 24342
rect 9128 24278 9180 24284
rect 8850 24032 8906 24041
rect 8850 23967 8906 23976
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8864 22094 8892 23967
rect 9416 23236 9444 26200
rect 9692 24274 9720 26302
rect 9770 26200 9826 26302
rect 10138 26200 10194 27000
rect 10506 26200 10562 27000
rect 10874 26200 10930 27000
rect 11242 26200 11298 27000
rect 11610 26200 11666 27000
rect 11978 26200 12034 27000
rect 12346 26200 12402 27000
rect 12714 26200 12770 27000
rect 13082 26330 13138 27000
rect 13082 26302 13400 26330
rect 13082 26200 13138 26302
rect 9954 24848 10010 24857
rect 9954 24783 10010 24792
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9496 24200 9548 24206
rect 9496 24142 9548 24148
rect 9586 24168 9642 24177
rect 9324 23208 9444 23236
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 9036 22568 9088 22574
rect 9036 22510 9088 22516
rect 9048 22098 9076 22510
rect 8772 22066 8892 22094
rect 9036 22092 9088 22098
rect 8772 18834 8800 22066
rect 9036 22034 9088 22040
rect 9048 21554 9076 22034
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 9048 20466 9076 21490
rect 9232 21146 9260 23122
rect 9324 23118 9352 23208
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9312 21888 9364 21894
rect 9310 21856 9312 21865
rect 9364 21856 9366 21865
rect 9310 21791 9366 21800
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9416 21486 9444 21626
rect 9312 21480 9364 21486
rect 9312 21422 9364 21428
rect 9404 21480 9456 21486
rect 9404 21422 9456 21428
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9324 20942 9352 21422
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9312 20800 9364 20806
rect 9312 20742 9364 20748
rect 9324 20641 9352 20742
rect 9310 20632 9366 20641
rect 9310 20567 9366 20576
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 8852 20324 8904 20330
rect 8852 20266 8904 20272
rect 8864 18970 8892 20266
rect 9048 19378 9076 20402
rect 9310 20088 9366 20097
rect 9310 20023 9366 20032
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 9048 19258 9076 19314
rect 8956 19230 9076 19258
rect 8852 18964 8904 18970
rect 8852 18906 8904 18912
rect 8760 18828 8812 18834
rect 8760 18770 8812 18776
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8772 17066 8800 18634
rect 8956 18290 8984 19230
rect 9140 18766 9168 19654
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9232 18329 9260 19450
rect 9324 18630 9352 20023
rect 9508 19854 9536 24142
rect 9586 24103 9642 24112
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9416 18834 9444 19246
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9218 18320 9274 18329
rect 8944 18284 8996 18290
rect 9218 18255 9274 18264
rect 8944 18226 8996 18232
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8864 17649 8892 18090
rect 8956 17746 8984 18226
rect 9402 17912 9458 17921
rect 9128 17876 9180 17882
rect 9402 17847 9458 17856
rect 9128 17818 9180 17824
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8850 17640 8906 17649
rect 8850 17575 8906 17584
rect 8956 17202 8984 17682
rect 9140 17678 9168 17818
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 9416 17241 9444 17847
rect 9508 17610 9536 18770
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9402 17232 9458 17241
rect 8944 17196 8996 17202
rect 9402 17167 9458 17176
rect 8944 17138 8996 17144
rect 8760 17060 8812 17066
rect 8760 17002 8812 17008
rect 9310 16824 9366 16833
rect 9310 16759 9366 16768
rect 9324 16726 9352 16759
rect 9312 16720 9364 16726
rect 9312 16662 9364 16668
rect 9600 16658 9628 24103
rect 9968 22094 9996 24783
rect 10152 23798 10180 26200
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 9876 22066 9996 22094
rect 9678 21856 9734 21865
rect 9678 21791 9734 21800
rect 9692 19009 9720 21791
rect 9678 19000 9734 19009
rect 9678 18935 9734 18944
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9784 18170 9812 18906
rect 9692 18142 9812 18170
rect 9692 16794 9720 18142
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9784 17270 9812 18022
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 9588 16652 9640 16658
rect 9876 16640 9904 22066
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 10060 21690 10088 21830
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10048 21072 10100 21078
rect 10048 21014 10100 21020
rect 10060 20398 10088 21014
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 10140 17604 10192 17610
rect 10140 17546 10192 17552
rect 10060 17134 10088 17546
rect 10152 17270 10180 17546
rect 10140 17264 10192 17270
rect 10140 17206 10192 17212
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 9968 16708 9996 17070
rect 10152 16998 10180 17206
rect 10048 16992 10100 16998
rect 10046 16960 10048 16969
rect 10140 16992 10192 16998
rect 10100 16960 10102 16969
rect 10140 16934 10192 16940
rect 10046 16895 10102 16904
rect 10140 16720 10192 16726
rect 9968 16680 10140 16708
rect 10140 16662 10192 16668
rect 9876 16612 9996 16640
rect 9588 16594 9640 16600
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 7852 16476 8156 16504
rect 7852 16250 7880 16476
rect 8588 16402 8616 16526
rect 8758 16416 8814 16425
rect 8588 16374 8758 16402
rect 7950 16348 8258 16357
rect 8758 16351 8814 16360
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8220 16114 8248 16186
rect 8666 16144 8722 16153
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 8208 16108 8260 16114
rect 8666 16079 8668 16088
rect 8208 16050 8260 16056
rect 8720 16079 8722 16088
rect 8668 16050 8720 16056
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7654 15056 7710 15065
rect 7654 14991 7710 15000
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 6550 13968 6606 13977
rect 6550 13903 6606 13912
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 5538 12200 5594 12209
rect 5538 12135 5594 12144
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 8496 9586 8524 15846
rect 8772 15706 8800 16351
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 9126 16008 9182 16017
rect 9508 15994 9536 16118
rect 9600 16114 9628 16594
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9784 16289 9812 16390
rect 9770 16280 9826 16289
rect 9770 16215 9826 16224
rect 9876 16114 9904 16390
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9508 15966 9720 15994
rect 9126 15943 9128 15952
rect 9180 15943 9182 15952
rect 9128 15914 9180 15920
rect 9692 15881 9720 15966
rect 9678 15872 9734 15881
rect 9678 15807 9734 15816
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 9968 15502 9996 16612
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10152 16250 10180 16390
rect 10244 16289 10272 24006
rect 10520 23186 10548 26200
rect 10598 23896 10654 23905
rect 10598 23831 10654 23840
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10416 22704 10468 22710
rect 10416 22646 10468 22652
rect 10428 21554 10456 22646
rect 10416 21548 10468 21554
rect 10416 21490 10468 21496
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10428 20806 10456 21082
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10520 20806 10548 20946
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10508 20800 10560 20806
rect 10508 20742 10560 20748
rect 10336 20602 10364 20742
rect 10324 20596 10376 20602
rect 10324 20538 10376 20544
rect 10322 19544 10378 19553
rect 10322 19479 10378 19488
rect 10336 18970 10364 19479
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10414 18456 10470 18465
rect 10414 18391 10470 18400
rect 10428 16833 10456 18391
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10520 17610 10548 18294
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10612 17354 10640 23831
rect 10888 23798 10916 26200
rect 11256 24274 11284 26200
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 10876 23792 10928 23798
rect 10876 23734 10928 23740
rect 11518 23760 11574 23769
rect 11518 23695 11574 23704
rect 11336 22500 11388 22506
rect 11336 22442 11388 22448
rect 11152 22432 11204 22438
rect 10966 22400 11022 22409
rect 11152 22374 11204 22380
rect 11244 22432 11296 22438
rect 11244 22374 11296 22380
rect 10966 22335 11022 22344
rect 10980 21962 11008 22335
rect 11060 22092 11112 22098
rect 11060 22034 11112 22040
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10704 21350 10732 21422
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10876 21344 10928 21350
rect 10876 21286 10928 21292
rect 10796 21078 10824 21286
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 10888 20806 10916 21286
rect 11072 21010 11100 22034
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 11164 20874 11192 22374
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 11152 20868 11204 20874
rect 11152 20810 11204 20816
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10980 20602 11008 20810
rect 10968 20596 11020 20602
rect 10968 20538 11020 20544
rect 11164 20505 11192 20810
rect 11150 20496 11206 20505
rect 11150 20431 11206 20440
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10796 20074 10824 20198
rect 10796 20046 11100 20074
rect 10796 19514 10824 20046
rect 11072 19922 11100 20046
rect 11256 19938 11284 22374
rect 11348 22098 11376 22442
rect 11336 22092 11388 22098
rect 11336 22034 11388 22040
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 11440 21554 11468 21898
rect 11428 21548 11480 21554
rect 11428 21490 11480 21496
rect 11440 20874 11468 21490
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 11440 20534 11468 20810
rect 11428 20528 11480 20534
rect 11428 20470 11480 20476
rect 10968 19916 11020 19922
rect 10968 19858 11020 19864
rect 11060 19916 11112 19922
rect 11256 19910 11468 19938
rect 11060 19858 11112 19864
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10782 19408 10838 19417
rect 10782 19343 10838 19352
rect 10796 19258 10824 19343
rect 10520 17326 10640 17354
rect 10704 19230 10824 19258
rect 10414 16824 10470 16833
rect 10414 16759 10470 16768
rect 10322 16552 10378 16561
rect 10322 16487 10378 16496
rect 10230 16280 10286 16289
rect 10140 16244 10192 16250
rect 10230 16215 10286 16224
rect 10140 16186 10192 16192
rect 10336 15978 10364 16487
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10046 15600 10102 15609
rect 10046 15535 10102 15544
rect 10060 15502 10088 15535
rect 9496 15496 9548 15502
rect 9496 15438 9548 15444
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9508 15162 9536 15438
rect 10060 15162 10088 15438
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10520 15026 10548 17326
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10520 14618 10548 14962
rect 10612 14958 10640 16934
rect 10704 16182 10732 19230
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10796 18222 10824 19110
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10888 16590 10916 19654
rect 10980 19174 11008 19858
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 11164 18902 11192 19110
rect 11256 18970 11284 19790
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10796 15910 10824 16390
rect 10980 16046 11008 18226
rect 11164 17882 11192 18838
rect 11334 18592 11390 18601
rect 11334 18527 11390 18536
rect 11348 18358 11376 18527
rect 11336 18352 11388 18358
rect 11336 18294 11388 18300
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11256 16590 11284 16730
rect 11348 16658 11376 18294
rect 11440 17542 11468 19910
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10704 14958 10732 15370
rect 11164 15366 11192 16390
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10704 14414 10732 14894
rect 11164 14618 11192 14962
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10704 13190 10732 14350
rect 11532 14006 11560 23695
rect 11624 23186 11652 26200
rect 11704 24336 11756 24342
rect 11704 24278 11756 24284
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11624 20097 11652 22646
rect 11610 20088 11666 20097
rect 11610 20023 11666 20032
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11624 19378 11652 19790
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11716 18714 11744 24278
rect 11992 23662 12020 26200
rect 12360 24342 12388 26200
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12348 24336 12400 24342
rect 12348 24278 12400 24284
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11796 23316 11848 23322
rect 11796 23258 11848 23264
rect 11808 23118 11836 23258
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 12070 22944 12126 22953
rect 12070 22879 12126 22888
rect 11794 22536 11850 22545
rect 11794 22471 11850 22480
rect 11888 22500 11940 22506
rect 11624 18686 11744 18714
rect 11624 16969 11652 18686
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11716 18154 11744 18566
rect 11704 18148 11756 18154
rect 11704 18090 11756 18096
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11716 17202 11744 17682
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11610 16960 11666 16969
rect 11610 16895 11666 16904
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11624 15366 11652 16594
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11716 16046 11744 16526
rect 11808 16454 11836 22471
rect 11888 22442 11940 22448
rect 11900 21162 11928 22442
rect 12084 22234 12112 22879
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12072 22228 12124 22234
rect 12072 22170 12124 22176
rect 12164 22228 12216 22234
rect 12164 22170 12216 22176
rect 11980 21888 12032 21894
rect 12176 21876 12204 22170
rect 12268 22098 12296 22510
rect 12452 22386 12480 24142
rect 12532 23248 12584 23254
rect 12532 23190 12584 23196
rect 12360 22358 12480 22386
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 12032 21848 12204 21876
rect 12256 21888 12308 21894
rect 11980 21830 12032 21836
rect 12256 21830 12308 21836
rect 12268 21554 12296 21830
rect 12256 21548 12308 21554
rect 12256 21490 12308 21496
rect 12254 21312 12310 21321
rect 12254 21247 12310 21256
rect 11900 21134 12020 21162
rect 11886 21040 11942 21049
rect 11886 20975 11942 20984
rect 11900 19145 11928 20975
rect 11992 19310 12020 21134
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12176 19786 12204 20470
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12176 19514 12204 19722
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12268 19334 12296 21247
rect 12360 20482 12388 22358
rect 12438 22264 12494 22273
rect 12544 22234 12572 23190
rect 12636 22778 12664 24550
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12622 22400 12678 22409
rect 12622 22335 12678 22344
rect 12438 22199 12494 22208
rect 12532 22228 12584 22234
rect 12452 21078 12480 22199
rect 12532 22170 12584 22176
rect 12636 22098 12664 22335
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12440 21072 12492 21078
rect 12440 21014 12492 21020
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12452 20754 12480 20878
rect 12636 20754 12664 21422
rect 12728 21321 12756 26200
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12820 23594 12848 24074
rect 12808 23588 12860 23594
rect 12808 23530 12860 23536
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 13004 22506 13032 22578
rect 12992 22500 13044 22506
rect 12992 22442 13044 22448
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 13372 22216 13400 26302
rect 13450 26200 13506 27000
rect 13818 26200 13874 27000
rect 14186 26330 14242 27000
rect 13924 26302 14242 26330
rect 13464 23254 13492 26200
rect 13728 25084 13780 25090
rect 13728 25026 13780 25032
rect 13740 23866 13768 25026
rect 13832 24041 13860 26200
rect 13818 24032 13874 24041
rect 13818 23967 13874 23976
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 13636 23520 13688 23526
rect 13636 23462 13688 23468
rect 13648 23322 13676 23462
rect 13636 23316 13688 23322
rect 13636 23258 13688 23264
rect 13452 23248 13504 23254
rect 13452 23190 13504 23196
rect 13924 23186 13952 26302
rect 14186 26200 14242 26302
rect 14554 26200 14610 27000
rect 14922 26200 14978 27000
rect 15290 26200 15346 27000
rect 15658 26200 15714 27000
rect 16026 26330 16082 27000
rect 16394 26330 16450 27000
rect 16026 26302 16252 26330
rect 16026 26200 16082 26302
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 14002 23352 14058 23361
rect 14002 23287 14058 23296
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13452 23044 13504 23050
rect 13452 22986 13504 22992
rect 13280 22188 13400 22216
rect 13176 21684 13228 21690
rect 13176 21626 13228 21632
rect 13188 21457 13216 21626
rect 13174 21448 13230 21457
rect 13280 21434 13308 22188
rect 13464 22094 13492 22986
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 13556 22710 13584 22918
rect 13544 22704 13596 22710
rect 13544 22646 13596 22652
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 13648 22438 13676 22578
rect 13636 22432 13688 22438
rect 13740 22420 13768 23054
rect 13740 22392 13860 22420
rect 13636 22374 13688 22380
rect 13372 22066 13492 22094
rect 13636 22092 13688 22098
rect 13372 21690 13400 22066
rect 13636 22034 13688 22040
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13360 21684 13412 21690
rect 13360 21626 13412 21632
rect 13452 21480 13504 21486
rect 13280 21406 13400 21434
rect 13452 21422 13504 21428
rect 13174 21383 13230 21392
rect 12808 21344 12860 21350
rect 12714 21312 12770 21321
rect 12808 21286 12860 21292
rect 12714 21247 12770 21256
rect 12452 20726 12664 20754
rect 12438 20632 12494 20641
rect 12438 20567 12440 20576
rect 12492 20567 12494 20576
rect 12532 20596 12584 20602
rect 12440 20538 12492 20544
rect 12716 20596 12768 20602
rect 12584 20556 12716 20584
rect 12532 20538 12584 20544
rect 12716 20538 12768 20544
rect 12360 20454 12664 20482
rect 12820 20466 12848 21286
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 13266 20904 13322 20913
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 12452 20210 12480 20266
rect 12452 20182 12572 20210
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 12072 19304 12124 19310
rect 12268 19306 12480 19334
rect 12072 19246 12124 19252
rect 11886 19136 11942 19145
rect 11886 19071 11942 19080
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11992 18630 12020 18702
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11900 17746 11928 18566
rect 12084 18426 12112 19246
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12176 18766 12204 19178
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11992 17921 12020 18226
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 11978 17912 12034 17921
rect 11978 17847 12034 17856
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11900 16969 11928 17274
rect 12084 17270 12112 17818
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 11980 16992 12032 16998
rect 11886 16960 11942 16969
rect 11980 16934 12032 16940
rect 11886 16895 11942 16904
rect 11992 16726 12020 16934
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 12176 16454 12204 18158
rect 12268 17882 12296 19110
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12360 18306 12388 18838
rect 12452 18766 12480 19306
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12360 18278 12480 18306
rect 12452 17882 12480 18278
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12348 17740 12400 17746
rect 12544 17728 12572 20182
rect 12636 17785 12664 20454
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 13004 20244 13032 20878
rect 13266 20839 13268 20848
rect 13320 20839 13322 20848
rect 13268 20810 13320 20816
rect 12728 20216 13032 20244
rect 12400 17700 12572 17728
rect 12622 17776 12678 17785
rect 12622 17711 12678 17720
rect 12348 17682 12400 17688
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 11992 16182 12020 16390
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11624 14482 11652 15302
rect 11716 14958 11744 15982
rect 11900 15706 11928 16118
rect 12072 15904 12124 15910
rect 12268 15881 12296 17478
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12544 16522 12572 17070
rect 12636 16969 12664 17274
rect 12622 16960 12678 16969
rect 12622 16895 12678 16904
rect 12532 16516 12584 16522
rect 12532 16458 12584 16464
rect 12544 16182 12572 16458
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12728 16130 12756 20216
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12806 19408 12862 19417
rect 12806 19343 12862 19352
rect 12820 16425 12848 19343
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13372 18834 13400 21406
rect 13464 19990 13492 21422
rect 13556 20777 13584 21898
rect 13648 21146 13676 22034
rect 13832 21185 13860 22392
rect 14016 22094 14044 23287
rect 13924 22066 14044 22094
rect 13924 21865 13952 22066
rect 13910 21856 13966 21865
rect 13910 21791 13966 21800
rect 13818 21176 13874 21185
rect 13636 21140 13688 21146
rect 13818 21111 13874 21120
rect 13636 21082 13688 21088
rect 13726 20904 13782 20913
rect 13726 20839 13782 20848
rect 14004 20868 14056 20874
rect 13636 20800 13688 20806
rect 13542 20768 13598 20777
rect 13636 20742 13688 20748
rect 13542 20703 13598 20712
rect 13544 20528 13596 20534
rect 13544 20470 13596 20476
rect 13556 19990 13584 20470
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 13544 19984 13596 19990
rect 13544 19926 13596 19932
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13464 19174 13492 19722
rect 13556 19446 13584 19926
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 12992 18692 13044 18698
rect 12992 18634 13044 18640
rect 13004 18290 13032 18634
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 13004 17134 13032 17546
rect 13280 17270 13308 17818
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13268 16720 13320 16726
rect 13266 16688 13268 16697
rect 13320 16688 13322 16697
rect 13266 16623 13322 16632
rect 12806 16416 12862 16425
rect 12806 16351 12862 16360
rect 12348 16040 12400 16046
rect 12348 15982 12400 15988
rect 12072 15846 12124 15852
rect 12254 15872 12310 15881
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 12084 14958 12112 15846
rect 12254 15807 12310 15816
rect 12360 15366 12388 15982
rect 12544 15434 12572 16118
rect 12728 16102 12848 16130
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12728 15570 12756 15982
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12348 15360 12400 15366
rect 12348 15302 12400 15308
rect 12544 15094 12572 15370
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 11992 14482 12020 14894
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11886 14376 11942 14385
rect 11886 14311 11942 14320
rect 11520 14000 11572 14006
rect 11520 13942 11572 13948
rect 11900 13870 11928 14311
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 12084 13258 12112 14894
rect 12544 14278 12572 15030
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12544 13530 12572 14214
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12544 13258 12572 13466
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 10060 9042 10088 13126
rect 12544 12986 12572 13194
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 12544 8906 12572 12922
rect 12728 12918 12756 13330
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12820 12753 12848 16102
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13372 14113 13400 18226
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13464 17066 13492 17682
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13450 16688 13506 16697
rect 13450 16623 13506 16632
rect 13464 16046 13492 16623
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13452 14816 13504 14822
rect 13450 14784 13452 14793
rect 13504 14784 13506 14793
rect 13450 14719 13506 14728
rect 13450 14648 13506 14657
rect 13450 14583 13506 14592
rect 13358 14104 13414 14113
rect 13358 14039 13414 14048
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13372 13394 13400 14039
rect 13464 13870 13492 14583
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13360 12776 13412 12782
rect 12806 12744 12862 12753
rect 13360 12718 13412 12724
rect 12806 12679 12862 12688
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 13372 11830 13400 12718
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13464 11694 13492 13398
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 6840 2650 6868 8842
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 13556 8498 13584 17002
rect 13648 15042 13676 20742
rect 13740 18873 13768 20839
rect 14004 20810 14056 20816
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 19514 13860 20198
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13924 19514 13952 19790
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13912 19508 13964 19514
rect 13912 19450 13964 19456
rect 13910 19000 13966 19009
rect 13910 18935 13966 18944
rect 13726 18864 13782 18873
rect 13726 18799 13782 18808
rect 13728 18692 13780 18698
rect 13728 18634 13780 18640
rect 13740 17746 13768 18634
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13832 17218 13860 17818
rect 13740 17190 13860 17218
rect 13740 16658 13768 17190
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13832 15502 13860 17070
rect 13924 16726 13952 18935
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 14016 16640 14044 20810
rect 14108 20806 14136 24686
rect 14568 24138 14596 26200
rect 14556 24132 14608 24138
rect 14556 24074 14608 24080
rect 14936 23746 14964 26200
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 15028 23866 15056 24074
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 14844 23718 14964 23746
rect 14740 23656 14792 23662
rect 14740 23598 14792 23604
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14292 22438 14320 23054
rect 14372 23044 14424 23050
rect 14372 22986 14424 22992
rect 14384 22545 14412 22986
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14660 22778 14688 22918
rect 14752 22778 14780 23598
rect 14844 23322 14872 23718
rect 14924 23656 14976 23662
rect 14924 23598 14976 23604
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14370 22536 14426 22545
rect 14370 22471 14426 22480
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 14370 22400 14426 22409
rect 14292 22030 14320 22374
rect 14752 22386 14780 22714
rect 14370 22335 14426 22344
rect 14660 22358 14780 22386
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14096 20800 14148 20806
rect 14096 20742 14148 20748
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 14108 17202 14136 19926
rect 14200 19854 14228 21490
rect 14292 20262 14320 21966
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14292 20097 14320 20198
rect 14278 20088 14334 20097
rect 14278 20023 14334 20032
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14280 19440 14332 19446
rect 14280 19382 14332 19388
rect 14292 18970 14320 19382
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 14384 18358 14412 22335
rect 14660 22234 14688 22358
rect 14936 22250 14964 23598
rect 14648 22228 14700 22234
rect 14844 22222 14964 22250
rect 14844 22216 14872 22222
rect 14648 22170 14700 22176
rect 14752 22188 14872 22216
rect 14752 22094 14780 22188
rect 15120 22114 15148 24142
rect 14660 22066 14780 22094
rect 14844 22086 15148 22114
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 14476 21146 14504 21354
rect 14554 21312 14610 21321
rect 14554 21247 14610 21256
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14568 20074 14596 21247
rect 14476 20046 14596 20074
rect 14476 19514 14504 20046
rect 14556 19984 14608 19990
rect 14556 19926 14608 19932
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14476 18426 14504 18566
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14278 18048 14334 18057
rect 14278 17983 14334 17992
rect 14292 17542 14320 17983
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14476 16998 14504 17478
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14016 16612 14136 16640
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 13912 15904 13964 15910
rect 13912 15846 13964 15852
rect 13924 15706 13952 15846
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13910 15464 13966 15473
rect 13910 15399 13966 15408
rect 13924 15366 13952 15399
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13648 15014 13768 15042
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13648 14618 13676 14826
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13740 14074 13768 15014
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13832 14550 13860 14962
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13924 14414 13952 15302
rect 14016 15094 14044 16050
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13832 13818 13860 14010
rect 13740 13802 13952 13818
rect 13728 13796 13952 13802
rect 13780 13790 13952 13796
rect 13728 13738 13780 13744
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13740 13190 13768 13466
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12442 13768 13126
rect 13924 12442 13952 13790
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 13740 11830 13768 12378
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 14108 11626 14136 16612
rect 14568 16266 14596 19926
rect 14384 16238 14596 16266
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 14200 13258 14228 15506
rect 14292 14482 14320 15506
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14292 14006 14320 14418
rect 14384 14074 14412 16238
rect 14660 16130 14688 22066
rect 14738 21584 14794 21593
rect 14738 21519 14794 21528
rect 14752 21010 14780 21519
rect 14740 21004 14792 21010
rect 14740 20946 14792 20952
rect 14738 20224 14794 20233
rect 14738 20159 14794 20168
rect 14752 19417 14780 20159
rect 14844 19514 14872 22086
rect 15014 21584 15070 21593
rect 15014 21519 15070 21528
rect 15200 21548 15252 21554
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 14738 19408 14794 19417
rect 14738 19343 14794 19352
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14936 18834 14964 19314
rect 14924 18828 14976 18834
rect 14924 18770 14976 18776
rect 14936 18442 14964 18770
rect 14844 18414 14964 18442
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 14752 17746 14780 18294
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 14752 17202 14780 17546
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14752 16794 14780 16934
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14844 16522 14872 18414
rect 14924 17740 14976 17746
rect 14924 17682 14976 17688
rect 14936 16658 14964 17682
rect 15028 17082 15056 21519
rect 15200 21490 15252 21496
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15120 20262 15148 21422
rect 15108 20256 15160 20262
rect 15108 20198 15160 20204
rect 15120 19310 15148 20198
rect 15212 19786 15240 21490
rect 15304 20058 15332 26200
rect 15384 23860 15436 23866
rect 15384 23802 15436 23808
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15200 19780 15252 19786
rect 15200 19722 15252 19728
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15212 18986 15240 19722
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15304 19417 15332 19654
rect 15290 19408 15346 19417
rect 15290 19343 15346 19352
rect 15212 18958 15332 18986
rect 15304 18698 15332 18958
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15120 17785 15148 18226
rect 15106 17776 15162 17785
rect 15212 17746 15240 18566
rect 15106 17711 15162 17720
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15028 17054 15148 17082
rect 14924 16652 14976 16658
rect 14924 16594 14976 16600
rect 14832 16516 14884 16522
rect 14476 16102 14688 16130
rect 14752 16476 14832 16504
rect 14476 15434 14504 16102
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14464 15428 14516 15434
rect 14464 15370 14516 15376
rect 14568 14482 14596 15982
rect 14646 15736 14702 15745
rect 14646 15671 14702 15680
rect 14660 14618 14688 15671
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14556 14476 14608 14482
rect 14608 14436 14688 14464
rect 14556 14418 14608 14424
rect 14660 14074 14688 14436
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14280 14000 14332 14006
rect 14752 13954 14780 16476
rect 14832 16458 14884 16464
rect 15016 16516 15068 16522
rect 15016 16458 15068 16464
rect 15028 15910 15056 16458
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 15028 15434 15056 15846
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14830 14920 14886 14929
rect 14830 14855 14886 14864
rect 14844 14822 14872 14855
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14936 14618 14964 15098
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 15028 14346 15056 15370
rect 15120 15026 15148 17054
rect 15212 16697 15240 17138
rect 15304 17134 15332 18634
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15198 16688 15254 16697
rect 15198 16623 15254 16632
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 14280 13942 14332 13948
rect 14292 13394 14320 13942
rect 14476 13926 14780 13954
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14292 12986 14320 13330
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14292 12782 14320 12922
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 14476 9178 14504 13926
rect 15028 13920 15056 14282
rect 15212 14278 15240 15982
rect 15396 15094 15424 23802
rect 15672 22817 15700 26200
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 16040 24274 16068 24890
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 16120 23724 16172 23730
rect 16120 23666 16172 23672
rect 15934 23624 15990 23633
rect 15934 23559 15990 23568
rect 15844 23520 15896 23526
rect 15844 23462 15896 23468
rect 15856 23050 15884 23462
rect 15844 23044 15896 23050
rect 15844 22986 15896 22992
rect 15658 22808 15714 22817
rect 15856 22778 15884 22986
rect 15658 22743 15714 22752
rect 15844 22772 15896 22778
rect 15844 22714 15896 22720
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15660 22160 15712 22166
rect 15660 22102 15712 22108
rect 15672 21486 15700 22102
rect 15476 21480 15528 21486
rect 15660 21480 15712 21486
rect 15476 21422 15528 21428
rect 15566 21448 15622 21457
rect 15488 20942 15516 21422
rect 15660 21422 15712 21428
rect 15566 21383 15622 21392
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15488 20806 15516 20878
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15488 18970 15516 20742
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15488 18358 15516 18770
rect 15476 18352 15528 18358
rect 15476 18294 15528 18300
rect 15474 17776 15530 17785
rect 15474 17711 15530 17720
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15108 13932 15160 13938
rect 15028 13892 15108 13920
rect 15028 13258 15056 13892
rect 15108 13874 15160 13880
rect 15488 13870 15516 17711
rect 15580 16028 15608 21383
rect 15764 19122 15792 22578
rect 15856 21962 15884 22714
rect 15948 22030 15976 23559
rect 16028 22636 16080 22642
rect 16028 22578 16080 22584
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15844 21956 15896 21962
rect 15844 21898 15896 21904
rect 15856 21332 15884 21898
rect 15948 21554 15976 21966
rect 16040 21729 16068 22578
rect 16026 21720 16082 21729
rect 16026 21655 16082 21664
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 16028 21344 16080 21350
rect 15856 21304 16028 21332
rect 16028 21286 16080 21292
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 15936 20868 15988 20874
rect 15936 20810 15988 20816
rect 15856 20641 15884 20810
rect 15842 20632 15898 20641
rect 15842 20567 15898 20576
rect 15948 20505 15976 20810
rect 15934 20496 15990 20505
rect 15844 20460 15896 20466
rect 15934 20431 15990 20440
rect 15844 20402 15896 20408
rect 15856 19417 15884 20402
rect 15934 20360 15990 20369
rect 15934 20295 15990 20304
rect 15948 20262 15976 20295
rect 16040 20262 16068 21286
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16040 20074 16068 20198
rect 15948 20046 16068 20074
rect 15842 19408 15898 19417
rect 15842 19343 15898 19352
rect 15764 19094 15884 19122
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 15764 18426 15792 18906
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15672 17513 15700 17546
rect 15658 17504 15714 17513
rect 15658 17439 15714 17448
rect 15764 16182 15792 18362
rect 15856 17921 15884 19094
rect 15948 18222 15976 20046
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16040 18698 16068 19246
rect 16028 18692 16080 18698
rect 16028 18634 16080 18640
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15842 17912 15898 17921
rect 15842 17847 15898 17856
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15936 17740 15988 17746
rect 15936 17682 15988 17688
rect 15752 16176 15804 16182
rect 15752 16118 15804 16124
rect 15580 16000 15792 16028
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15658 13696 15714 13705
rect 15658 13631 15714 13640
rect 15106 13560 15162 13569
rect 15106 13495 15162 13504
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 14568 11898 14596 13194
rect 15028 12918 15056 13194
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 15028 12442 15056 12854
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 15028 11354 15056 12378
rect 15120 11898 15148 13495
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 15488 12306 15516 12718
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15580 11014 15608 12174
rect 15672 11898 15700 13631
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15764 11150 15792 16000
rect 15856 15638 15884 17682
rect 15948 17134 15976 17682
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 16040 16794 16068 18634
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 16132 14074 16160 23666
rect 16224 21978 16252 26302
rect 16316 26302 16450 26330
rect 16316 23322 16344 26302
rect 16394 26200 16450 26302
rect 16762 26200 16818 27000
rect 17130 26200 17186 27000
rect 17498 26200 17554 27000
rect 17866 26330 17922 27000
rect 17604 26302 17922 26330
rect 16396 24336 16448 24342
rect 16396 24278 16448 24284
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16224 21950 16344 21978
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16224 20330 16252 21830
rect 16316 21486 16344 21950
rect 16304 21480 16356 21486
rect 16304 21422 16356 21428
rect 16408 20369 16436 24278
rect 16578 24032 16634 24041
rect 16578 23967 16634 23976
rect 16592 22642 16620 23967
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16488 22500 16540 22506
rect 16488 22442 16540 22448
rect 16500 22166 16528 22442
rect 16684 22438 16712 22918
rect 16580 22432 16632 22438
rect 16580 22374 16632 22380
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16488 22160 16540 22166
rect 16592 22148 16620 22374
rect 16592 22120 16712 22148
rect 16488 22102 16540 22108
rect 16684 21894 16712 22120
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16488 21616 16540 21622
rect 16488 21558 16540 21564
rect 16500 20942 16528 21558
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16670 20496 16726 20505
rect 16488 20460 16540 20466
rect 16670 20431 16726 20440
rect 16488 20402 16540 20408
rect 16394 20360 16450 20369
rect 16212 20324 16264 20330
rect 16394 20295 16450 20304
rect 16212 20266 16264 20272
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16408 19990 16436 20198
rect 16500 20097 16528 20402
rect 16486 20088 16542 20097
rect 16486 20023 16542 20032
rect 16396 19984 16448 19990
rect 16396 19926 16448 19932
rect 16212 19780 16264 19786
rect 16212 19722 16264 19728
rect 16396 19780 16448 19786
rect 16396 19722 16448 19728
rect 16224 18873 16252 19722
rect 16304 19712 16356 19718
rect 16302 19680 16304 19689
rect 16356 19680 16358 19689
rect 16302 19615 16358 19624
rect 16408 19514 16436 19722
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16500 19378 16528 20023
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 19553 16620 19654
rect 16578 19544 16634 19553
rect 16578 19479 16634 19488
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 16210 18864 16266 18873
rect 16210 18799 16266 18808
rect 16212 18692 16264 18698
rect 16212 18634 16264 18640
rect 16224 18222 16252 18634
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16224 18086 16252 18158
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16224 17513 16252 18022
rect 16210 17504 16266 17513
rect 16210 17439 16266 17448
rect 16316 16969 16344 19110
rect 16408 17354 16436 19110
rect 16500 18834 16528 19314
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16578 18592 16634 18601
rect 16578 18527 16634 18536
rect 16486 18456 16542 18465
rect 16486 18391 16488 18400
rect 16540 18391 16542 18400
rect 16488 18362 16540 18368
rect 16592 18358 16620 18527
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 17882 16528 18022
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16408 17326 16528 17354
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16302 16960 16358 16969
rect 16302 16895 16358 16904
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 13530 16068 13670
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 16132 12170 16160 13126
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 16120 11280 16172 11286
rect 16118 11248 16120 11257
rect 16172 11248 16174 11257
rect 16118 11183 16174 11192
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15764 10810 15792 11086
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 16224 9450 16252 16050
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16316 15638 16344 15846
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16408 13394 16436 17206
rect 16500 15026 16528 17326
rect 16592 15434 16620 17682
rect 16684 16794 16712 20431
rect 16776 19310 16804 26200
rect 16856 24676 16908 24682
rect 16856 24618 16908 24624
rect 16868 23526 16896 24618
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 16960 24410 16988 24550
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16960 23526 16988 24006
rect 17038 23896 17094 23905
rect 17144 23882 17172 26200
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17144 23854 17264 23882
rect 17038 23831 17094 23840
rect 17052 23633 17080 23831
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17038 23624 17094 23633
rect 17038 23559 17094 23568
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16948 23248 17000 23254
rect 16948 23190 17000 23196
rect 16856 22976 16908 22982
rect 16960 22953 16988 23190
rect 17144 23186 17172 23666
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 17132 23044 17184 23050
rect 17132 22986 17184 22992
rect 16856 22918 16908 22924
rect 16946 22944 17002 22953
rect 16868 22545 16896 22918
rect 16946 22879 17002 22888
rect 16854 22536 16910 22545
rect 16854 22471 16910 22480
rect 17040 22228 17092 22234
rect 17040 22170 17092 22176
rect 17052 22098 17080 22170
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16868 18902 16896 21830
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16960 20777 16988 21422
rect 17052 21026 17080 21830
rect 17144 21418 17172 22986
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 17052 20998 17172 21026
rect 17040 20868 17092 20874
rect 17040 20810 17092 20816
rect 16946 20768 17002 20777
rect 16946 20703 17002 20712
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 16960 19854 16988 19994
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16856 18896 16908 18902
rect 16856 18838 16908 18844
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16776 15722 16804 18226
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16684 15694 16804 15722
rect 16868 15706 16896 16934
rect 16856 15700 16908 15706
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16500 14482 16528 14758
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16500 13394 16528 14418
rect 16592 14278 16620 15370
rect 16684 14890 16712 15694
rect 16856 15642 16908 15648
rect 16764 15632 16816 15638
rect 16764 15574 16816 15580
rect 16776 15094 16804 15574
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 16316 12170 16344 12854
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16304 12164 16356 12170
rect 16304 12106 16356 12112
rect 16408 11150 16436 12378
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16408 10810 16436 11086
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 16592 10198 16620 12786
rect 16960 11354 16988 17138
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16960 10810 16988 11086
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 17052 10606 17080 20810
rect 17144 19009 17172 20998
rect 17130 19000 17186 19009
rect 17236 18970 17264 23854
rect 17316 23792 17368 23798
rect 17316 23734 17368 23740
rect 17328 22094 17356 23734
rect 17420 23497 17448 24006
rect 17406 23488 17462 23497
rect 17406 23423 17462 23432
rect 17408 23180 17460 23186
rect 17408 23122 17460 23128
rect 17420 23050 17448 23122
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17328 22066 17448 22094
rect 17420 21554 17448 22066
rect 17512 21894 17540 26200
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 17408 21548 17460 21554
rect 17460 21508 17540 21536
rect 17408 21490 17460 21496
rect 17316 21412 17368 21418
rect 17316 21354 17368 21360
rect 17328 19310 17356 21354
rect 17406 21312 17462 21321
rect 17406 21247 17462 21256
rect 17420 21078 17448 21247
rect 17408 21072 17460 21078
rect 17408 21014 17460 21020
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 17130 18935 17186 18944
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17144 17882 17172 18566
rect 17236 18154 17264 18566
rect 17224 18148 17276 18154
rect 17224 18090 17276 18096
rect 17222 17912 17278 17921
rect 17132 17876 17184 17882
rect 17222 17847 17224 17856
rect 17132 17818 17184 17824
rect 17276 17847 17278 17856
rect 17224 17818 17276 17824
rect 17328 17814 17356 19246
rect 17316 17808 17368 17814
rect 17316 17750 17368 17756
rect 17222 17096 17278 17105
rect 17222 17031 17224 17040
rect 17276 17031 17278 17040
rect 17224 17002 17276 17008
rect 17132 16584 17184 16590
rect 17132 16526 17184 16532
rect 17144 14958 17172 16526
rect 17420 16522 17448 20742
rect 17512 18766 17540 21508
rect 17604 20806 17632 26302
rect 17866 26200 17922 26302
rect 18234 26330 18290 27000
rect 18234 26302 18368 26330
rect 18234 26200 18290 26302
rect 18052 24336 18104 24342
rect 17958 24304 18014 24313
rect 18236 24336 18288 24342
rect 18104 24296 18236 24324
rect 18052 24278 18104 24284
rect 18236 24278 18288 24284
rect 17958 24239 17960 24248
rect 18012 24239 18014 24248
rect 17960 24210 18012 24216
rect 17684 24064 17736 24070
rect 17684 24006 17736 24012
rect 17774 24032 17830 24041
rect 17696 23866 17724 24006
rect 17774 23967 17830 23976
rect 17684 23860 17736 23866
rect 17788 23848 17816 23967
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17788 23820 18092 23848
rect 17684 23802 17736 23808
rect 18064 23730 18092 23820
rect 17868 23724 17920 23730
rect 17868 23666 17920 23672
rect 18052 23724 18104 23730
rect 18052 23666 18104 23672
rect 17776 23588 17828 23594
rect 17776 23530 17828 23536
rect 17788 22574 17816 23530
rect 17880 23186 17908 23666
rect 17960 23316 18012 23322
rect 17960 23258 18012 23264
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 17972 23118 18000 23258
rect 18064 23118 18092 23666
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 18052 23112 18104 23118
rect 18052 23054 18104 23060
rect 17868 22976 17920 22982
rect 17868 22918 17920 22924
rect 17776 22568 17828 22574
rect 17776 22510 17828 22516
rect 17880 22250 17908 22918
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17788 22222 17908 22250
rect 17788 22166 17816 22222
rect 17776 22160 17828 22166
rect 17776 22102 17828 22108
rect 17868 22160 17920 22166
rect 17868 22102 17920 22108
rect 17880 21894 17908 22102
rect 18052 22094 18104 22098
rect 18052 22092 18276 22094
rect 18104 22066 18276 22092
rect 18052 22034 18104 22040
rect 18248 21894 18276 22066
rect 17684 21888 17736 21894
rect 17684 21830 17736 21836
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 17696 21690 17724 21830
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17682 21176 17738 21185
rect 17682 21111 17738 21120
rect 17880 21128 17908 21830
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 18340 21593 18368 26302
rect 18602 26200 18658 27000
rect 18970 26200 19026 27000
rect 19338 26200 19394 27000
rect 19706 26200 19762 27000
rect 20074 26330 20130 27000
rect 20442 26330 20498 27000
rect 20810 26330 20866 27000
rect 21178 26330 21234 27000
rect 19812 26302 20130 26330
rect 20180 26314 20498 26330
rect 19812 26217 19840 26302
rect 19798 26208 19854 26217
rect 18616 23225 18644 26200
rect 18984 24721 19012 26200
rect 18970 24712 19026 24721
rect 18970 24647 19026 24656
rect 19156 24404 19208 24410
rect 19156 24346 19208 24352
rect 18788 24268 18840 24274
rect 18788 24210 18840 24216
rect 18800 23662 18828 24210
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18602 23216 18658 23225
rect 18420 23180 18472 23186
rect 18602 23151 18658 23160
rect 18696 23180 18748 23186
rect 18420 23122 18472 23128
rect 18696 23122 18748 23128
rect 18432 22778 18460 23122
rect 18602 23080 18658 23089
rect 18512 23044 18564 23050
rect 18602 23015 18604 23024
rect 18512 22986 18564 22992
rect 18656 23015 18658 23024
rect 18604 22986 18656 22992
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 18524 22545 18552 22986
rect 18510 22536 18566 22545
rect 18510 22471 18566 22480
rect 18708 22409 18736 23122
rect 18694 22400 18750 22409
rect 18694 22335 18750 22344
rect 18786 22264 18842 22273
rect 18420 22228 18472 22234
rect 18786 22199 18842 22208
rect 18420 22170 18472 22176
rect 18326 21584 18382 21593
rect 18326 21519 18382 21528
rect 18432 21457 18460 22170
rect 18604 21956 18656 21962
rect 18604 21898 18656 21904
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 18418 21448 18474 21457
rect 18328 21412 18380 21418
rect 18418 21383 18474 21392
rect 18328 21354 18380 21360
rect 17960 21140 18012 21146
rect 17696 21078 17724 21111
rect 17880 21100 17960 21128
rect 17684 21072 17736 21078
rect 17684 21014 17736 21020
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17592 20596 17644 20602
rect 17592 20538 17644 20544
rect 17604 20058 17632 20538
rect 17696 20398 17724 20878
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17696 18834 17724 20334
rect 17880 19334 17908 21100
rect 17960 21082 18012 21088
rect 18340 21010 18368 21354
rect 18512 21140 18564 21146
rect 18512 21082 18564 21088
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18524 20534 18552 21082
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18512 19984 18564 19990
rect 18512 19926 18564 19932
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 18328 19372 18380 19378
rect 17880 19306 18000 19334
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 17776 18896 17828 18902
rect 17776 18838 17828 18844
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17500 18760 17552 18766
rect 17500 18702 17552 18708
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17696 18222 17724 18566
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17512 16697 17540 17478
rect 17498 16688 17554 16697
rect 17498 16623 17554 16632
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17236 15570 17264 16390
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17420 15450 17448 16458
rect 17500 15972 17552 15978
rect 17500 15914 17552 15920
rect 17328 15434 17448 15450
rect 17316 15428 17448 15434
rect 17368 15422 17448 15428
rect 17316 15370 17368 15376
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 17236 15094 17264 15302
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 17236 14346 17264 15030
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 17144 9518 17172 14010
rect 17236 13258 17264 14282
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 17236 12918 17264 13194
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17328 11354 17356 13670
rect 17420 12306 17448 13874
rect 17512 13530 17540 15914
rect 17604 14074 17632 18022
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17696 17270 17724 17478
rect 17684 17264 17736 17270
rect 17684 17206 17736 17212
rect 17696 16522 17724 17206
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17696 15434 17724 16458
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17682 14104 17738 14113
rect 17592 14068 17644 14074
rect 17682 14039 17738 14048
rect 17592 14010 17644 14016
rect 17696 14006 17724 14039
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17604 13190 17632 13738
rect 17788 13376 17816 18838
rect 17880 17678 17908 18906
rect 17972 18630 18000 19306
rect 18248 19320 18328 19334
rect 18248 19314 18380 19320
rect 18248 19306 18368 19314
rect 18052 18896 18104 18902
rect 18050 18864 18052 18873
rect 18104 18864 18106 18873
rect 18050 18799 18106 18808
rect 18248 18698 18276 19306
rect 18420 18896 18472 18902
rect 18420 18838 18472 18844
rect 18328 18828 18380 18834
rect 18328 18770 18380 18776
rect 18236 18692 18288 18698
rect 18236 18634 18288 18640
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18340 17202 18368 18770
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18142 17096 18198 17105
rect 18142 17031 18198 17040
rect 18326 17096 18382 17105
rect 18326 17031 18328 17040
rect 18156 16998 18184 17031
rect 18380 17031 18382 17040
rect 18328 17002 18380 17008
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17880 14006 17908 15846
rect 18432 15416 18460 18838
rect 18524 18834 18552 19926
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18524 18290 18552 18634
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18616 17626 18644 21898
rect 18708 21146 18736 21898
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18708 20602 18736 20946
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18708 19514 18736 19858
rect 18696 19508 18748 19514
rect 18696 19450 18748 19456
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18340 15388 18460 15416
rect 18524 17598 18644 17626
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17696 13348 17816 13376
rect 17592 13184 17644 13190
rect 17592 13126 17644 13132
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17512 12442 17540 12718
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17604 12102 17632 12854
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17500 11824 17552 11830
rect 17604 11812 17632 12038
rect 17552 11784 17632 11812
rect 17500 11766 17552 11772
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17696 10810 17724 13348
rect 17880 11218 17908 13398
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18340 12782 18368 15388
rect 18418 15328 18474 15337
rect 18418 15263 18474 15272
rect 18432 14385 18460 15263
rect 18418 14376 18474 14385
rect 18418 14311 18474 14320
rect 18524 13734 18552 17598
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 15638 18644 17478
rect 18604 15632 18656 15638
rect 18604 15574 18656 15580
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18616 14482 18644 14758
rect 18708 14550 18736 18158
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18708 13394 18736 14486
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18326 12608 18382 12617
rect 18326 12543 18382 12552
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 18340 10674 18368 12543
rect 18432 11218 18460 12786
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18616 11694 18644 12650
rect 18708 12322 18736 12718
rect 18800 12442 18828 22199
rect 18970 21992 19026 22001
rect 18970 21927 19026 21936
rect 18984 21894 19012 21927
rect 18880 21888 18932 21894
rect 18880 21830 18932 21836
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18892 21672 18920 21830
rect 18892 21644 19012 21672
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18892 15910 18920 21490
rect 18984 19990 19012 21644
rect 19168 21622 19196 24346
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19260 22778 19288 24006
rect 19352 23254 19380 26200
rect 19340 23248 19392 23254
rect 19340 23190 19392 23196
rect 19720 23168 19748 26200
rect 20074 26200 20130 26302
rect 20168 26308 20498 26314
rect 20220 26302 20498 26308
rect 20168 26250 20220 26256
rect 20442 26200 20498 26302
rect 20732 26302 20866 26330
rect 19798 26143 19854 26152
rect 20352 25016 20404 25022
rect 20352 24958 20404 24964
rect 19800 24064 19852 24070
rect 19800 24006 19852 24012
rect 19812 23526 19840 24006
rect 20260 23588 20312 23594
rect 20260 23530 20312 23536
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19628 23140 19748 23168
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19352 22030 19380 23054
rect 19628 22681 19656 23140
rect 19708 23044 19760 23050
rect 19708 22986 19760 22992
rect 19720 22710 19748 22986
rect 19812 22982 19840 23462
rect 19800 22976 19852 22982
rect 19800 22918 19852 22924
rect 19708 22704 19760 22710
rect 19614 22672 19670 22681
rect 19708 22646 19760 22652
rect 19614 22607 19670 22616
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 19432 22500 19484 22506
rect 19432 22442 19484 22448
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 19156 21616 19208 21622
rect 19156 21558 19208 21564
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 18972 19984 19024 19990
rect 18972 19926 19024 19932
rect 18984 17105 19012 19926
rect 19076 18834 19104 20810
rect 19156 20528 19208 20534
rect 19260 20505 19288 21490
rect 19352 21350 19380 21966
rect 19444 21962 19472 22442
rect 19432 21956 19484 21962
rect 19432 21898 19484 21904
rect 19524 21956 19576 21962
rect 19524 21898 19576 21904
rect 19444 21865 19472 21898
rect 19430 21856 19486 21865
rect 19430 21791 19486 21800
rect 19536 21729 19564 21898
rect 19522 21720 19578 21729
rect 19522 21655 19578 21664
rect 19812 21570 19840 22578
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19904 22166 19932 22510
rect 19892 22160 19944 22166
rect 19892 22102 19944 22108
rect 19444 21542 19840 21570
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 20942 19380 21286
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19156 20470 19208 20476
rect 19246 20496 19302 20505
rect 19168 20058 19196 20470
rect 19246 20431 19302 20440
rect 19248 20392 19300 20398
rect 19352 20380 19380 20878
rect 19300 20352 19380 20380
rect 19248 20334 19300 20340
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19168 19378 19196 19994
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19168 18426 19196 19110
rect 19260 18766 19288 20334
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19156 18420 19208 18426
rect 19156 18362 19208 18368
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 18970 17096 19026 17105
rect 18970 17031 19026 17040
rect 19168 16182 19196 18090
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19260 16454 19288 17070
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19156 16176 19208 16182
rect 19156 16118 19208 16124
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18984 15366 19012 15982
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18892 14906 18920 15098
rect 18984 15094 19012 15302
rect 18972 15088 19024 15094
rect 18972 15030 19024 15036
rect 18892 14890 19012 14906
rect 18892 14884 19024 14890
rect 18892 14878 18972 14884
rect 18972 14826 19024 14832
rect 19076 14822 19104 16050
rect 19154 15736 19210 15745
rect 19352 15706 19380 18090
rect 19444 16833 19472 21542
rect 19708 21480 19760 21486
rect 20180 21434 20208 22578
rect 20272 21894 20300 23530
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20272 21554 20300 21830
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 19708 21422 19760 21428
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19536 18290 19564 18634
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19430 16824 19486 16833
rect 19430 16759 19486 16768
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19444 16250 19472 16458
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19154 15671 19210 15680
rect 19340 15700 19392 15706
rect 19168 15162 19196 15671
rect 19340 15642 19392 15648
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 14657 19104 14758
rect 19062 14648 19118 14657
rect 18972 14612 19024 14618
rect 19062 14583 19118 14592
rect 19248 14612 19300 14618
rect 18972 14554 19024 14560
rect 19248 14554 19300 14560
rect 18984 14498 19012 14554
rect 19260 14498 19288 14554
rect 18984 14470 19288 14498
rect 19156 14408 19208 14414
rect 18970 14376 19026 14385
rect 18970 14311 19026 14320
rect 19076 14368 19156 14396
rect 18880 14272 18932 14278
rect 18878 14240 18880 14249
rect 18932 14240 18934 14249
rect 18878 14175 18934 14184
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18892 12918 18920 13262
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18708 12294 18828 12322
rect 18694 12200 18750 12209
rect 18694 12135 18696 12144
rect 18748 12135 18750 12144
rect 18696 12106 18748 12112
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 18800 11558 18828 12294
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18892 12102 18920 12242
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18880 11824 18932 11830
rect 18880 11766 18932 11772
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18420 11212 18472 11218
rect 18420 11154 18472 11160
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18340 10266 18368 10610
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 18064 9178 18092 9318
rect 14464 9172 14516 9178
rect 14464 9114 14516 9120
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 15106 8392 15162 8401
rect 15106 8327 15162 8336
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 15120 8022 15148 8327
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 18708 7886 18736 11290
rect 18892 10674 18920 11766
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18984 4078 19012 14311
rect 19076 14006 19104 14368
rect 19156 14350 19208 14356
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19168 13462 19196 14214
rect 19352 14074 19380 14894
rect 19628 14618 19656 19654
rect 19720 19378 19748 21422
rect 19812 21406 20208 21434
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19708 19236 19760 19242
rect 19708 19178 19760 19184
rect 19720 19009 19748 19178
rect 19706 19000 19762 19009
rect 19706 18935 19762 18944
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19720 18057 19748 18158
rect 19706 18048 19762 18057
rect 19706 17983 19762 17992
rect 19812 17921 19840 21406
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19892 20392 19944 20398
rect 19892 20334 19944 20340
rect 19904 19446 19932 20334
rect 19892 19440 19944 19446
rect 19892 19382 19944 19388
rect 19904 19310 19932 19382
rect 19892 19304 19944 19310
rect 19892 19246 19944 19252
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19798 17912 19854 17921
rect 19798 17847 19854 17856
rect 19798 17776 19854 17785
rect 19798 17711 19800 17720
rect 19852 17711 19854 17720
rect 19800 17682 19852 17688
rect 19708 17536 19760 17542
rect 19760 17496 19840 17524
rect 19708 17478 19760 17484
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19720 16522 19748 17002
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19616 14340 19668 14346
rect 19616 14282 19668 14288
rect 19628 14249 19656 14282
rect 19614 14240 19670 14249
rect 19614 14175 19670 14184
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19156 13456 19208 13462
rect 19156 13398 19208 13404
rect 19062 13288 19118 13297
rect 19062 13223 19118 13232
rect 19076 13190 19104 13223
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19168 12646 19196 12718
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19076 8430 19104 12582
rect 19352 12238 19380 14010
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19444 13462 19472 13942
rect 19720 13530 19748 16050
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19248 12164 19300 12170
rect 19248 12106 19300 12112
rect 19260 11286 19288 12106
rect 19352 11898 19380 12174
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19444 11762 19472 13262
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19536 12782 19564 13126
rect 19812 12782 19840 17496
rect 19904 14346 19932 18022
rect 19996 15502 20024 21286
rect 20272 21162 20300 21490
rect 20180 21134 20300 21162
rect 20076 19780 20128 19786
rect 20076 19722 20128 19728
rect 20088 17338 20116 19722
rect 20180 17542 20208 21134
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20272 20602 20300 20810
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20272 20058 20300 20538
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 20272 18358 20300 18634
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 20076 17128 20128 17134
rect 20076 17070 20128 17076
rect 20088 16250 20116 17070
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 20180 16114 20208 16458
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20076 15972 20128 15978
rect 20076 15914 20128 15920
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 20088 14521 20116 15914
rect 20166 15736 20222 15745
rect 20166 15671 20222 15680
rect 20074 14512 20130 14521
rect 20074 14447 20130 14456
rect 19892 14340 19944 14346
rect 19892 14282 19944 14288
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19432 11756 19484 11762
rect 19432 11698 19484 11704
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19352 10742 19380 11630
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19430 10296 19486 10305
rect 19430 10231 19432 10240
rect 19484 10231 19486 10240
rect 19432 10202 19484 10208
rect 19246 10024 19302 10033
rect 19246 9959 19302 9968
rect 19064 8424 19116 8430
rect 19064 8366 19116 8372
rect 19260 8362 19288 9959
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19352 9110 19380 9590
rect 19430 9480 19486 9489
rect 19430 9415 19432 9424
rect 19484 9415 19486 9424
rect 19432 9386 19484 9392
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 19536 3074 19564 12038
rect 19720 11558 19748 12242
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11830 19840 12038
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19812 11354 19840 11494
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19616 11280 19668 11286
rect 19616 11222 19668 11228
rect 19628 10062 19656 11222
rect 19706 11112 19762 11121
rect 19706 11047 19708 11056
rect 19760 11047 19762 11056
rect 19708 11018 19760 11024
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19904 8634 19932 12378
rect 19996 10674 20024 14282
rect 20180 12434 20208 15671
rect 20272 13002 20300 17682
rect 20364 17354 20392 24958
rect 20732 23746 20760 26302
rect 20810 26200 20866 26302
rect 21008 26302 21234 26330
rect 21272 26376 21324 26382
rect 21546 26330 21602 27000
rect 21324 26324 21602 26330
rect 21272 26318 21602 26324
rect 21284 26302 21602 26318
rect 20812 24200 20864 24206
rect 20812 24142 20864 24148
rect 20824 23798 20852 24142
rect 20904 24132 20956 24138
rect 20904 24074 20956 24080
rect 20640 23718 20760 23746
rect 20812 23792 20864 23798
rect 20812 23734 20864 23740
rect 20640 23361 20668 23718
rect 20720 23656 20772 23662
rect 20720 23598 20772 23604
rect 20626 23352 20682 23361
rect 20626 23287 20682 23296
rect 20732 23254 20760 23598
rect 20720 23248 20772 23254
rect 20720 23190 20772 23196
rect 20824 23118 20852 23734
rect 20916 23662 20944 24074
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20812 23112 20864 23118
rect 20916 23089 20944 23598
rect 21008 23186 21036 26302
rect 21178 26200 21234 26302
rect 21546 26200 21602 26302
rect 21914 26200 21970 27000
rect 22190 26344 22246 26353
rect 22190 26279 22246 26288
rect 21732 24336 21784 24342
rect 21732 24278 21784 24284
rect 21744 23594 21772 24278
rect 21928 24177 21956 26200
rect 22204 26058 22232 26279
rect 22282 26200 22338 27000
rect 22650 26330 22706 27000
rect 23018 26330 23074 27000
rect 23386 26330 23442 27000
rect 24490 26330 24546 27000
rect 22388 26302 22706 26330
rect 22296 26058 22324 26200
rect 22204 26030 22324 26058
rect 22006 25664 22062 25673
rect 22006 25599 22062 25608
rect 22020 24410 22048 25599
rect 22008 24404 22060 24410
rect 22008 24346 22060 24352
rect 21914 24168 21970 24177
rect 21914 24103 21970 24112
rect 22020 23730 22048 24346
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22296 23662 22324 24142
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 21732 23588 21784 23594
rect 21732 23530 21784 23536
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 20996 23180 21048 23186
rect 20996 23122 21048 23128
rect 21272 23112 21324 23118
rect 20812 23054 20864 23060
rect 20902 23080 20958 23089
rect 21272 23054 21324 23060
rect 20902 23015 20958 23024
rect 21284 22778 21312 23054
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 20444 22704 20496 22710
rect 20444 22646 20496 22652
rect 20456 21146 20484 22646
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20364 17326 20484 17354
rect 20456 16250 20484 17326
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20548 16130 20576 22714
rect 20812 22432 20864 22438
rect 20812 22374 20864 22380
rect 20720 22094 20772 22098
rect 20824 22094 20852 22374
rect 21284 22094 21312 22714
rect 21652 22556 21680 23462
rect 22296 23186 22324 23598
rect 22388 23497 22416 26302
rect 22650 26200 22706 26302
rect 22756 26302 23074 26330
rect 22756 24290 22784 26302
rect 23018 26200 23074 26302
rect 23124 26302 23442 26330
rect 23124 24664 23152 26302
rect 23386 26200 23442 26302
rect 24320 26302 24546 26330
rect 23478 26072 23534 26081
rect 23478 26007 23534 26016
rect 23388 24744 23440 24750
rect 23388 24686 23440 24692
rect 22480 24262 22784 24290
rect 22848 24636 23152 24664
rect 22374 23488 22430 23497
rect 22374 23423 22430 23432
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 21652 22528 21864 22556
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21376 22273 21404 22374
rect 21362 22264 21418 22273
rect 21362 22199 21418 22208
rect 20720 22092 20852 22094
rect 20772 22066 20852 22092
rect 20720 22034 20772 22040
rect 20824 20602 20852 22066
rect 21192 22066 21312 22094
rect 21730 22128 21786 22137
rect 21192 21962 21220 22066
rect 21730 22063 21786 22072
rect 21546 21992 21602 22001
rect 21180 21956 21232 21962
rect 21546 21927 21602 21936
rect 21180 21898 21232 21904
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20718 20360 20774 20369
rect 20718 20295 20774 20304
rect 20732 18970 20760 20295
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20824 19718 20852 20198
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20916 18698 20944 20946
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 21008 19825 21036 20810
rect 21100 20806 21128 21626
rect 21088 20800 21140 20806
rect 21088 20742 21140 20748
rect 21192 20262 21220 21898
rect 21454 21856 21510 21865
rect 21454 21791 21510 21800
rect 21468 21486 21496 21791
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 21456 21480 21508 21486
rect 21456 21422 21508 21428
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21192 20074 21220 20198
rect 21100 20058 21220 20074
rect 21088 20052 21220 20058
rect 21140 20046 21220 20052
rect 21088 19994 21140 20000
rect 20994 19816 21050 19825
rect 20994 19751 21050 19760
rect 20996 19440 21048 19446
rect 20996 19382 21048 19388
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 21008 18442 21036 19382
rect 21100 19174 21128 19994
rect 21178 19544 21234 19553
rect 21178 19479 21234 19488
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 21100 18698 21128 19110
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 20824 18414 21036 18442
rect 20824 18306 20852 18414
rect 20904 18352 20956 18358
rect 20732 18278 20852 18306
rect 20902 18320 20904 18329
rect 20956 18320 20958 18329
rect 20732 18154 20760 18278
rect 20902 18255 20958 18264
rect 21008 18170 21036 18414
rect 21100 18222 21128 18634
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20812 18148 20864 18154
rect 20812 18090 20864 18096
rect 20916 18142 21036 18170
rect 21088 18216 21140 18222
rect 21088 18158 21140 18164
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 20640 16998 20668 17818
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20456 16102 20576 16130
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20364 14074 20392 14554
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20272 12974 20392 13002
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20088 12406 20208 12434
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 20088 9654 20116 12406
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 8634 20024 9318
rect 19892 8628 19944 8634
rect 19892 8570 19944 8576
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20272 7410 20300 12582
rect 20364 12306 20392 12974
rect 20352 12300 20404 12306
rect 20352 12242 20404 12248
rect 20456 11150 20484 16102
rect 20536 15904 20588 15910
rect 20536 15846 20588 15852
rect 20548 15706 20576 15846
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20548 11234 20576 15302
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20640 13530 20668 14010
rect 20732 13938 20760 14826
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20720 13728 20772 13734
rect 20720 13670 20772 13676
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20640 13258 20668 13466
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20640 12102 20668 12650
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20548 11206 20668 11234
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20260 7404 20312 7410
rect 20260 7346 20312 7352
rect 20168 4072 20220 4078
rect 20168 4014 20220 4020
rect 19536 3058 19656 3074
rect 19536 3052 19668 3058
rect 19536 3046 19616 3052
rect 19616 2994 19668 3000
rect 19524 2984 19576 2990
rect 19524 2926 19576 2932
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 19536 2650 19564 2926
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 6920 2440 6972 2446
rect 6748 2388 6920 2394
rect 6748 2382 6972 2388
rect 6748 2366 6960 2382
rect 6748 800 6776 2366
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 20180 800 20208 4014
rect 20548 3534 20576 11018
rect 20640 9042 20668 11206
rect 20732 10674 20760 13670
rect 20824 13190 20852 18090
rect 20916 16182 20944 18142
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 20904 14544 20956 14550
rect 20904 14486 20956 14492
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20718 10432 20774 10441
rect 20718 10367 20774 10376
rect 20732 10266 20760 10367
rect 20720 10260 20772 10266
rect 20720 10202 20772 10208
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9654 20760 9998
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20824 9586 20852 11290
rect 20916 11150 20944 14486
rect 21008 13870 21036 18022
rect 21100 17610 21128 18158
rect 21088 17604 21140 17610
rect 21088 17546 21140 17552
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 21100 17202 21128 17274
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 21008 11558 21036 11766
rect 21100 11626 21128 15982
rect 21192 15570 21220 19479
rect 21284 17134 21312 21422
rect 21560 20505 21588 21927
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21546 20496 21602 20505
rect 21546 20431 21602 20440
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 21364 19780 21416 19786
rect 21364 19722 21416 19728
rect 21376 19446 21404 19722
rect 21364 19440 21416 19446
rect 21364 19382 21416 19388
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21376 18290 21404 18906
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21468 17728 21496 20334
rect 21548 20324 21600 20330
rect 21548 20266 21600 20272
rect 21560 19310 21588 20266
rect 21548 19304 21600 19310
rect 21548 19246 21600 19252
rect 21376 17700 21496 17728
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 15570 21312 16390
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21272 15564 21324 15570
rect 21272 15506 21324 15512
rect 21376 15450 21404 17700
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21468 17134 21496 17546
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21652 16538 21680 20742
rect 21744 19174 21772 22063
rect 21836 21010 21864 22528
rect 22020 21894 22048 22986
rect 22192 22568 22244 22574
rect 22190 22536 22192 22545
rect 22284 22568 22336 22574
rect 22244 22536 22246 22545
rect 22284 22510 22336 22516
rect 22190 22471 22246 22480
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 21928 21146 21956 21490
rect 21916 21140 21968 21146
rect 21916 21082 21968 21088
rect 22020 21078 22048 21830
rect 22008 21072 22060 21078
rect 22008 21014 22060 21020
rect 21824 21004 21876 21010
rect 21824 20946 21876 20952
rect 21916 21004 21968 21010
rect 21916 20946 21968 20952
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21836 19786 21864 20198
rect 21928 20058 21956 20946
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 21824 19780 21876 19786
rect 21824 19722 21876 19728
rect 21822 19544 21878 19553
rect 21822 19479 21824 19488
rect 21876 19479 21878 19488
rect 21824 19450 21876 19456
rect 21824 19236 21876 19242
rect 21824 19178 21876 19184
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21836 17338 21864 19178
rect 21928 18834 21956 19994
rect 22006 19544 22062 19553
rect 22006 19479 22062 19488
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 21928 18290 21956 18634
rect 22020 18630 22048 19479
rect 22112 19145 22140 21966
rect 22192 21548 22244 21554
rect 22192 21490 22244 21496
rect 22204 20777 22232 21490
rect 22190 20768 22246 20777
rect 22190 20703 22246 20712
rect 22192 20528 22244 20534
rect 22192 20470 22244 20476
rect 22204 19553 22232 20470
rect 22296 20330 22324 22510
rect 22480 22030 22508 24262
rect 22652 24132 22704 24138
rect 22652 24074 22704 24080
rect 22664 23662 22692 24074
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22652 23656 22704 23662
rect 22652 23598 22704 23604
rect 22572 22982 22600 23598
rect 22848 23338 22876 24636
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23216 24070 23244 24210
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23400 23769 23428 24686
rect 23386 23760 23442 23769
rect 23386 23695 23442 23704
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22756 23310 22876 23338
rect 22650 23080 22706 23089
rect 22650 23015 22706 23024
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22374 21584 22430 21593
rect 22374 21519 22430 21528
rect 22388 20398 22416 21519
rect 22466 21448 22522 21457
rect 22466 21383 22522 21392
rect 22376 20392 22428 20398
rect 22376 20334 22428 20340
rect 22284 20324 22336 20330
rect 22284 20266 22336 20272
rect 22480 19768 22508 21383
rect 22664 21332 22692 23015
rect 22756 22438 22784 23310
rect 23388 23248 23440 23254
rect 22834 23216 22890 23225
rect 23388 23190 23440 23196
rect 22834 23151 22890 23160
rect 23296 23180 23348 23186
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 22848 22234 22876 23151
rect 23296 23122 23348 23128
rect 23204 23112 23256 23118
rect 23204 23054 23256 23060
rect 23216 22506 23244 23054
rect 23308 22642 23336 23122
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 23204 22500 23256 22506
rect 23204 22442 23256 22448
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 23204 22228 23256 22234
rect 23204 22170 23256 22176
rect 23216 22030 23244 22170
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 22756 21622 22784 21966
rect 22744 21616 22796 21622
rect 22744 21558 22796 21564
rect 22572 21304 22692 21332
rect 22572 20534 22600 21304
rect 22756 21146 22784 21558
rect 23308 21554 23336 22578
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22744 21140 22796 21146
rect 22744 21082 22796 21088
rect 22664 20992 22692 21082
rect 22664 20964 22784 20992
rect 22650 20904 22706 20913
rect 22650 20839 22652 20848
rect 22704 20839 22706 20848
rect 22652 20810 22704 20816
rect 22756 20534 22784 20964
rect 22836 20800 22888 20806
rect 22836 20742 22888 20748
rect 22560 20528 22612 20534
rect 22560 20470 22612 20476
rect 22744 20528 22796 20534
rect 22744 20470 22796 20476
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22652 20392 22704 20398
rect 22652 20334 22704 20340
rect 22572 19961 22600 20334
rect 22558 19952 22614 19961
rect 22558 19887 22614 19896
rect 22480 19740 22600 19768
rect 22466 19680 22522 19689
rect 22466 19615 22522 19624
rect 22190 19544 22246 19553
rect 22480 19514 22508 19615
rect 22190 19479 22192 19488
rect 22244 19479 22246 19488
rect 22468 19508 22520 19514
rect 22192 19450 22244 19456
rect 22468 19450 22520 19456
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22098 19136 22154 19145
rect 22098 19071 22154 19080
rect 22296 18902 22324 19314
rect 22284 18896 22336 18902
rect 22284 18838 22336 18844
rect 22008 18624 22060 18630
rect 22376 18624 22428 18630
rect 22008 18566 22060 18572
rect 22282 18592 22338 18601
rect 22376 18566 22428 18572
rect 22282 18527 22338 18536
rect 21916 18284 21968 18290
rect 21916 18226 21968 18232
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21652 16510 21772 16538
rect 21640 16448 21692 16454
rect 21640 16390 21692 16396
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21284 15422 21404 15450
rect 21180 14884 21232 14890
rect 21180 14826 21232 14832
rect 21192 14074 21220 14826
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21192 12782 21220 13466
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21192 11762 21220 12718
rect 21284 11898 21312 15422
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21376 12434 21404 15302
rect 21468 15094 21496 16050
rect 21652 15434 21680 16390
rect 21744 16046 21772 16510
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21640 15428 21692 15434
rect 21640 15370 21692 15376
rect 21456 15088 21508 15094
rect 21456 15030 21508 15036
rect 21468 14618 21496 15030
rect 21836 14958 21864 17274
rect 21914 16688 21970 16697
rect 21914 16623 21970 16632
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21546 14512 21602 14521
rect 21546 14447 21602 14456
rect 21456 13864 21508 13870
rect 21456 13806 21508 13812
rect 21468 13530 21496 13806
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21560 12918 21588 14447
rect 21928 14006 21956 16623
rect 22020 14414 22048 18226
rect 22192 17808 22244 17814
rect 22192 17750 22244 17756
rect 22098 17504 22154 17513
rect 22098 17439 22154 17448
rect 22112 17270 22140 17439
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 22204 17066 22232 17750
rect 22296 17542 22324 18527
rect 22388 17882 22416 18566
rect 22572 17898 22600 19740
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22480 17870 22600 17898
rect 22664 17882 22692 20334
rect 22742 19952 22798 19961
rect 22742 19887 22798 19896
rect 22756 19009 22784 19887
rect 22848 19281 22876 20742
rect 23308 20466 23336 21490
rect 23400 20874 23428 23190
rect 23492 22234 23520 26007
rect 23846 24440 23902 24449
rect 24320 24410 24348 26302
rect 24490 26200 24546 26302
rect 24858 26200 24914 27000
rect 25042 26480 25098 26489
rect 25042 26415 25098 26424
rect 24766 25256 24822 25265
rect 24766 25191 24822 25200
rect 24398 24984 24454 24993
rect 24398 24919 24454 24928
rect 24412 24410 24440 24919
rect 23846 24375 23902 24384
rect 24308 24404 24360 24410
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23584 23866 23612 24006
rect 23572 23860 23624 23866
rect 23572 23802 23624 23808
rect 23584 22710 23612 23802
rect 23860 23633 23888 24375
rect 24308 24346 24360 24352
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 23940 24132 23992 24138
rect 23940 24074 23992 24080
rect 23952 23798 23980 24074
rect 24320 23866 24348 24346
rect 24412 24206 24440 24346
rect 24400 24200 24452 24206
rect 24400 24142 24452 24148
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24308 23860 24360 23866
rect 24308 23802 24360 23808
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 23846 23624 23902 23633
rect 23846 23559 23902 23568
rect 24504 23322 24532 24006
rect 24780 23798 24808 25191
rect 24860 24676 24912 24682
rect 24860 24618 24912 24624
rect 24584 23792 24636 23798
rect 24584 23734 24636 23740
rect 24768 23792 24820 23798
rect 24768 23734 24820 23740
rect 24596 23526 24624 23734
rect 24584 23520 24636 23526
rect 24584 23462 24636 23468
rect 24492 23316 24544 23322
rect 24492 23258 24544 23264
rect 23664 23044 23716 23050
rect 23664 22986 23716 22992
rect 23676 22778 23704 22986
rect 24032 22976 24084 22982
rect 24032 22918 24084 22924
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23572 22704 23624 22710
rect 23572 22646 23624 22652
rect 23480 22228 23532 22234
rect 23480 22170 23532 22176
rect 23480 22092 23532 22098
rect 23480 22034 23532 22040
rect 23492 20942 23520 22034
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23388 20868 23440 20874
rect 23388 20810 23440 20816
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23308 19922 23336 20402
rect 23296 19916 23348 19922
rect 23296 19858 23348 19864
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 22940 19378 22968 19790
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 23112 19712 23164 19718
rect 23112 19654 23164 19660
rect 23032 19553 23060 19654
rect 23018 19544 23074 19553
rect 23018 19479 23074 19488
rect 23124 19417 23152 19654
rect 23110 19408 23166 19417
rect 22928 19372 22980 19378
rect 23308 19378 23336 19858
rect 23492 19718 23520 20878
rect 23584 19990 23612 22646
rect 23676 21622 23704 22714
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23676 20874 23704 21558
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23664 20868 23716 20874
rect 23664 20810 23716 20816
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23572 19984 23624 19990
rect 23572 19926 23624 19932
rect 23388 19712 23440 19718
rect 23388 19654 23440 19660
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23110 19343 23166 19352
rect 23296 19372 23348 19378
rect 22928 19314 22980 19320
rect 23296 19314 23348 19320
rect 22834 19272 22890 19281
rect 22834 19207 22890 19216
rect 22940 19156 22968 19314
rect 22848 19128 22968 19156
rect 22742 19000 22798 19009
rect 22848 18970 22876 19128
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22742 18935 22798 18944
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 23020 18964 23072 18970
rect 23020 18906 23072 18912
rect 23032 18850 23060 18906
rect 22836 18828 22888 18834
rect 22836 18770 22888 18776
rect 22940 18822 23060 18850
rect 22652 17876 22704 17882
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22388 17066 22416 17818
rect 22480 17377 22508 17870
rect 22652 17818 22704 17824
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22466 17368 22522 17377
rect 22466 17303 22522 17312
rect 22572 17202 22600 17682
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22466 17096 22522 17105
rect 22192 17060 22244 17066
rect 22192 17002 22244 17008
rect 22376 17060 22428 17066
rect 22466 17031 22522 17040
rect 22560 17060 22612 17066
rect 22376 17002 22428 17008
rect 22098 16960 22154 16969
rect 22098 16895 22154 16904
rect 22112 15094 22140 16895
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22204 15026 22232 16730
rect 22284 16652 22336 16658
rect 22284 16594 22336 16600
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22296 14958 22324 16594
rect 22376 15904 22428 15910
rect 22376 15846 22428 15852
rect 22284 14952 22336 14958
rect 22284 14894 22336 14900
rect 22296 14618 22324 14894
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 21916 14000 21968 14006
rect 21916 13942 21968 13948
rect 22098 13968 22154 13977
rect 22296 13938 22324 14554
rect 22098 13903 22100 13912
rect 22152 13903 22154 13912
rect 22284 13932 22336 13938
rect 22100 13874 22152 13880
rect 22284 13874 22336 13880
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21548 12912 21600 12918
rect 21548 12854 21600 12860
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 21376 12406 21496 12434
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 21088 11620 21140 11626
rect 21088 11562 21140 11568
rect 20996 11552 21048 11558
rect 20996 11494 21048 11500
rect 20994 11384 21050 11393
rect 20994 11319 21050 11328
rect 21008 11286 21036 11319
rect 20996 11280 21048 11286
rect 20996 11222 21048 11228
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 21284 11082 21312 11834
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21088 10736 21140 10742
rect 21088 10678 21140 10684
rect 20812 9580 20864 9586
rect 20812 9522 20864 9528
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20916 9382 20944 9522
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20628 9036 20680 9042
rect 20628 8978 20680 8984
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20732 7478 20760 7686
rect 20720 7472 20772 7478
rect 20720 7414 20772 7420
rect 20916 5302 20944 8910
rect 21100 7410 21128 10678
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 21192 6798 21220 10406
rect 21284 10130 21312 10406
rect 21376 10130 21404 12242
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 21364 10124 21416 10130
rect 21364 10066 21416 10072
rect 21468 8974 21496 12406
rect 21652 12238 21680 12786
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21560 11762 21588 12106
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21560 11150 21588 11698
rect 21640 11620 21692 11626
rect 21640 11562 21692 11568
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 21560 9586 21588 11086
rect 21652 10266 21680 11562
rect 21744 11218 21772 13466
rect 21732 11212 21784 11218
rect 21732 11154 21784 11160
rect 21732 11076 21784 11082
rect 21732 11018 21784 11024
rect 21640 10260 21692 10266
rect 21640 10202 21692 10208
rect 21744 9994 21772 11018
rect 21836 10418 21864 13806
rect 22296 13394 22324 13874
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 22284 13388 22336 13394
rect 22284 13330 22336 13336
rect 21928 12850 21956 13330
rect 22282 13152 22338 13161
rect 22282 13087 22338 13096
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21928 12306 21956 12786
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22020 11694 22048 12378
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 21928 10742 21956 10950
rect 21916 10736 21968 10742
rect 21916 10678 21968 10684
rect 22112 10674 22140 12922
rect 22296 12918 22324 13087
rect 22284 12912 22336 12918
rect 22190 12880 22246 12889
rect 22284 12854 22336 12860
rect 22190 12815 22246 12824
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 21836 10390 22048 10418
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 21744 9722 21772 9930
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 21548 9580 21600 9586
rect 21548 9522 21600 9528
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21836 5710 21864 10202
rect 21916 9988 21968 9994
rect 21916 9930 21968 9936
rect 21928 9586 21956 9930
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 22020 8616 22048 10390
rect 21928 8588 22048 8616
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 20904 5296 20956 5302
rect 20904 5238 20956 5244
rect 21928 4146 21956 8588
rect 22204 8514 22232 12815
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22296 12442 22324 12718
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22282 12336 22338 12345
rect 22282 12271 22338 12280
rect 22296 9518 22324 12271
rect 22388 11150 22416 15846
rect 22480 15473 22508 17031
rect 22560 17002 22612 17008
rect 22572 16046 22600 17002
rect 22664 16658 22692 17818
rect 22744 17604 22796 17610
rect 22744 17546 22796 17552
rect 22756 17338 22784 17546
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22744 15972 22796 15978
rect 22744 15914 22796 15920
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22466 15464 22522 15473
rect 22466 15399 22522 15408
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22480 14618 22508 15098
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22468 13252 22520 13258
rect 22468 13194 22520 13200
rect 22480 12986 22508 13194
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22466 12880 22522 12889
rect 22466 12815 22522 12824
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22480 10690 22508 12815
rect 22572 10810 22600 15846
rect 22756 15434 22784 15914
rect 22848 15450 22876 18770
rect 22940 18698 22968 18822
rect 23018 18728 23074 18737
rect 22928 18692 22980 18698
rect 23018 18663 23020 18672
rect 22928 18634 22980 18640
rect 23072 18663 23074 18672
rect 23020 18634 23072 18640
rect 23308 18426 23336 19314
rect 23400 19258 23428 19654
rect 23400 19230 23520 19258
rect 23388 19168 23440 19174
rect 23386 19136 23388 19145
rect 23440 19136 23442 19145
rect 23386 19071 23442 19080
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23112 18352 23164 18358
rect 23110 18320 23112 18329
rect 23164 18320 23166 18329
rect 23110 18255 23166 18264
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23018 17776 23074 17785
rect 23308 17746 23336 18362
rect 23492 18170 23520 19230
rect 23400 18142 23520 18170
rect 23018 17711 23074 17720
rect 23296 17740 23348 17746
rect 22928 17536 22980 17542
rect 22928 17478 22980 17484
rect 22940 17270 22968 17478
rect 22928 17264 22980 17270
rect 22928 17206 22980 17212
rect 22940 16998 22968 17206
rect 23032 17105 23060 17711
rect 23296 17682 23348 17688
rect 23204 17672 23256 17678
rect 23204 17614 23256 17620
rect 23018 17096 23074 17105
rect 23216 17082 23244 17614
rect 23216 17054 23336 17082
rect 23018 17031 23074 17040
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23308 16794 23336 17054
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 23308 15978 23336 16390
rect 23296 15972 23348 15978
rect 23296 15914 23348 15920
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 22744 15428 22796 15434
rect 22848 15422 22968 15450
rect 22744 15370 22796 15376
rect 22836 15360 22888 15366
rect 22834 15328 22836 15337
rect 22888 15328 22890 15337
rect 22834 15263 22890 15272
rect 22742 15056 22798 15065
rect 22742 14991 22798 15000
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22664 12434 22692 14758
rect 22756 14278 22784 14991
rect 22940 14906 22968 15422
rect 23308 15162 23336 15914
rect 23296 15156 23348 15162
rect 23296 15098 23348 15104
rect 22848 14878 22968 14906
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22742 13832 22798 13841
rect 22742 13767 22798 13776
rect 22756 13394 22784 13767
rect 22744 13388 22796 13394
rect 22744 13330 22796 13336
rect 22744 13252 22796 13258
rect 22744 13194 22796 13200
rect 22756 13161 22784 13194
rect 22742 13152 22798 13161
rect 22742 13087 22798 13096
rect 22848 12866 22876 14878
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23400 14482 23428 18142
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23492 17814 23520 18022
rect 23480 17808 23532 17814
rect 23480 17750 23532 17756
rect 23480 17604 23532 17610
rect 23480 17546 23532 17552
rect 23492 16289 23520 17546
rect 23572 17536 23624 17542
rect 23572 17478 23624 17484
rect 23478 16280 23534 16289
rect 23478 16215 23534 16224
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23294 14240 23350 14249
rect 23294 14175 23350 14184
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22928 13388 22980 13394
rect 22928 13330 22980 13336
rect 22756 12838 22876 12866
rect 22756 12782 22784 12838
rect 22744 12776 22796 12782
rect 22940 12730 22968 13330
rect 22744 12718 22796 12724
rect 22848 12702 22968 12730
rect 22664 12406 22784 12434
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22388 10662 22508 10690
rect 22284 9512 22336 9518
rect 22284 9454 22336 9460
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22020 8498 22232 8514
rect 22008 8492 22232 8498
rect 22060 8486 22232 8492
rect 22008 8434 22060 8440
rect 22006 7032 22062 7041
rect 22006 6967 22062 6976
rect 22020 5914 22048 6967
rect 22296 6322 22324 9114
rect 22388 8634 22416 10662
rect 22468 10532 22520 10538
rect 22468 10474 22520 10480
rect 22480 9586 22508 10474
rect 22468 9580 22520 9586
rect 22468 9522 22520 9528
rect 22468 9444 22520 9450
rect 22468 9386 22520 9392
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22388 7886 22416 8570
rect 22480 8498 22508 9386
rect 22664 9110 22692 11086
rect 22652 9104 22704 9110
rect 22652 9046 22704 9052
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22664 7546 22692 8910
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22284 6316 22336 6322
rect 22284 6258 22336 6264
rect 22008 5908 22060 5914
rect 22008 5850 22060 5856
rect 22376 5772 22428 5778
rect 22376 5714 22428 5720
rect 22388 4826 22416 5714
rect 22650 5536 22706 5545
rect 22650 5471 22706 5480
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22664 4622 22692 5471
rect 22756 5234 22784 12406
rect 22848 11082 22876 12702
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23308 12434 23336 14175
rect 23386 13424 23442 13433
rect 23386 13359 23442 13368
rect 23400 12646 23428 13359
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23308 12406 23428 12434
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22836 11076 22888 11082
rect 22836 11018 22888 11024
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22836 10192 22888 10198
rect 22836 10134 22888 10140
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 21916 4140 21968 4146
rect 21916 4082 21968 4088
rect 22100 4004 22152 4010
rect 22100 3946 22152 3952
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 22008 3460 22060 3466
rect 22008 3402 22060 3408
rect 22020 1170 22048 3402
rect 22112 1601 22140 3946
rect 22848 2774 22876 10134
rect 23294 9752 23350 9761
rect 23294 9687 23350 9696
rect 23308 9654 23336 9687
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23400 7426 23428 12406
rect 23492 7954 23520 15302
rect 23584 10062 23612 17478
rect 23676 16250 23704 20538
rect 23768 20534 23796 21286
rect 23848 20868 23900 20874
rect 23848 20810 23900 20816
rect 23756 20528 23808 20534
rect 23756 20470 23808 20476
rect 23860 20398 23888 20810
rect 23848 20392 23900 20398
rect 23848 20334 23900 20340
rect 23860 19530 23888 20334
rect 23860 19514 23980 19530
rect 23860 19508 23992 19514
rect 23860 19502 23940 19508
rect 23940 19450 23992 19456
rect 23848 19440 23900 19446
rect 23848 19382 23900 19388
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23768 15502 23796 18226
rect 23860 17746 23888 19382
rect 23848 17740 23900 17746
rect 23848 17682 23900 17688
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23860 16522 23888 16934
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 23940 16516 23992 16522
rect 23940 16458 23992 16464
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 23952 15201 23980 16458
rect 24044 16182 24072 22918
rect 24596 22778 24624 23462
rect 24766 23080 24822 23089
rect 24766 23015 24822 23024
rect 24780 22982 24808 23015
rect 24768 22976 24820 22982
rect 24768 22918 24820 22924
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24872 22098 24900 24618
rect 24952 24608 25004 24614
rect 24952 24550 25004 24556
rect 24860 22092 24912 22098
rect 24860 22034 24912 22040
rect 24216 21888 24268 21894
rect 24584 21888 24636 21894
rect 24216 21830 24268 21836
rect 24582 21856 24584 21865
rect 24676 21888 24728 21894
rect 24636 21856 24638 21865
rect 24124 19916 24176 19922
rect 24124 19858 24176 19864
rect 24032 16176 24084 16182
rect 24032 16118 24084 16124
rect 23938 15192 23994 15201
rect 24136 15162 24164 19858
rect 24228 17218 24256 21830
rect 24676 21830 24728 21836
rect 24582 21791 24638 21800
rect 24584 20800 24636 20806
rect 24584 20742 24636 20748
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24400 18216 24452 18222
rect 24398 18184 24400 18193
rect 24452 18184 24454 18193
rect 24398 18119 24454 18128
rect 24504 17762 24532 18566
rect 24308 17740 24360 17746
rect 24308 17682 24360 17688
rect 24412 17734 24532 17762
rect 24320 17338 24348 17682
rect 24308 17332 24360 17338
rect 24308 17274 24360 17280
rect 24228 17190 24348 17218
rect 23938 15127 23994 15136
rect 24124 15156 24176 15162
rect 24124 15098 24176 15104
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23676 14550 23704 15030
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23676 14006 23704 14486
rect 24136 14362 24164 15098
rect 24044 14334 24164 14362
rect 24320 14346 24348 17190
rect 24308 14340 24360 14346
rect 24044 14074 24072 14334
rect 24308 14282 24360 14288
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23664 14000 23716 14006
rect 23664 13942 23716 13948
rect 23676 13462 23704 13942
rect 23664 13456 23716 13462
rect 23664 13398 23716 13404
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23768 12986 23796 13330
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 23940 11756 23992 11762
rect 23940 11698 23992 11704
rect 23848 10124 23900 10130
rect 23848 10066 23900 10072
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 23860 9926 23888 10066
rect 23848 9920 23900 9926
rect 23848 9862 23900 9868
rect 23952 8090 23980 11698
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 23480 7948 23532 7954
rect 23480 7890 23532 7896
rect 23480 7744 23532 7750
rect 23480 7686 23532 7692
rect 23308 7398 23428 7426
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23308 5778 23336 7398
rect 23388 7268 23440 7274
rect 23388 7210 23440 7216
rect 23296 5772 23348 5778
rect 23296 5714 23348 5720
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23400 4622 23428 7210
rect 23492 5710 23520 7686
rect 23664 5840 23716 5846
rect 23664 5782 23716 5788
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23388 4616 23440 4622
rect 23388 4558 23440 4564
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23492 3534 23520 5510
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23584 3058 23612 4422
rect 23676 3534 23704 5782
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 24136 3058 24164 14214
rect 24214 12744 24270 12753
rect 24214 12679 24216 12688
rect 24268 12679 24270 12688
rect 24216 12650 24268 12656
rect 24412 11150 24440 17734
rect 24596 17678 24624 20742
rect 24688 20058 24716 21830
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24676 20052 24728 20058
rect 24676 19994 24728 20000
rect 24872 18873 24900 20742
rect 24858 18864 24914 18873
rect 24858 18799 24914 18808
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24584 17672 24636 17678
rect 24490 17640 24546 17649
rect 24584 17614 24636 17620
rect 24490 17575 24492 17584
rect 24544 17575 24546 17584
rect 24492 17546 24544 17552
rect 24872 17320 24900 18566
rect 24964 18426 24992 24550
rect 25056 22574 25084 26415
rect 25226 26200 25282 27000
rect 26148 24880 26200 24886
rect 26148 24822 26200 24828
rect 25412 24064 25464 24070
rect 25412 24006 25464 24012
rect 25044 22568 25096 22574
rect 25044 22510 25096 22516
rect 25136 22432 25188 22438
rect 25136 22374 25188 22380
rect 25148 22098 25176 22374
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25136 22092 25188 22098
rect 25136 22034 25188 22040
rect 25148 21486 25176 22034
rect 25228 21616 25280 21622
rect 25228 21558 25280 21564
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25044 21004 25096 21010
rect 25044 20946 25096 20952
rect 25056 19514 25084 20946
rect 25240 20874 25268 21558
rect 25228 20868 25280 20874
rect 25228 20810 25280 20816
rect 25240 20534 25268 20810
rect 25228 20528 25280 20534
rect 25228 20470 25280 20476
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 24872 17292 24992 17320
rect 24858 17232 24914 17241
rect 24858 17167 24860 17176
rect 24912 17167 24914 17176
rect 24860 17138 24912 17144
rect 24674 16416 24730 16425
rect 24674 16351 24730 16360
rect 24688 16182 24716 16351
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 24504 13870 24532 14418
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24504 12306 24532 13806
rect 24596 12306 24624 16050
rect 24766 15872 24822 15881
rect 24766 15807 24822 15816
rect 24780 12866 24808 15807
rect 24964 14618 24992 17292
rect 25056 17202 25084 19450
rect 25240 19310 25268 20198
rect 25332 19310 25360 22170
rect 25228 19304 25280 19310
rect 25228 19246 25280 19252
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25240 18834 25268 19246
rect 25228 18828 25280 18834
rect 25228 18770 25280 18776
rect 25228 18692 25280 18698
rect 25228 18634 25280 18640
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 25044 15972 25096 15978
rect 25044 15914 25096 15920
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24872 12986 24900 14350
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24780 12850 24900 12866
rect 24768 12844 24900 12850
rect 24820 12838 24900 12844
rect 24768 12786 24820 12792
rect 24766 12608 24822 12617
rect 24766 12543 24822 12552
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24674 12200 24730 12209
rect 24674 12135 24730 12144
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24584 11008 24636 11014
rect 24584 10950 24636 10956
rect 24596 10606 24624 10950
rect 24688 10606 24716 12135
rect 24780 11694 24808 12543
rect 24872 12442 24900 12838
rect 24860 12436 24912 12442
rect 25056 12434 25084 15914
rect 25136 14612 25188 14618
rect 25136 14554 25188 14560
rect 25148 14006 25176 14554
rect 25136 14000 25188 14006
rect 25136 13942 25188 13948
rect 25240 13394 25268 18634
rect 25424 17218 25452 24006
rect 25504 23656 25556 23662
rect 25504 23598 25556 23604
rect 25516 18222 25544 23598
rect 25964 22976 26016 22982
rect 25964 22918 26016 22924
rect 25504 18216 25556 18222
rect 25504 18158 25556 18164
rect 25872 17604 25924 17610
rect 25872 17546 25924 17552
rect 25424 17190 25544 17218
rect 25412 15700 25464 15706
rect 25412 15642 25464 15648
rect 25320 13864 25372 13870
rect 25320 13806 25372 13812
rect 25228 13388 25280 13394
rect 25228 13330 25280 13336
rect 25228 13252 25280 13258
rect 25228 13194 25280 13200
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 24860 12378 24912 12384
rect 24964 12406 25084 12434
rect 24860 11824 24912 11830
rect 24858 11792 24860 11801
rect 24912 11792 24914 11801
rect 24858 11727 24914 11736
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24858 11384 24914 11393
rect 24858 11319 24914 11328
rect 24872 11218 24900 11319
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24766 10976 24822 10985
rect 24766 10911 24822 10920
rect 24584 10600 24636 10606
rect 24584 10542 24636 10548
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24674 10160 24730 10169
rect 24674 10095 24730 10104
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 24596 6798 24624 9318
rect 24688 8362 24716 10095
rect 24780 9518 24808 10911
rect 24860 10736 24912 10742
rect 24860 10678 24912 10684
rect 24872 10577 24900 10678
rect 24858 10568 24914 10577
rect 24858 10503 24914 10512
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 24964 9450 24992 12406
rect 25148 12102 25176 12582
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 25044 11280 25096 11286
rect 25044 11222 25096 11228
rect 24952 9444 25004 9450
rect 24952 9386 25004 9392
rect 24858 9344 24914 9353
rect 24858 9279 24914 9288
rect 24872 9042 24900 9279
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 24950 8528 25006 8537
rect 24950 8463 24952 8472
rect 25004 8463 25006 8472
rect 24952 8434 25004 8440
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24872 7834 24900 8298
rect 24950 8120 25006 8129
rect 24950 8055 25006 8064
rect 24964 7954 24992 8055
rect 24952 7948 25004 7954
rect 24952 7890 25004 7896
rect 25056 7886 25084 11222
rect 25134 8936 25190 8945
rect 25134 8871 25190 8880
rect 25044 7880 25096 7886
rect 24872 7806 24992 7834
rect 25044 7822 25096 7828
rect 24766 7712 24822 7721
rect 24766 7647 24822 7656
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24674 6488 24730 6497
rect 24674 6423 24730 6432
rect 24688 5166 24716 6423
rect 24780 6254 24808 7647
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 24872 7313 24900 7414
rect 24858 7304 24914 7313
rect 24858 7239 24914 7248
rect 24858 6896 24914 6905
rect 24858 6831 24860 6840
rect 24912 6831 24914 6840
rect 24860 6802 24912 6808
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24872 6089 24900 6326
rect 24858 6080 24914 6089
rect 24858 6015 24914 6024
rect 24964 5778 24992 7806
rect 25148 7478 25176 8871
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 25044 6724 25096 6730
rect 25044 6666 25096 6672
rect 24952 5772 25004 5778
rect 24952 5714 25004 5720
rect 24950 5672 25006 5681
rect 24950 5607 24952 5616
rect 25004 5607 25006 5616
rect 24952 5578 25004 5584
rect 24766 5264 24822 5273
rect 24766 5199 24822 5208
rect 24676 5160 24728 5166
rect 24676 5102 24728 5108
rect 24780 4078 24808 5199
rect 24952 5092 25004 5098
rect 24952 5034 25004 5040
rect 24964 4865 24992 5034
rect 24950 4856 25006 4865
rect 24950 4791 25006 4800
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 24964 4457 24992 4490
rect 24950 4448 25006 4457
rect 24950 4383 25006 4392
rect 25056 4146 25084 6666
rect 25240 6662 25268 13194
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25044 4140 25096 4146
rect 25044 4082 25096 4088
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 25226 4040 25282 4049
rect 24952 4004 25004 4010
rect 25226 3975 25282 3984
rect 24952 3946 25004 3952
rect 24964 3641 24992 3946
rect 24950 3632 25006 3641
rect 24950 3567 25006 3576
rect 25136 3460 25188 3466
rect 25136 3402 25188 3408
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 24124 3052 24176 3058
rect 24124 2994 24176 3000
rect 22756 2746 22876 2774
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 22192 2644 22244 2650
rect 22192 2586 22244 2592
rect 22204 2009 22232 2586
rect 22756 2446 22784 2746
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 24596 2446 24624 3334
rect 25148 3233 25176 3402
rect 25134 3224 25190 3233
rect 25134 3159 25190 3168
rect 25240 3126 25268 3975
rect 25332 3194 25360 13806
rect 25424 10062 25452 15642
rect 25516 11898 25544 17190
rect 25688 17060 25740 17066
rect 25688 17002 25740 17008
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 25504 11892 25556 11898
rect 25504 11834 25556 11840
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 25608 6322 25636 16594
rect 25700 7342 25728 17002
rect 25780 15564 25832 15570
rect 25780 15506 25832 15512
rect 25688 7336 25740 7342
rect 25688 7278 25740 7284
rect 25596 6316 25648 6322
rect 25596 6258 25648 6264
rect 25792 4146 25820 15506
rect 25884 7818 25912 17546
rect 25976 11257 26004 22918
rect 26056 19780 26108 19786
rect 26056 19722 26108 19728
rect 26068 11558 26096 19722
rect 26160 14618 26188 24822
rect 26148 14612 26200 14618
rect 26148 14554 26200 14560
rect 26056 11552 26108 11558
rect 26056 11494 26108 11500
rect 25962 11248 26018 11257
rect 25962 11183 26018 11192
rect 25872 7812 25924 7818
rect 25872 7754 25924 7760
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 24860 3120 24912 3126
rect 24860 3062 24912 3068
rect 25228 3120 25280 3126
rect 25228 3062 25280 3068
rect 24872 2825 24900 3062
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 24858 2816 24914 2825
rect 24858 2751 24914 2760
rect 22744 2440 22796 2446
rect 22744 2382 22796 2388
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24950 2408 25006 2417
rect 23388 2372 23440 2378
rect 24950 2343 24952 2352
rect 23388 2314 23440 2320
rect 25004 2343 25006 2352
rect 24952 2314 25004 2320
rect 22190 2000 22246 2009
rect 22190 1935 22246 1944
rect 22098 1592 22154 1601
rect 22098 1527 22154 1536
rect 22098 1184 22154 1193
rect 22020 1142 22098 1170
rect 22098 1119 22154 1128
rect 6734 0 6790 800
rect 20166 0 20222 800
rect 23400 377 23428 2314
rect 25056 785 25084 2926
rect 25042 776 25098 785
rect 25042 711 25098 720
rect 23386 368 23442 377
rect 23386 303 23442 312
<< via2 >>
rect 1306 23724 1362 23760
rect 1306 23704 1308 23724
rect 1308 23704 1360 23724
rect 1360 23704 1362 23724
rect 1306 22636 1362 22672
rect 1306 22616 1308 22636
rect 1308 22616 1360 22636
rect 1360 22616 1362 22636
rect 2134 26152 2190 26208
rect 1582 18808 1638 18864
rect 2778 24792 2834 24848
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 3422 25880 3478 25936
rect 3698 22072 3754 22128
rect 3606 21392 3662 21448
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2226 19896 2282 19952
rect 2318 19352 2374 19408
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 4158 24248 4214 24304
rect 4066 20848 4122 20904
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 4526 19760 4582 19816
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 4710 19216 4766 19272
rect 5262 24928 5318 24984
rect 4710 17720 4766 17776
rect 4618 14456 4674 14512
rect 4526 12824 4582 12880
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 5170 18672 5226 18728
rect 5538 20304 5594 20360
rect 5630 18164 5632 18184
rect 5632 18164 5684 18184
rect 5684 18164 5686 18184
rect 5630 18128 5686 18164
rect 6550 25064 6606 25120
rect 6366 24656 6422 24712
rect 6182 23568 6238 23624
rect 6274 22208 6330 22264
rect 5538 17196 5594 17232
rect 5538 17176 5540 17196
rect 5540 17176 5592 17196
rect 5592 17176 5594 17196
rect 5262 16652 5318 16688
rect 5262 16632 5264 16652
rect 5264 16632 5316 16652
rect 5316 16632 5318 16652
rect 6458 17856 6514 17912
rect 6918 23604 6920 23624
rect 6920 23604 6972 23624
rect 6972 23604 6974 23624
rect 6918 23568 6974 23604
rect 7102 23588 7158 23624
rect 7102 23568 7104 23588
rect 7104 23568 7156 23588
rect 7156 23568 7158 23588
rect 7102 22616 7158 22672
rect 7378 21972 7380 21992
rect 7380 21972 7432 21992
rect 7432 21972 7434 21992
rect 7378 21936 7434 21972
rect 7286 21528 7342 21584
rect 7194 17584 7250 17640
rect 7102 17040 7158 17096
rect 7562 23160 7618 23216
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7562 18944 7618 19000
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 8390 23024 8446 23080
rect 8666 22752 8722 22808
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 8482 21664 8538 21720
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7746 19080 7802 19136
rect 7470 17992 7526 18048
rect 7746 17992 7802 18048
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7838 17720 7894 17776
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 8574 19372 8630 19408
rect 8574 19352 8576 19372
rect 8576 19352 8628 19372
rect 8628 19352 8630 19372
rect 8850 23976 8906 24032
rect 9954 24792 10010 24848
rect 9310 21836 9312 21856
rect 9312 21836 9364 21856
rect 9364 21836 9366 21856
rect 9310 21800 9366 21836
rect 9310 20576 9366 20632
rect 9310 20032 9366 20088
rect 9586 24112 9642 24168
rect 9218 18264 9274 18320
rect 9402 17856 9458 17912
rect 8850 17584 8906 17640
rect 9402 17176 9458 17232
rect 9310 16768 9366 16824
rect 9678 21800 9734 21856
rect 9678 18944 9734 19000
rect 10046 16940 10048 16960
rect 10048 16940 10100 16960
rect 10100 16940 10102 16960
rect 10046 16904 10102 16940
rect 8758 16360 8814 16416
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 8666 16108 8722 16144
rect 8666 16088 8668 16108
rect 8668 16088 8720 16108
rect 8720 16088 8722 16108
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7654 15000 7710 15056
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 6550 13912 6606 13968
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 5538 12144 5594 12200
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 9126 15972 9182 16008
rect 9126 15952 9128 15972
rect 9128 15952 9180 15972
rect 9180 15952 9182 15972
rect 9770 16224 9826 16280
rect 9678 15816 9734 15872
rect 10598 23840 10654 23896
rect 10322 19488 10378 19544
rect 10414 18400 10470 18456
rect 11518 23704 11574 23760
rect 10966 22344 11022 22400
rect 11150 20440 11206 20496
rect 10782 19352 10838 19408
rect 10414 16768 10470 16824
rect 10322 16496 10378 16552
rect 10230 16224 10286 16280
rect 10046 15544 10102 15600
rect 11334 18536 11390 18592
rect 11610 20032 11666 20088
rect 12070 22888 12126 22944
rect 11794 22480 11850 22536
rect 11610 16904 11666 16960
rect 12254 21256 12310 21312
rect 11886 20984 11942 21040
rect 12438 22208 12494 22264
rect 12622 22344 12678 22400
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 13818 23976 13874 24032
rect 14002 23296 14058 23352
rect 13174 21392 13230 21448
rect 12714 21256 12770 21312
rect 12438 20596 12494 20632
rect 12438 20576 12440 20596
rect 12440 20576 12492 20596
rect 12492 20576 12494 20596
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 11886 19080 11942 19136
rect 11978 17856 12034 17912
rect 11886 16904 11942 16960
rect 13266 20868 13322 20904
rect 13266 20848 13268 20868
rect 13268 20848 13320 20868
rect 13320 20848 13322 20868
rect 12622 17720 12678 17776
rect 12622 16904 12678 16960
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12806 19352 12862 19408
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 13910 21800 13966 21856
rect 13818 21120 13874 21176
rect 13726 20848 13782 20904
rect 13542 20712 13598 20768
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13266 16668 13268 16688
rect 13268 16668 13320 16688
rect 13320 16668 13322 16688
rect 13266 16632 13322 16668
rect 12806 16360 12862 16416
rect 12254 15816 12310 15872
rect 11886 14320 11942 14376
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 13450 16632 13506 16688
rect 13450 14764 13452 14784
rect 13452 14764 13504 14784
rect 13504 14764 13506 14784
rect 13450 14728 13506 14764
rect 13450 14592 13506 14648
rect 13358 14048 13414 14104
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12806 12688 12862 12744
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 13910 18944 13966 19000
rect 13726 18808 13782 18864
rect 14370 22480 14426 22536
rect 14370 22344 14426 22400
rect 14278 20032 14334 20088
rect 14554 21256 14610 21312
rect 14278 17992 14334 18048
rect 13910 15408 13966 15464
rect 14738 21528 14794 21584
rect 14738 20168 14794 20224
rect 15014 21528 15070 21584
rect 14738 19352 14794 19408
rect 15290 19352 15346 19408
rect 15106 17720 15162 17776
rect 14646 15680 14702 15736
rect 14830 14864 14886 14920
rect 15198 16632 15254 16688
rect 15934 23568 15990 23624
rect 15658 22752 15714 22808
rect 15566 21392 15622 21448
rect 15474 17720 15530 17776
rect 16026 21664 16082 21720
rect 15842 20576 15898 20632
rect 15934 20440 15990 20496
rect 15934 20304 15990 20360
rect 15842 19352 15898 19408
rect 15658 17448 15714 17504
rect 15842 17856 15898 17912
rect 15658 13640 15714 13696
rect 15106 13504 15162 13560
rect 16578 23976 16634 24032
rect 16670 20440 16726 20496
rect 16394 20304 16450 20360
rect 16486 20032 16542 20088
rect 16302 19660 16304 19680
rect 16304 19660 16356 19680
rect 16356 19660 16358 19680
rect 16302 19624 16358 19660
rect 16578 19488 16634 19544
rect 16210 18808 16266 18864
rect 16210 17448 16266 17504
rect 16578 18536 16634 18592
rect 16486 18420 16542 18456
rect 16486 18400 16488 18420
rect 16488 18400 16540 18420
rect 16540 18400 16542 18420
rect 16302 16904 16358 16960
rect 16118 11228 16120 11248
rect 16120 11228 16172 11248
rect 16172 11228 16174 11248
rect 16118 11192 16174 11228
rect 17038 23840 17094 23896
rect 17038 23568 17094 23624
rect 16946 22888 17002 22944
rect 16854 22480 16910 22536
rect 16946 20712 17002 20768
rect 17130 18944 17186 19000
rect 17406 23432 17462 23488
rect 17406 21256 17462 21312
rect 17222 17876 17278 17912
rect 17222 17856 17224 17876
rect 17224 17856 17276 17876
rect 17276 17856 17278 17876
rect 17222 17060 17278 17096
rect 17222 17040 17224 17060
rect 17224 17040 17276 17060
rect 17276 17040 17278 17060
rect 17958 24268 18014 24304
rect 17958 24248 17960 24268
rect 17960 24248 18012 24268
rect 18012 24248 18014 24268
rect 17774 23976 17830 24032
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17682 21120 17738 21176
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 18970 24656 19026 24712
rect 18602 23160 18658 23216
rect 18602 23044 18658 23080
rect 18602 23024 18604 23044
rect 18604 23024 18656 23044
rect 18656 23024 18658 23044
rect 18510 22480 18566 22536
rect 18694 22344 18750 22400
rect 18786 22208 18842 22264
rect 18326 21528 18382 21584
rect 18418 21392 18474 21448
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17498 16632 17554 16688
rect 17682 14048 17738 14104
rect 18050 18844 18052 18864
rect 18052 18844 18104 18864
rect 18104 18844 18106 18864
rect 18050 18808 18106 18844
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18142 17040 18198 17096
rect 18326 17060 18382 17096
rect 18326 17040 18328 17060
rect 18328 17040 18380 17060
rect 18380 17040 18382 17060
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18418 15272 18474 15328
rect 18418 14320 18474 14376
rect 18326 12552 18382 12608
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18970 21936 19026 21992
rect 19798 26152 19854 26208
rect 19614 22616 19670 22672
rect 19430 21800 19486 21856
rect 19522 21664 19578 21720
rect 19246 20440 19302 20496
rect 18970 17040 19026 17096
rect 19154 15680 19210 15736
rect 19430 16768 19486 16824
rect 19062 14592 19118 14648
rect 18970 14320 19026 14376
rect 18878 14220 18880 14240
rect 18880 14220 18932 14240
rect 18932 14220 18934 14240
rect 18878 14184 18934 14220
rect 18694 12164 18750 12200
rect 18694 12144 18696 12164
rect 18696 12144 18748 12164
rect 18748 12144 18750 12164
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 15106 8336 15162 8392
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 19706 18944 19762 19000
rect 19706 17992 19762 18048
rect 19798 17856 19854 17912
rect 19798 17740 19854 17776
rect 19798 17720 19800 17740
rect 19800 17720 19852 17740
rect 19852 17720 19854 17740
rect 19614 14184 19670 14240
rect 19062 13232 19118 13288
rect 20166 15680 20222 15736
rect 20074 14456 20130 14512
rect 19430 10260 19486 10296
rect 19430 10240 19432 10260
rect 19432 10240 19484 10260
rect 19484 10240 19486 10260
rect 19246 9968 19302 10024
rect 19430 9444 19486 9480
rect 19430 9424 19432 9444
rect 19432 9424 19484 9444
rect 19484 9424 19486 9444
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 19706 11076 19762 11112
rect 19706 11056 19708 11076
rect 19708 11056 19760 11076
rect 19760 11056 19762 11076
rect 20626 23296 20682 23352
rect 22190 26288 22246 26344
rect 22006 25608 22062 25664
rect 21914 24112 21970 24168
rect 20902 23024 20958 23080
rect 23478 26016 23534 26072
rect 22374 23432 22430 23488
rect 21362 22208 21418 22264
rect 21730 22072 21786 22128
rect 21546 21936 21602 21992
rect 20718 20304 20774 20360
rect 21454 21800 21510 21856
rect 20994 19760 21050 19816
rect 21178 19488 21234 19544
rect 20902 18300 20904 18320
rect 20904 18300 20956 18320
rect 20956 18300 20958 18320
rect 20902 18264 20958 18300
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 20718 10376 20774 10432
rect 21546 20440 21602 20496
rect 22190 22516 22192 22536
rect 22192 22516 22244 22536
rect 22244 22516 22246 22536
rect 22190 22480 22246 22516
rect 21822 19508 21878 19544
rect 21822 19488 21824 19508
rect 21824 19488 21876 19508
rect 21876 19488 21878 19508
rect 22006 19488 22062 19544
rect 22190 20712 22246 20768
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 23386 23704 23442 23760
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22650 23024 22706 23080
rect 22374 21528 22430 21584
rect 22466 21392 22522 21448
rect 22834 23160 22890 23216
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22650 20868 22706 20904
rect 22650 20848 22652 20868
rect 22652 20848 22704 20868
rect 22704 20848 22706 20868
rect 22558 19896 22614 19952
rect 22466 19624 22522 19680
rect 22190 19508 22246 19544
rect 22190 19488 22192 19508
rect 22192 19488 22244 19508
rect 22244 19488 22246 19508
rect 22098 19080 22154 19136
rect 22282 18536 22338 18592
rect 21914 16632 21970 16688
rect 21546 14456 21602 14512
rect 22098 17448 22154 17504
rect 22742 19896 22798 19952
rect 23846 24384 23902 24440
rect 25042 26424 25098 26480
rect 24766 25200 24822 25256
rect 24398 24928 24454 24984
rect 23846 23568 23902 23624
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 23018 19488 23074 19544
rect 23110 19352 23166 19408
rect 22834 19216 22890 19272
rect 22742 18944 22798 19000
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22466 17312 22522 17368
rect 22466 17040 22522 17096
rect 22098 16904 22154 16960
rect 22098 13932 22154 13968
rect 22098 13912 22100 13932
rect 22100 13912 22152 13932
rect 22152 13912 22154 13932
rect 20994 11328 21050 11384
rect 22282 13096 22338 13152
rect 22190 12824 22246 12880
rect 22282 12280 22338 12336
rect 22466 15408 22522 15464
rect 22466 12824 22522 12880
rect 23018 18692 23074 18728
rect 23018 18672 23020 18692
rect 23020 18672 23072 18692
rect 23072 18672 23074 18692
rect 23386 19116 23388 19136
rect 23388 19116 23440 19136
rect 23440 19116 23442 19136
rect 23386 19080 23442 19116
rect 23110 18300 23112 18320
rect 23112 18300 23164 18320
rect 23164 18300 23166 18320
rect 23110 18264 23166 18300
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23018 17720 23074 17776
rect 23018 17040 23074 17096
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 22834 15308 22836 15328
rect 22836 15308 22888 15328
rect 22888 15308 22890 15328
rect 22834 15272 22890 15308
rect 22742 15000 22798 15056
rect 22742 13776 22798 13832
rect 22742 13096 22798 13152
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 23478 16224 23534 16280
rect 23294 14184 23350 14240
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22006 6976 22062 7032
rect 22650 5480 22706 5536
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 23386 13368 23442 13424
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23294 9696 23350 9752
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 24766 23024 24822 23080
rect 24582 21836 24584 21856
rect 24584 21836 24636 21856
rect 24636 21836 24638 21856
rect 23938 15136 23994 15192
rect 24582 21800 24638 21836
rect 24398 18164 24400 18184
rect 24400 18164 24452 18184
rect 24452 18164 24454 18184
rect 24398 18128 24454 18164
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 24214 12708 24270 12744
rect 24214 12688 24216 12708
rect 24216 12688 24268 12708
rect 24268 12688 24270 12708
rect 24858 18808 24914 18864
rect 24490 17604 24546 17640
rect 24490 17584 24492 17604
rect 24492 17584 24544 17604
rect 24544 17584 24546 17604
rect 24858 17196 24914 17232
rect 24858 17176 24860 17196
rect 24860 17176 24912 17196
rect 24912 17176 24914 17196
rect 24674 16360 24730 16416
rect 24766 15816 24822 15872
rect 24766 12552 24822 12608
rect 24674 12144 24730 12200
rect 24858 11772 24860 11792
rect 24860 11772 24912 11792
rect 24912 11772 24914 11792
rect 24858 11736 24914 11772
rect 24858 11328 24914 11384
rect 24766 10920 24822 10976
rect 24674 10104 24730 10160
rect 24858 10512 24914 10568
rect 24858 9288 24914 9344
rect 24950 8492 25006 8528
rect 24950 8472 24952 8492
rect 24952 8472 25004 8492
rect 25004 8472 25006 8492
rect 24950 8064 25006 8120
rect 25134 8880 25190 8936
rect 24766 7656 24822 7712
rect 24674 6432 24730 6488
rect 24858 7248 24914 7304
rect 24858 6860 24914 6896
rect 24858 6840 24860 6860
rect 24860 6840 24912 6860
rect 24912 6840 24914 6860
rect 24858 6024 24914 6080
rect 24950 5636 25006 5672
rect 24950 5616 24952 5636
rect 24952 5616 25004 5636
rect 25004 5616 25006 5636
rect 24766 5208 24822 5264
rect 24950 4800 25006 4856
rect 24950 4392 25006 4448
rect 25226 3984 25282 4040
rect 24950 3576 25006 3632
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 25134 3168 25190 3224
rect 25962 11192 26018 11248
rect 24858 2760 24914 2816
rect 24950 2372 25006 2408
rect 24950 2352 24952 2372
rect 24952 2352 25004 2372
rect 25004 2352 25006 2372
rect 22190 1944 22246 2000
rect 22098 1536 22154 1592
rect 22098 1128 22154 1184
rect 25042 720 25098 776
rect 23386 312 23442 368
<< metal3 >>
rect 25037 26482 25103 26485
rect 26200 26482 27000 26512
rect 25037 26480 27000 26482
rect 25037 26424 25042 26480
rect 25098 26424 27000 26480
rect 25037 26422 27000 26424
rect 25037 26419 25103 26422
rect 26200 26392 27000 26422
rect 22185 26346 22251 26349
rect 2270 26344 22251 26346
rect 2270 26288 22190 26344
rect 22246 26288 22251 26344
rect 2270 26286 22251 26288
rect 2129 26210 2195 26213
rect 2270 26210 2330 26286
rect 22185 26283 22251 26286
rect 2129 26208 2330 26210
rect 2129 26152 2134 26208
rect 2190 26152 2330 26208
rect 2129 26150 2330 26152
rect 2129 26147 2195 26150
rect 4838 26148 4844 26212
rect 4908 26210 4914 26212
rect 19793 26210 19859 26213
rect 4908 26208 19859 26210
rect 4908 26152 19798 26208
rect 19854 26152 19859 26208
rect 4908 26150 19859 26152
rect 4908 26148 4914 26150
rect 19793 26147 19859 26150
rect 23473 26074 23539 26077
rect 26200 26074 27000 26104
rect 23473 26072 27000 26074
rect 23473 26016 23478 26072
rect 23534 26016 27000 26072
rect 23473 26014 27000 26016
rect 23473 26011 23539 26014
rect 26200 25984 27000 26014
rect 0 25938 800 25968
rect 3417 25938 3483 25941
rect 0 25936 3483 25938
rect 0 25880 3422 25936
rect 3478 25880 3483 25936
rect 0 25878 3483 25880
rect 0 25848 800 25878
rect 3417 25875 3483 25878
rect 22001 25666 22067 25669
rect 26200 25666 27000 25696
rect 22001 25664 27000 25666
rect 22001 25608 22006 25664
rect 22062 25608 27000 25664
rect 22001 25606 27000 25608
rect 22001 25603 22067 25606
rect 26200 25576 27000 25606
rect 24761 25258 24827 25261
rect 26200 25258 27000 25288
rect 24761 25256 27000 25258
rect 24761 25200 24766 25256
rect 24822 25200 27000 25256
rect 24761 25198 27000 25200
rect 24761 25195 24827 25198
rect 26200 25168 27000 25198
rect 6545 25122 6611 25125
rect 19374 25122 19380 25124
rect 6545 25120 19380 25122
rect 6545 25064 6550 25120
rect 6606 25064 19380 25120
rect 6545 25062 19380 25064
rect 6545 25059 6611 25062
rect 19374 25060 19380 25062
rect 19444 25060 19450 25124
rect 5257 24986 5323 24989
rect 24393 24986 24459 24989
rect 5257 24984 24459 24986
rect 5257 24928 5262 24984
rect 5318 24928 24398 24984
rect 24454 24928 24459 24984
rect 5257 24926 24459 24928
rect 5257 24923 5323 24926
rect 24393 24923 24459 24926
rect 0 24850 800 24880
rect 2773 24850 2839 24853
rect 0 24848 2839 24850
rect 0 24792 2778 24848
rect 2834 24792 2839 24848
rect 0 24790 2839 24792
rect 0 24760 800 24790
rect 2773 24787 2839 24790
rect 9949 24850 10015 24853
rect 26200 24850 27000 24880
rect 9949 24848 27000 24850
rect 9949 24792 9954 24848
rect 10010 24792 27000 24848
rect 9949 24790 27000 24792
rect 9949 24787 10015 24790
rect 26200 24760 27000 24790
rect 6361 24714 6427 24717
rect 18965 24714 19031 24717
rect 6361 24712 19031 24714
rect 6361 24656 6366 24712
rect 6422 24656 18970 24712
rect 19026 24656 19031 24712
rect 6361 24654 19031 24656
rect 6361 24651 6427 24654
rect 18965 24651 19031 24654
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 23841 24442 23907 24445
rect 26200 24442 27000 24472
rect 23841 24440 27000 24442
rect 23841 24384 23846 24440
rect 23902 24384 27000 24440
rect 23841 24382 27000 24384
rect 23841 24379 23907 24382
rect 26200 24352 27000 24382
rect 4153 24306 4219 24309
rect 17953 24306 18019 24309
rect 4153 24304 18019 24306
rect 4153 24248 4158 24304
rect 4214 24248 17958 24304
rect 18014 24248 18019 24304
rect 4153 24246 18019 24248
rect 4153 24243 4219 24246
rect 17953 24243 18019 24246
rect 9581 24170 9647 24173
rect 21909 24170 21975 24173
rect 9581 24168 21975 24170
rect 9581 24112 9586 24168
rect 9642 24112 21914 24168
rect 21970 24112 21975 24168
rect 9581 24110 21975 24112
rect 9581 24107 9647 24110
rect 21909 24107 21975 24110
rect 8845 24034 8911 24037
rect 13813 24034 13879 24037
rect 8845 24032 13879 24034
rect 8845 23976 8850 24032
rect 8906 23976 13818 24032
rect 13874 23976 13879 24032
rect 8845 23974 13879 23976
rect 8845 23971 8911 23974
rect 13813 23971 13879 23974
rect 16573 24034 16639 24037
rect 17769 24034 17835 24037
rect 26200 24034 27000 24064
rect 16573 24032 17835 24034
rect 16573 23976 16578 24032
rect 16634 23976 17774 24032
rect 17830 23976 17835 24032
rect 16573 23974 17835 23976
rect 16573 23971 16639 23974
rect 17769 23971 17835 23974
rect 22050 23974 27000 24034
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 10593 23898 10659 23901
rect 17033 23898 17099 23901
rect 22050 23898 22110 23974
rect 26200 23944 27000 23974
rect 10593 23896 17099 23898
rect 10593 23840 10598 23896
rect 10654 23840 17038 23896
rect 17094 23840 17099 23896
rect 10593 23838 17099 23840
rect 10593 23835 10659 23838
rect 17033 23835 17099 23838
rect 18462 23838 22110 23898
rect 0 23762 800 23792
rect 1301 23762 1367 23765
rect 0 23760 1367 23762
rect 0 23704 1306 23760
rect 1362 23704 1367 23760
rect 0 23702 1367 23704
rect 0 23672 800 23702
rect 1301 23699 1367 23702
rect 11513 23762 11579 23765
rect 18462 23762 18522 23838
rect 11513 23760 18522 23762
rect 11513 23704 11518 23760
rect 11574 23704 18522 23760
rect 11513 23702 18522 23704
rect 23381 23762 23447 23765
rect 23381 23760 24042 23762
rect 23381 23704 23386 23760
rect 23442 23704 24042 23760
rect 23381 23702 24042 23704
rect 11513 23699 11579 23702
rect 23381 23699 23447 23702
rect 6177 23626 6243 23629
rect 6913 23626 6979 23629
rect 6177 23624 6979 23626
rect 6177 23568 6182 23624
rect 6238 23568 6918 23624
rect 6974 23568 6979 23624
rect 6177 23566 6979 23568
rect 6177 23563 6243 23566
rect 6913 23563 6979 23566
rect 7097 23626 7163 23629
rect 15929 23626 15995 23629
rect 7097 23624 15995 23626
rect 7097 23568 7102 23624
rect 7158 23568 15934 23624
rect 15990 23568 15995 23624
rect 7097 23566 15995 23568
rect 7097 23563 7163 23566
rect 15929 23563 15995 23566
rect 17033 23626 17099 23629
rect 23841 23626 23907 23629
rect 17033 23624 23907 23626
rect 17033 23568 17038 23624
rect 17094 23568 23846 23624
rect 23902 23568 23907 23624
rect 17033 23566 23907 23568
rect 23982 23626 24042 23702
rect 26200 23626 27000 23656
rect 23982 23566 27000 23626
rect 17033 23563 17099 23566
rect 23841 23563 23907 23566
rect 26200 23536 27000 23566
rect 17401 23490 17467 23493
rect 17534 23490 17540 23492
rect 17401 23488 17540 23490
rect 17401 23432 17406 23488
rect 17462 23432 17540 23488
rect 17401 23430 17540 23432
rect 17401 23427 17467 23430
rect 17534 23428 17540 23430
rect 17604 23428 17610 23492
rect 22134 23428 22140 23492
rect 22204 23490 22210 23492
rect 22369 23490 22435 23493
rect 22204 23488 22435 23490
rect 22204 23432 22374 23488
rect 22430 23432 22435 23488
rect 22204 23430 22435 23432
rect 22204 23428 22210 23430
rect 22369 23427 22435 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 13997 23354 14063 23357
rect 20621 23354 20687 23357
rect 13997 23352 20687 23354
rect 13997 23296 14002 23352
rect 14058 23296 20626 23352
rect 20682 23296 20687 23352
rect 13997 23294 20687 23296
rect 13997 23291 14063 23294
rect 20621 23291 20687 23294
rect 7557 23218 7623 23221
rect 18597 23218 18663 23221
rect 7557 23216 18663 23218
rect 7557 23160 7562 23216
rect 7618 23160 18602 23216
rect 18658 23160 18663 23216
rect 7557 23158 18663 23160
rect 7557 23155 7623 23158
rect 18597 23155 18663 23158
rect 22829 23218 22895 23221
rect 26200 23218 27000 23248
rect 22829 23216 27000 23218
rect 22829 23160 22834 23216
rect 22890 23160 27000 23216
rect 22829 23158 27000 23160
rect 22829 23155 22895 23158
rect 26200 23128 27000 23158
rect 8385 23082 8451 23085
rect 18597 23082 18663 23085
rect 8385 23080 18663 23082
rect 8385 23024 8390 23080
rect 8446 23024 18602 23080
rect 18658 23024 18663 23080
rect 8385 23022 18663 23024
rect 8385 23019 8451 23022
rect 18597 23019 18663 23022
rect 20897 23082 20963 23085
rect 22645 23082 22711 23085
rect 24761 23082 24827 23085
rect 20897 23080 24827 23082
rect 20897 23024 20902 23080
rect 20958 23024 22650 23080
rect 22706 23024 24766 23080
rect 24822 23024 24827 23080
rect 20897 23022 24827 23024
rect 20897 23019 20963 23022
rect 22645 23019 22711 23022
rect 24761 23019 24827 23022
rect 12065 22946 12131 22949
rect 16941 22946 17007 22949
rect 12065 22944 17007 22946
rect 12065 22888 12070 22944
rect 12126 22888 16946 22944
rect 17002 22888 17007 22944
rect 12065 22886 17007 22888
rect 12065 22883 12131 22886
rect 16941 22883 17007 22886
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 8661 22810 8727 22813
rect 15653 22810 15719 22813
rect 8661 22808 15719 22810
rect 8661 22752 8666 22808
rect 8722 22752 15658 22808
rect 15714 22752 15719 22808
rect 8661 22750 15719 22752
rect 8661 22747 8727 22750
rect 15653 22747 15719 22750
rect 20110 22748 20116 22812
rect 20180 22810 20186 22812
rect 26200 22810 27000 22840
rect 20180 22750 27000 22810
rect 20180 22748 20186 22750
rect 26200 22720 27000 22750
rect 0 22674 800 22704
rect 1301 22674 1367 22677
rect 0 22672 1367 22674
rect 0 22616 1306 22672
rect 1362 22616 1367 22672
rect 0 22614 1367 22616
rect 0 22584 800 22614
rect 1301 22611 1367 22614
rect 7097 22674 7163 22677
rect 19609 22674 19675 22677
rect 7097 22672 19675 22674
rect 7097 22616 7102 22672
rect 7158 22616 19614 22672
rect 19670 22616 19675 22672
rect 7097 22614 19675 22616
rect 7097 22611 7163 22614
rect 19609 22611 19675 22614
rect 11789 22538 11855 22541
rect 14365 22538 14431 22541
rect 16849 22540 16915 22541
rect 16798 22538 16804 22540
rect 11789 22536 14431 22538
rect 11789 22480 11794 22536
rect 11850 22480 14370 22536
rect 14426 22480 14431 22536
rect 11789 22478 14431 22480
rect 16758 22478 16804 22538
rect 16868 22536 16915 22540
rect 16910 22480 16915 22536
rect 11789 22475 11855 22478
rect 14365 22475 14431 22478
rect 16798 22476 16804 22478
rect 16868 22476 16915 22480
rect 16849 22475 16915 22476
rect 18505 22538 18571 22541
rect 18638 22538 18644 22540
rect 18505 22536 18644 22538
rect 18505 22480 18510 22536
rect 18566 22480 18644 22536
rect 18505 22478 18644 22480
rect 18505 22475 18571 22478
rect 18638 22476 18644 22478
rect 18708 22476 18714 22540
rect 22185 22538 22251 22541
rect 22185 22536 23490 22538
rect 22185 22480 22190 22536
rect 22246 22480 23490 22536
rect 22185 22478 23490 22480
rect 22185 22475 22251 22478
rect 10961 22402 11027 22405
rect 12617 22402 12683 22405
rect 10961 22400 12683 22402
rect 10961 22344 10966 22400
rect 11022 22344 12622 22400
rect 12678 22344 12683 22400
rect 10961 22342 12683 22344
rect 10961 22339 11027 22342
rect 12617 22339 12683 22342
rect 14365 22402 14431 22405
rect 18689 22402 18755 22405
rect 14365 22400 18755 22402
rect 14365 22344 14370 22400
rect 14426 22344 18694 22400
rect 18750 22344 18755 22400
rect 14365 22342 18755 22344
rect 23430 22402 23490 22478
rect 26200 22402 27000 22432
rect 23430 22342 27000 22402
rect 14365 22339 14431 22342
rect 18689 22339 18755 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 26200 22312 27000 22342
rect 22946 22271 23262 22272
rect 6269 22266 6335 22269
rect 12433 22266 12499 22269
rect 6269 22264 12499 22266
rect 6269 22208 6274 22264
rect 6330 22208 12438 22264
rect 12494 22208 12499 22264
rect 6269 22206 12499 22208
rect 6269 22203 6335 22206
rect 12433 22203 12499 22206
rect 18781 22266 18847 22269
rect 21357 22266 21423 22269
rect 18781 22264 21423 22266
rect 18781 22208 18786 22264
rect 18842 22208 21362 22264
rect 21418 22208 21423 22264
rect 18781 22206 21423 22208
rect 18781 22203 18847 22206
rect 21357 22203 21423 22206
rect 3693 22130 3759 22133
rect 21725 22130 21791 22133
rect 3693 22128 21791 22130
rect 3693 22072 3698 22128
rect 3754 22072 21730 22128
rect 21786 22072 21791 22128
rect 3693 22070 21791 22072
rect 3693 22067 3759 22070
rect 21725 22067 21791 22070
rect 7373 21994 7439 21997
rect 18965 21994 19031 21997
rect 7373 21992 19031 21994
rect 7373 21936 7378 21992
rect 7434 21936 18970 21992
rect 19026 21936 19031 21992
rect 7373 21934 19031 21936
rect 7373 21931 7439 21934
rect 18965 21931 19031 21934
rect 21541 21994 21607 21997
rect 26200 21994 27000 22024
rect 21541 21992 27000 21994
rect 21541 21936 21546 21992
rect 21602 21936 27000 21992
rect 21541 21934 27000 21936
rect 21541 21931 21607 21934
rect 26200 21904 27000 21934
rect 9305 21858 9371 21861
rect 9438 21858 9444 21860
rect 9305 21856 9444 21858
rect 9305 21800 9310 21856
rect 9366 21800 9444 21856
rect 9305 21798 9444 21800
rect 9305 21795 9371 21798
rect 9438 21796 9444 21798
rect 9508 21796 9514 21860
rect 9673 21858 9739 21861
rect 13905 21858 13971 21861
rect 9673 21856 13971 21858
rect 9673 21800 9678 21856
rect 9734 21800 13910 21856
rect 13966 21800 13971 21856
rect 9673 21798 13971 21800
rect 9673 21795 9739 21798
rect 13905 21795 13971 21798
rect 19425 21858 19491 21861
rect 21449 21858 21515 21861
rect 24577 21860 24643 21861
rect 19425 21856 21515 21858
rect 19425 21800 19430 21856
rect 19486 21800 21454 21856
rect 21510 21800 21515 21856
rect 19425 21798 21515 21800
rect 19425 21795 19491 21798
rect 21449 21795 21515 21798
rect 24526 21796 24532 21860
rect 24596 21858 24643 21860
rect 24596 21856 24688 21858
rect 24638 21800 24688 21856
rect 24596 21798 24688 21800
rect 24596 21796 24643 21798
rect 24577 21795 24643 21796
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 8477 21722 8543 21725
rect 16021 21722 16087 21725
rect 8477 21720 16087 21722
rect 8477 21664 8482 21720
rect 8538 21664 16026 21720
rect 16082 21664 16087 21720
rect 8477 21662 16087 21664
rect 8477 21659 8543 21662
rect 16021 21659 16087 21662
rect 19517 21722 19583 21725
rect 19742 21722 19748 21724
rect 19517 21720 19748 21722
rect 19517 21664 19522 21720
rect 19578 21664 19748 21720
rect 19517 21662 19748 21664
rect 19517 21659 19583 21662
rect 19742 21660 19748 21662
rect 19812 21660 19818 21724
rect 7281 21586 7347 21589
rect 14733 21586 14799 21589
rect 7281 21584 14799 21586
rect 7281 21528 7286 21584
rect 7342 21528 14738 21584
rect 14794 21528 14799 21584
rect 7281 21526 14799 21528
rect 7281 21523 7347 21526
rect 14733 21523 14799 21526
rect 15009 21586 15075 21589
rect 18321 21586 18387 21589
rect 15009 21584 18387 21586
rect 15009 21528 15014 21584
rect 15070 21528 18326 21584
rect 18382 21528 18387 21584
rect 15009 21526 18387 21528
rect 15009 21523 15075 21526
rect 18321 21523 18387 21526
rect 22369 21586 22435 21589
rect 26200 21586 27000 21616
rect 22369 21584 27000 21586
rect 22369 21528 22374 21584
rect 22430 21528 27000 21584
rect 22369 21526 27000 21528
rect 22369 21523 22435 21526
rect 26200 21496 27000 21526
rect 3601 21450 3667 21453
rect 13169 21450 13235 21453
rect 3601 21448 13235 21450
rect 3601 21392 3606 21448
rect 3662 21392 13174 21448
rect 13230 21392 13235 21448
rect 3601 21390 13235 21392
rect 3601 21387 3667 21390
rect 13169 21387 13235 21390
rect 15561 21450 15627 21453
rect 18413 21450 18479 21453
rect 15561 21448 18479 21450
rect 15561 21392 15566 21448
rect 15622 21392 18418 21448
rect 18474 21392 18479 21448
rect 15561 21390 18479 21392
rect 15561 21387 15627 21390
rect 18413 21387 18479 21390
rect 22461 21450 22527 21453
rect 22461 21448 23490 21450
rect 22461 21392 22466 21448
rect 22522 21392 23490 21448
rect 22461 21390 23490 21392
rect 22461 21387 22527 21390
rect 12249 21314 12315 21317
rect 12709 21314 12775 21317
rect 12249 21312 12775 21314
rect 12249 21256 12254 21312
rect 12310 21256 12714 21312
rect 12770 21256 12775 21312
rect 12249 21254 12775 21256
rect 12249 21251 12315 21254
rect 12709 21251 12775 21254
rect 14549 21314 14615 21317
rect 17401 21314 17467 21317
rect 14549 21312 17467 21314
rect 14549 21256 14554 21312
rect 14610 21256 17406 21312
rect 17462 21256 17467 21312
rect 14549 21254 17467 21256
rect 14549 21251 14615 21254
rect 17401 21251 17467 21254
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 13813 21178 13879 21181
rect 17677 21178 17743 21181
rect 13813 21176 17743 21178
rect 13813 21120 13818 21176
rect 13874 21120 17682 21176
rect 17738 21120 17743 21176
rect 13813 21118 17743 21120
rect 23430 21178 23490 21390
rect 26200 21178 27000 21208
rect 23430 21118 27000 21178
rect 13813 21115 13879 21118
rect 17677 21115 17743 21118
rect 26200 21088 27000 21118
rect 11881 21042 11947 21045
rect 11881 21040 24226 21042
rect 11881 20984 11886 21040
rect 11942 20984 24226 21040
rect 11881 20982 24226 20984
rect 11881 20979 11947 20982
rect 4061 20906 4127 20909
rect 13261 20906 13327 20909
rect 4061 20904 13327 20906
rect 4061 20848 4066 20904
rect 4122 20848 13266 20904
rect 13322 20848 13327 20904
rect 4061 20846 13327 20848
rect 4061 20843 4127 20846
rect 13261 20843 13327 20846
rect 13721 20906 13787 20909
rect 13721 20904 16130 20906
rect 13721 20848 13726 20904
rect 13782 20848 16130 20904
rect 13721 20846 16130 20848
rect 13721 20843 13787 20846
rect 13537 20770 13603 20773
rect 13670 20770 13676 20772
rect 13537 20768 13676 20770
rect 13537 20712 13542 20768
rect 13598 20712 13676 20768
rect 13537 20710 13676 20712
rect 13537 20707 13603 20710
rect 13670 20708 13676 20710
rect 13740 20708 13746 20772
rect 16070 20770 16130 20846
rect 16430 20844 16436 20908
rect 16500 20906 16506 20908
rect 22645 20906 22711 20909
rect 16500 20904 22711 20906
rect 16500 20848 22650 20904
rect 22706 20848 22711 20904
rect 16500 20846 22711 20848
rect 16500 20844 16506 20846
rect 22645 20843 22711 20846
rect 16941 20770 17007 20773
rect 16070 20768 17007 20770
rect 16070 20712 16946 20768
rect 17002 20712 17007 20768
rect 16070 20710 17007 20712
rect 16941 20707 17007 20710
rect 22185 20770 22251 20773
rect 22318 20770 22324 20772
rect 22185 20768 22324 20770
rect 22185 20712 22190 20768
rect 22246 20712 22324 20768
rect 22185 20710 22324 20712
rect 22185 20707 22251 20710
rect 22318 20708 22324 20710
rect 22388 20708 22394 20772
rect 24166 20770 24226 20982
rect 26200 20770 27000 20800
rect 24166 20710 27000 20770
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 26200 20680 27000 20710
rect 17946 20639 18262 20640
rect 9305 20634 9371 20637
rect 12433 20634 12499 20637
rect 9305 20632 12499 20634
rect 9305 20576 9310 20632
rect 9366 20576 12438 20632
rect 12494 20576 12499 20632
rect 9305 20574 12499 20576
rect 9305 20571 9371 20574
rect 12433 20571 12499 20574
rect 15837 20636 15903 20637
rect 15837 20632 15884 20636
rect 15948 20634 15954 20636
rect 15837 20576 15842 20632
rect 15837 20572 15884 20576
rect 15948 20574 15994 20634
rect 15948 20572 15954 20574
rect 15837 20571 15903 20572
rect 11145 20498 11211 20501
rect 15929 20498 15995 20501
rect 11145 20496 15995 20498
rect 11145 20440 11150 20496
rect 11206 20440 15934 20496
rect 15990 20440 15995 20496
rect 11145 20438 15995 20440
rect 11145 20435 11211 20438
rect 15929 20435 15995 20438
rect 16665 20498 16731 20501
rect 19241 20498 19307 20501
rect 16665 20496 19307 20498
rect 16665 20440 16670 20496
rect 16726 20440 19246 20496
rect 19302 20440 19307 20496
rect 16665 20438 19307 20440
rect 16665 20435 16731 20438
rect 19241 20435 19307 20438
rect 20846 20436 20852 20500
rect 20916 20498 20922 20500
rect 21541 20498 21607 20501
rect 20916 20496 21607 20498
rect 20916 20440 21546 20496
rect 21602 20440 21607 20496
rect 20916 20438 21607 20440
rect 20916 20436 20922 20438
rect 21541 20435 21607 20438
rect 5533 20362 5599 20365
rect 15929 20362 15995 20365
rect 5533 20360 15995 20362
rect 5533 20304 5538 20360
rect 5594 20304 15934 20360
rect 15990 20304 15995 20360
rect 5533 20302 15995 20304
rect 5533 20299 5599 20302
rect 15929 20299 15995 20302
rect 16389 20362 16455 20365
rect 20713 20362 20779 20365
rect 26200 20362 27000 20392
rect 16389 20360 20779 20362
rect 16389 20304 16394 20360
rect 16450 20304 20718 20360
rect 20774 20304 20779 20360
rect 16389 20302 20779 20304
rect 16389 20299 16455 20302
rect 20713 20299 20779 20302
rect 22050 20302 27000 20362
rect 14733 20226 14799 20229
rect 22050 20226 22110 20302
rect 26200 20272 27000 20302
rect 14733 20224 22110 20226
rect 14733 20168 14738 20224
rect 14794 20168 22110 20224
rect 14733 20166 22110 20168
rect 14733 20163 14799 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 9305 20090 9371 20093
rect 11605 20090 11671 20093
rect 9305 20088 11671 20090
rect 9305 20032 9310 20088
rect 9366 20032 11610 20088
rect 11666 20032 11671 20088
rect 9305 20030 11671 20032
rect 9305 20027 9371 20030
rect 11605 20027 11671 20030
rect 14273 20090 14339 20093
rect 16481 20090 16547 20093
rect 14273 20088 16547 20090
rect 14273 20032 14278 20088
rect 14334 20032 16486 20088
rect 16542 20032 16547 20088
rect 14273 20030 16547 20032
rect 14273 20027 14339 20030
rect 16481 20027 16547 20030
rect 2221 19954 2287 19957
rect 16430 19954 16436 19956
rect 2221 19952 16436 19954
rect 2221 19896 2226 19952
rect 2282 19896 16436 19952
rect 2221 19894 16436 19896
rect 2221 19891 2287 19894
rect 16430 19892 16436 19894
rect 16500 19892 16506 19956
rect 19558 19892 19564 19956
rect 19628 19954 19634 19956
rect 22553 19954 22619 19957
rect 19628 19952 22619 19954
rect 19628 19896 22558 19952
rect 22614 19896 22619 19952
rect 19628 19894 22619 19896
rect 19628 19892 19634 19894
rect 22553 19891 22619 19894
rect 22737 19954 22803 19957
rect 26200 19954 27000 19984
rect 22737 19952 27000 19954
rect 22737 19896 22742 19952
rect 22798 19896 27000 19952
rect 22737 19894 27000 19896
rect 22737 19891 22803 19894
rect 26200 19864 27000 19894
rect 4521 19818 4587 19821
rect 20989 19818 21055 19821
rect 4521 19816 21055 19818
rect 4521 19760 4526 19816
rect 4582 19760 20994 19816
rect 21050 19760 21055 19816
rect 4521 19758 21055 19760
rect 4521 19755 4587 19758
rect 20989 19755 21055 19758
rect 16297 19682 16363 19685
rect 8342 19680 16363 19682
rect 8342 19624 16302 19680
rect 16358 19624 16363 19680
rect 8342 19622 16363 19624
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 2313 19410 2379 19413
rect 8342 19410 8402 19622
rect 16297 19619 16363 19622
rect 20662 19620 20668 19684
rect 20732 19682 20738 19684
rect 22461 19682 22527 19685
rect 20732 19680 22527 19682
rect 20732 19624 22466 19680
rect 22522 19624 22527 19680
rect 20732 19622 22527 19624
rect 20732 19620 20738 19622
rect 22461 19619 22527 19622
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 10317 19546 10383 19549
rect 16573 19546 16639 19549
rect 10317 19544 16639 19546
rect 10317 19488 10322 19544
rect 10378 19488 16578 19544
rect 16634 19488 16639 19544
rect 10317 19486 16639 19488
rect 10317 19483 10383 19486
rect 16573 19483 16639 19486
rect 21173 19546 21239 19549
rect 21817 19546 21883 19549
rect 21173 19544 21883 19546
rect 21173 19488 21178 19544
rect 21234 19488 21822 19544
rect 21878 19488 21883 19544
rect 21173 19486 21883 19488
rect 21173 19483 21239 19486
rect 21817 19483 21883 19486
rect 22001 19546 22067 19549
rect 22185 19546 22251 19549
rect 22001 19544 22251 19546
rect 22001 19488 22006 19544
rect 22062 19488 22190 19544
rect 22246 19488 22251 19544
rect 22001 19486 22251 19488
rect 22001 19483 22067 19486
rect 22185 19483 22251 19486
rect 23013 19546 23079 19549
rect 26200 19546 27000 19576
rect 23013 19544 27000 19546
rect 23013 19488 23018 19544
rect 23074 19488 27000 19544
rect 23013 19486 27000 19488
rect 23013 19483 23079 19486
rect 26200 19456 27000 19486
rect 2313 19408 8402 19410
rect 2313 19352 2318 19408
rect 2374 19352 8402 19408
rect 2313 19350 8402 19352
rect 8569 19410 8635 19413
rect 10777 19410 10843 19413
rect 8569 19408 10843 19410
rect 8569 19352 8574 19408
rect 8630 19352 10782 19408
rect 10838 19352 10843 19408
rect 8569 19350 10843 19352
rect 2313 19347 2379 19350
rect 8569 19347 8635 19350
rect 10777 19347 10843 19350
rect 12801 19410 12867 19413
rect 14733 19410 14799 19413
rect 12801 19408 14799 19410
rect 12801 19352 12806 19408
rect 12862 19352 14738 19408
rect 14794 19352 14799 19408
rect 12801 19350 14799 19352
rect 12801 19347 12867 19350
rect 14733 19347 14799 19350
rect 15142 19348 15148 19412
rect 15212 19410 15218 19412
rect 15285 19410 15351 19413
rect 15212 19408 15351 19410
rect 15212 19352 15290 19408
rect 15346 19352 15351 19408
rect 15212 19350 15351 19352
rect 15212 19348 15218 19350
rect 15285 19347 15351 19350
rect 15837 19410 15903 19413
rect 16062 19410 16068 19412
rect 15837 19408 16068 19410
rect 15837 19352 15842 19408
rect 15898 19352 16068 19408
rect 15837 19350 16068 19352
rect 15837 19347 15903 19350
rect 16062 19348 16068 19350
rect 16132 19348 16138 19412
rect 16430 19348 16436 19412
rect 16500 19410 16506 19412
rect 23105 19410 23171 19413
rect 16500 19408 23171 19410
rect 16500 19352 23110 19408
rect 23166 19352 23171 19408
rect 16500 19350 23171 19352
rect 16500 19348 16506 19350
rect 23105 19347 23171 19350
rect 4705 19274 4771 19277
rect 22829 19274 22895 19277
rect 4705 19272 22895 19274
rect 4705 19216 4710 19272
rect 4766 19216 22834 19272
rect 22890 19216 22895 19272
rect 4705 19214 22895 19216
rect 4705 19211 4771 19214
rect 22829 19211 22895 19214
rect 7741 19138 7807 19141
rect 11881 19138 11947 19141
rect 7741 19136 11947 19138
rect 7741 19080 7746 19136
rect 7802 19080 11886 19136
rect 11942 19080 11947 19136
rect 7741 19078 11947 19080
rect 7741 19075 7807 19078
rect 11881 19075 11947 19078
rect 21030 19076 21036 19140
rect 21100 19138 21106 19140
rect 22093 19138 22159 19141
rect 21100 19136 22159 19138
rect 21100 19080 22098 19136
rect 22154 19080 22159 19136
rect 21100 19078 22159 19080
rect 21100 19076 21106 19078
rect 22093 19075 22159 19078
rect 23381 19138 23447 19141
rect 26200 19138 27000 19168
rect 23381 19136 27000 19138
rect 23381 19080 23386 19136
rect 23442 19080 27000 19136
rect 23381 19078 27000 19080
rect 23381 19075 23447 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 26200 19048 27000 19078
rect 22946 19007 23262 19008
rect 7557 19002 7623 19005
rect 9673 19002 9739 19005
rect 7557 19000 9739 19002
rect 7557 18944 7562 19000
rect 7618 18944 9678 19000
rect 9734 18944 9739 19000
rect 7557 18942 9739 18944
rect 7557 18939 7623 18942
rect 9673 18939 9739 18942
rect 13905 19002 13971 19005
rect 17125 19002 17191 19005
rect 13905 19000 17191 19002
rect 13905 18944 13910 19000
rect 13966 18944 17130 19000
rect 17186 18944 17191 19000
rect 13905 18942 17191 18944
rect 13905 18939 13971 18942
rect 17125 18939 17191 18942
rect 19701 19002 19767 19005
rect 22737 19002 22803 19005
rect 19701 19000 22803 19002
rect 19701 18944 19706 19000
rect 19762 18944 22742 19000
rect 22798 18944 22803 19000
rect 19701 18942 22803 18944
rect 19701 18939 19767 18942
rect 22737 18939 22803 18942
rect 1577 18866 1643 18869
rect 13721 18866 13787 18869
rect 1577 18864 13787 18866
rect 1577 18808 1582 18864
rect 1638 18808 13726 18864
rect 13782 18808 13787 18864
rect 1577 18806 13787 18808
rect 1577 18803 1643 18806
rect 13721 18803 13787 18806
rect 16205 18866 16271 18869
rect 16614 18866 16620 18868
rect 16205 18864 16620 18866
rect 16205 18808 16210 18864
rect 16266 18808 16620 18864
rect 16205 18806 16620 18808
rect 16205 18803 16271 18806
rect 16614 18804 16620 18806
rect 16684 18804 16690 18868
rect 18045 18866 18111 18869
rect 19006 18866 19012 18868
rect 18045 18864 19012 18866
rect 18045 18808 18050 18864
rect 18106 18808 19012 18864
rect 18045 18806 19012 18808
rect 18045 18803 18111 18806
rect 19006 18804 19012 18806
rect 19076 18804 19082 18868
rect 22686 18804 22692 18868
rect 22756 18866 22762 18868
rect 24853 18866 24919 18869
rect 22756 18864 24919 18866
rect 22756 18808 24858 18864
rect 24914 18808 24919 18864
rect 22756 18806 24919 18808
rect 22756 18804 22762 18806
rect 24853 18803 24919 18806
rect 5165 18730 5231 18733
rect 23013 18730 23079 18733
rect 26200 18730 27000 18760
rect 5165 18728 23079 18730
rect 5165 18672 5170 18728
rect 5226 18672 23018 18728
rect 23074 18672 23079 18728
rect 5165 18670 23079 18672
rect 5165 18667 5231 18670
rect 23013 18667 23079 18670
rect 23246 18670 27000 18730
rect 11329 18594 11395 18597
rect 16573 18594 16639 18597
rect 11329 18592 16639 18594
rect 11329 18536 11334 18592
rect 11390 18536 16578 18592
rect 16634 18536 16639 18592
rect 11329 18534 16639 18536
rect 11329 18531 11395 18534
rect 16573 18531 16639 18534
rect 22277 18594 22343 18597
rect 23246 18594 23306 18670
rect 26200 18640 27000 18670
rect 22277 18592 23306 18594
rect 22277 18536 22282 18592
rect 22338 18536 23306 18592
rect 22277 18534 23306 18536
rect 22277 18531 22343 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 10409 18458 10475 18461
rect 16481 18458 16547 18461
rect 10409 18456 16547 18458
rect 10409 18400 10414 18456
rect 10470 18400 16486 18456
rect 16542 18400 16547 18456
rect 10409 18398 16547 18400
rect 10409 18395 10475 18398
rect 16481 18395 16547 18398
rect 9213 18322 9279 18325
rect 20897 18322 20963 18325
rect 9213 18320 20963 18322
rect 9213 18264 9218 18320
rect 9274 18264 20902 18320
rect 20958 18264 20963 18320
rect 9213 18262 20963 18264
rect 9213 18259 9279 18262
rect 20897 18259 20963 18262
rect 23105 18322 23171 18325
rect 26200 18322 27000 18352
rect 23105 18320 27000 18322
rect 23105 18264 23110 18320
rect 23166 18264 27000 18320
rect 23105 18262 27000 18264
rect 23105 18259 23171 18262
rect 26200 18232 27000 18262
rect 5625 18186 5691 18189
rect 24393 18186 24459 18189
rect 5625 18184 24459 18186
rect 5625 18128 5630 18184
rect 5686 18128 24398 18184
rect 24454 18128 24459 18184
rect 5625 18126 24459 18128
rect 5625 18123 5691 18126
rect 24393 18123 24459 18126
rect 7465 18050 7531 18053
rect 7741 18050 7807 18053
rect 7465 18048 7807 18050
rect 7465 17992 7470 18048
rect 7526 17992 7746 18048
rect 7802 17992 7807 18048
rect 7465 17990 7807 17992
rect 7465 17987 7531 17990
rect 7741 17987 7807 17990
rect 14273 18050 14339 18053
rect 19701 18050 19767 18053
rect 14273 18048 19767 18050
rect 14273 17992 14278 18048
rect 14334 17992 19706 18048
rect 19762 17992 19767 18048
rect 14273 17990 19767 17992
rect 14273 17987 14339 17990
rect 19701 17987 19767 17990
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 6453 17914 6519 17917
rect 9397 17914 9463 17917
rect 6453 17912 9463 17914
rect 6453 17856 6458 17912
rect 6514 17856 9402 17912
rect 9458 17856 9463 17912
rect 6453 17854 9463 17856
rect 6453 17851 6519 17854
rect 9397 17851 9463 17854
rect 11973 17914 12039 17917
rect 15837 17914 15903 17917
rect 17217 17914 17283 17917
rect 19793 17914 19859 17917
rect 26200 17914 27000 17944
rect 11973 17912 12864 17914
rect 11973 17856 11978 17912
rect 12034 17856 12864 17912
rect 11973 17854 12864 17856
rect 11973 17851 12039 17854
rect 4705 17778 4771 17781
rect 4838 17778 4844 17780
rect 4705 17776 4844 17778
rect 4705 17720 4710 17776
rect 4766 17720 4844 17776
rect 4705 17718 4844 17720
rect 4705 17715 4771 17718
rect 4838 17716 4844 17718
rect 4908 17716 4914 17780
rect 7833 17778 7899 17781
rect 12617 17778 12683 17781
rect 7833 17776 12683 17778
rect 7833 17720 7838 17776
rect 7894 17720 12622 17776
rect 12678 17720 12683 17776
rect 7833 17718 12683 17720
rect 12804 17778 12864 17854
rect 15837 17912 17283 17914
rect 15837 17856 15842 17912
rect 15898 17856 17222 17912
rect 17278 17856 17283 17912
rect 15837 17854 17283 17856
rect 15837 17851 15903 17854
rect 17217 17851 17283 17854
rect 17358 17912 19859 17914
rect 17358 17856 19798 17912
rect 19854 17856 19859 17912
rect 17358 17854 19859 17856
rect 15101 17778 15167 17781
rect 12804 17776 15167 17778
rect 12804 17720 15106 17776
rect 15162 17720 15167 17776
rect 12804 17718 15167 17720
rect 7833 17715 7899 17718
rect 12617 17715 12683 17718
rect 15101 17715 15167 17718
rect 15469 17778 15535 17781
rect 17358 17778 17418 17854
rect 19793 17851 19859 17854
rect 23430 17854 27000 17914
rect 15469 17776 17418 17778
rect 15469 17720 15474 17776
rect 15530 17720 17418 17776
rect 15469 17718 17418 17720
rect 15469 17715 15535 17718
rect 19374 17716 19380 17780
rect 19444 17778 19450 17780
rect 19793 17778 19859 17781
rect 19444 17776 19859 17778
rect 19444 17720 19798 17776
rect 19854 17720 19859 17776
rect 19444 17718 19859 17720
rect 19444 17716 19450 17718
rect 19793 17715 19859 17718
rect 23013 17778 23079 17781
rect 23430 17778 23490 17854
rect 26200 17824 27000 17854
rect 23013 17776 23490 17778
rect 23013 17720 23018 17776
rect 23074 17720 23490 17776
rect 23013 17718 23490 17720
rect 23013 17715 23079 17718
rect 7189 17642 7255 17645
rect 8845 17642 8911 17645
rect 24485 17642 24551 17645
rect 7189 17640 8402 17642
rect 7189 17584 7194 17640
rect 7250 17584 8402 17640
rect 7189 17582 8402 17584
rect 7189 17579 7255 17582
rect 8342 17506 8402 17582
rect 8845 17640 24551 17642
rect 8845 17584 8850 17640
rect 8906 17584 24490 17640
rect 24546 17584 24551 17640
rect 8845 17582 24551 17584
rect 8845 17579 8911 17582
rect 24485 17579 24551 17582
rect 15142 17506 15148 17508
rect 8342 17446 15148 17506
rect 15142 17444 15148 17446
rect 15212 17444 15218 17508
rect 15653 17506 15719 17509
rect 16205 17506 16271 17509
rect 15653 17504 16271 17506
rect 15653 17448 15658 17504
rect 15714 17448 16210 17504
rect 16266 17448 16271 17504
rect 15653 17446 16271 17448
rect 15653 17443 15719 17446
rect 16205 17443 16271 17446
rect 22093 17506 22159 17509
rect 26200 17506 27000 17536
rect 22093 17504 27000 17506
rect 22093 17448 22098 17504
rect 22154 17448 27000 17504
rect 22093 17446 27000 17448
rect 22093 17443 22159 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 26200 17416 27000 17446
rect 17946 17375 18262 17376
rect 22461 17372 22527 17373
rect 16798 17370 16804 17372
rect 8342 17310 16804 17370
rect 5533 17234 5599 17237
rect 8342 17234 8402 17310
rect 16798 17308 16804 17310
rect 16868 17308 16874 17372
rect 22461 17368 22508 17372
rect 22572 17370 22578 17372
rect 22461 17312 22466 17368
rect 22461 17308 22508 17312
rect 22572 17310 22618 17370
rect 22572 17308 22578 17310
rect 22461 17307 22527 17308
rect 5533 17232 8402 17234
rect 5533 17176 5538 17232
rect 5594 17176 8402 17232
rect 5533 17174 8402 17176
rect 9397 17234 9463 17237
rect 24853 17234 24919 17237
rect 9397 17232 24919 17234
rect 9397 17176 9402 17232
rect 9458 17176 24858 17232
rect 24914 17176 24919 17232
rect 9397 17174 24919 17176
rect 5533 17171 5599 17174
rect 9397 17171 9463 17174
rect 24853 17171 24919 17174
rect 7097 17098 7163 17101
rect 16430 17098 16436 17100
rect 7097 17096 16436 17098
rect 7097 17040 7102 17096
rect 7158 17040 16436 17096
rect 7097 17038 16436 17040
rect 7097 17035 7163 17038
rect 16430 17036 16436 17038
rect 16500 17036 16506 17100
rect 17217 17098 17283 17101
rect 18137 17098 18203 17101
rect 17217 17096 18203 17098
rect 17217 17040 17222 17096
rect 17278 17040 18142 17096
rect 18198 17040 18203 17096
rect 17217 17038 18203 17040
rect 17217 17035 17283 17038
rect 18137 17035 18203 17038
rect 18321 17098 18387 17101
rect 18965 17098 19031 17101
rect 18321 17096 19031 17098
rect 18321 17040 18326 17096
rect 18382 17040 18970 17096
rect 19026 17040 19031 17096
rect 18321 17038 19031 17040
rect 18321 17035 18387 17038
rect 18965 17035 19031 17038
rect 22461 17098 22527 17101
rect 23013 17098 23079 17101
rect 22461 17096 23079 17098
rect 22461 17040 22466 17096
rect 22522 17040 23018 17096
rect 23074 17040 23079 17096
rect 22461 17038 23079 17040
rect 22461 17035 22527 17038
rect 23013 17035 23079 17038
rect 23422 17036 23428 17100
rect 23492 17098 23498 17100
rect 26200 17098 27000 17128
rect 23492 17038 27000 17098
rect 23492 17036 23498 17038
rect 26200 17008 27000 17038
rect 10041 16962 10107 16965
rect 11605 16962 11671 16965
rect 10041 16960 11671 16962
rect 10041 16904 10046 16960
rect 10102 16904 11610 16960
rect 11666 16904 11671 16960
rect 10041 16902 11671 16904
rect 10041 16899 10107 16902
rect 11605 16899 11671 16902
rect 11881 16962 11947 16965
rect 12617 16962 12683 16965
rect 11881 16960 12683 16962
rect 11881 16904 11886 16960
rect 11942 16904 12622 16960
rect 12678 16904 12683 16960
rect 11881 16902 12683 16904
rect 11881 16899 11947 16902
rect 12617 16899 12683 16902
rect 16297 16962 16363 16965
rect 22093 16962 22159 16965
rect 16297 16960 22159 16962
rect 16297 16904 16302 16960
rect 16358 16904 22098 16960
rect 22154 16904 22159 16960
rect 16297 16902 22159 16904
rect 16297 16899 16363 16902
rect 22093 16899 22159 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 9305 16826 9371 16829
rect 10409 16826 10475 16829
rect 19425 16828 19491 16829
rect 19374 16826 19380 16828
rect 9305 16824 10475 16826
rect 9305 16768 9310 16824
rect 9366 16768 10414 16824
rect 10470 16768 10475 16824
rect 9305 16766 10475 16768
rect 19334 16766 19380 16826
rect 19444 16824 19491 16828
rect 19486 16768 19491 16824
rect 9305 16763 9371 16766
rect 10409 16763 10475 16766
rect 19374 16764 19380 16766
rect 19444 16764 19491 16768
rect 19425 16763 19491 16764
rect 5257 16690 5323 16693
rect 13261 16690 13327 16693
rect 5257 16688 13327 16690
rect 5257 16632 5262 16688
rect 5318 16632 13266 16688
rect 13322 16632 13327 16688
rect 5257 16630 13327 16632
rect 5257 16627 5323 16630
rect 13261 16627 13327 16630
rect 13445 16690 13511 16693
rect 15193 16690 15259 16693
rect 13445 16688 15259 16690
rect 13445 16632 13450 16688
rect 13506 16632 15198 16688
rect 15254 16632 15259 16688
rect 13445 16630 15259 16632
rect 13445 16627 13511 16630
rect 15193 16627 15259 16630
rect 17493 16690 17559 16693
rect 17718 16690 17724 16692
rect 17493 16688 17724 16690
rect 17493 16632 17498 16688
rect 17554 16632 17724 16688
rect 17493 16630 17724 16632
rect 17493 16627 17559 16630
rect 17718 16628 17724 16630
rect 17788 16628 17794 16692
rect 21909 16690 21975 16693
rect 26200 16690 27000 16720
rect 21909 16688 27000 16690
rect 21909 16632 21914 16688
rect 21970 16632 27000 16688
rect 21909 16630 27000 16632
rect 21909 16627 21975 16630
rect 26200 16600 27000 16630
rect 10317 16554 10383 16557
rect 19558 16554 19564 16556
rect 10317 16552 19564 16554
rect 10317 16496 10322 16552
rect 10378 16496 19564 16552
rect 10317 16494 19564 16496
rect 10317 16491 10383 16494
rect 19558 16492 19564 16494
rect 19628 16492 19634 16556
rect 8753 16418 8819 16421
rect 12801 16418 12867 16421
rect 8753 16416 12867 16418
rect 8753 16360 8758 16416
rect 8814 16360 12806 16416
rect 12862 16360 12867 16416
rect 8753 16358 12867 16360
rect 8753 16355 8819 16358
rect 12801 16355 12867 16358
rect 18454 16356 18460 16420
rect 18524 16418 18530 16420
rect 24669 16418 24735 16421
rect 18524 16416 24735 16418
rect 18524 16360 24674 16416
rect 24730 16360 24735 16416
rect 18524 16358 24735 16360
rect 18524 16356 18530 16358
rect 24669 16355 24735 16358
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 9765 16282 9831 16285
rect 10225 16282 10291 16285
rect 9765 16280 10291 16282
rect 9765 16224 9770 16280
rect 9826 16224 10230 16280
rect 10286 16224 10291 16280
rect 9765 16222 10291 16224
rect 9765 16219 9831 16222
rect 10225 16219 10291 16222
rect 23473 16282 23539 16285
rect 26200 16282 27000 16312
rect 23473 16280 27000 16282
rect 23473 16224 23478 16280
rect 23534 16224 27000 16280
rect 23473 16222 27000 16224
rect 23473 16219 23539 16222
rect 26200 16192 27000 16222
rect 8661 16146 8727 16149
rect 24526 16146 24532 16148
rect 8661 16144 24532 16146
rect 8661 16088 8666 16144
rect 8722 16088 24532 16144
rect 8661 16086 24532 16088
rect 8661 16083 8727 16086
rect 24526 16084 24532 16086
rect 24596 16084 24602 16148
rect 9121 16010 9187 16013
rect 22686 16010 22692 16012
rect 9121 16008 22692 16010
rect 9121 15952 9126 16008
rect 9182 15952 22692 16008
rect 9121 15950 22692 15952
rect 9121 15947 9187 15950
rect 22686 15948 22692 15950
rect 22756 15948 22762 16012
rect 9673 15874 9739 15877
rect 12249 15874 12315 15877
rect 9673 15872 12315 15874
rect 9673 15816 9678 15872
rect 9734 15816 12254 15872
rect 12310 15816 12315 15872
rect 9673 15814 12315 15816
rect 9673 15811 9739 15814
rect 12249 15811 12315 15814
rect 24761 15874 24827 15877
rect 26200 15874 27000 15904
rect 24761 15872 27000 15874
rect 24761 15816 24766 15872
rect 24822 15816 27000 15872
rect 24761 15814 27000 15816
rect 24761 15811 24827 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 26200 15784 27000 15814
rect 22946 15743 23262 15744
rect 14641 15738 14707 15741
rect 19149 15738 19215 15741
rect 14641 15736 19215 15738
rect 14641 15680 14646 15736
rect 14702 15680 19154 15736
rect 19210 15680 19215 15736
rect 14641 15678 19215 15680
rect 14641 15675 14707 15678
rect 19149 15675 19215 15678
rect 20161 15738 20227 15741
rect 20161 15736 22754 15738
rect 20161 15680 20166 15736
rect 20222 15680 22754 15736
rect 20161 15678 22754 15680
rect 20161 15675 20227 15678
rect 10041 15602 10107 15605
rect 22134 15602 22140 15604
rect 10041 15600 22140 15602
rect 10041 15544 10046 15600
rect 10102 15544 22140 15600
rect 10041 15542 22140 15544
rect 10041 15539 10107 15542
rect 22134 15540 22140 15542
rect 22204 15540 22210 15604
rect 13905 15466 13971 15469
rect 22461 15466 22527 15469
rect 13905 15464 22527 15466
rect 13905 15408 13910 15464
rect 13966 15408 22466 15464
rect 22522 15408 22527 15464
rect 13905 15406 22527 15408
rect 22694 15466 22754 15678
rect 26200 15466 27000 15496
rect 22694 15406 27000 15466
rect 13905 15403 13971 15406
rect 22461 15403 22527 15406
rect 26200 15376 27000 15406
rect 18413 15330 18479 15333
rect 22318 15330 22324 15332
rect 18413 15328 22324 15330
rect 18413 15272 18418 15328
rect 18474 15272 22324 15328
rect 18413 15270 22324 15272
rect 18413 15267 18479 15270
rect 22318 15268 22324 15270
rect 22388 15268 22394 15332
rect 22686 15268 22692 15332
rect 22756 15330 22762 15332
rect 22829 15330 22895 15333
rect 22756 15328 22895 15330
rect 22756 15272 22834 15328
rect 22890 15272 22895 15328
rect 22756 15270 22895 15272
rect 22756 15268 22762 15270
rect 22829 15267 22895 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 23933 15194 23999 15197
rect 22050 15192 23999 15194
rect 22050 15136 23938 15192
rect 23994 15136 23999 15192
rect 22050 15134 23999 15136
rect 7649 15058 7715 15061
rect 22050 15058 22110 15134
rect 23933 15131 23999 15134
rect 7649 15056 22110 15058
rect 7649 15000 7654 15056
rect 7710 15000 22110 15056
rect 7649 14998 22110 15000
rect 22737 15058 22803 15061
rect 26200 15058 27000 15088
rect 22737 15056 27000 15058
rect 22737 15000 22742 15056
rect 22798 15000 27000 15056
rect 22737 14998 27000 15000
rect 7649 14995 7715 14998
rect 22737 14995 22803 14998
rect 26200 14968 27000 14998
rect 14825 14922 14891 14925
rect 20662 14922 20668 14924
rect 14825 14920 20668 14922
rect 14825 14864 14830 14920
rect 14886 14864 20668 14920
rect 14825 14862 20668 14864
rect 14825 14859 14891 14862
rect 20662 14860 20668 14862
rect 20732 14860 20738 14924
rect 13445 14786 13511 14789
rect 19742 14786 19748 14788
rect 13445 14784 19748 14786
rect 13445 14728 13450 14784
rect 13506 14728 19748 14784
rect 13445 14726 19748 14728
rect 13445 14723 13511 14726
rect 19742 14724 19748 14726
rect 19812 14724 19818 14788
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 13445 14650 13511 14653
rect 18638 14650 18644 14652
rect 13445 14648 18644 14650
rect 13445 14592 13450 14648
rect 13506 14592 18644 14648
rect 13445 14590 18644 14592
rect 13445 14587 13511 14590
rect 18638 14588 18644 14590
rect 18708 14588 18714 14652
rect 18822 14588 18828 14652
rect 18892 14650 18898 14652
rect 19057 14650 19123 14653
rect 26200 14650 27000 14680
rect 18892 14648 19123 14650
rect 18892 14592 19062 14648
rect 19118 14592 19123 14648
rect 18892 14590 19123 14592
rect 18892 14588 18898 14590
rect 19057 14587 19123 14590
rect 23384 14590 27000 14650
rect 4613 14514 4679 14517
rect 20069 14514 20135 14517
rect 4613 14512 20135 14514
rect 4613 14456 4618 14512
rect 4674 14456 20074 14512
rect 20130 14456 20135 14512
rect 4613 14454 20135 14456
rect 4613 14451 4679 14454
rect 20069 14451 20135 14454
rect 21541 14514 21607 14517
rect 23384 14514 23444 14590
rect 26200 14560 27000 14590
rect 21541 14512 23444 14514
rect 21541 14456 21546 14512
rect 21602 14456 23444 14512
rect 21541 14454 23444 14456
rect 21541 14451 21607 14454
rect 11881 14378 11947 14381
rect 18413 14378 18479 14381
rect 11881 14376 18479 14378
rect 11881 14320 11886 14376
rect 11942 14320 18418 14376
rect 18474 14320 18479 14376
rect 11881 14318 18479 14320
rect 11881 14315 11947 14318
rect 18413 14315 18479 14318
rect 18822 14316 18828 14380
rect 18892 14378 18898 14380
rect 18965 14378 19031 14381
rect 18892 14376 19031 14378
rect 18892 14320 18970 14376
rect 19026 14320 19031 14376
rect 18892 14318 19031 14320
rect 18892 14316 18898 14318
rect 18965 14315 19031 14318
rect 18873 14242 18939 14245
rect 19609 14242 19675 14245
rect 18873 14240 19675 14242
rect 18873 14184 18878 14240
rect 18934 14184 19614 14240
rect 19670 14184 19675 14240
rect 18873 14182 19675 14184
rect 18873 14179 18939 14182
rect 19609 14179 19675 14182
rect 23289 14242 23355 14245
rect 26200 14242 27000 14272
rect 23289 14240 27000 14242
rect 23289 14184 23294 14240
rect 23350 14184 27000 14240
rect 23289 14182 27000 14184
rect 23289 14179 23355 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 26200 14152 27000 14182
rect 17946 14111 18262 14112
rect 13353 14106 13419 14109
rect 17677 14106 17743 14109
rect 13353 14104 17743 14106
rect 13353 14048 13358 14104
rect 13414 14048 17682 14104
rect 17738 14048 17743 14104
rect 13353 14046 17743 14048
rect 13353 14043 13419 14046
rect 17677 14043 17743 14046
rect 6545 13970 6611 13973
rect 22093 13970 22159 13973
rect 6545 13968 22159 13970
rect 6545 13912 6550 13968
rect 6606 13912 22098 13968
rect 22154 13912 22159 13968
rect 6545 13910 22159 13912
rect 6545 13907 6611 13910
rect 22093 13907 22159 13910
rect 22737 13834 22803 13837
rect 26200 13834 27000 13864
rect 22737 13832 27000 13834
rect 22737 13776 22742 13832
rect 22798 13776 27000 13832
rect 22737 13774 27000 13776
rect 22737 13771 22803 13774
rect 26200 13744 27000 13774
rect 15653 13698 15719 13701
rect 20110 13698 20116 13700
rect 15653 13696 20116 13698
rect 15653 13640 15658 13696
rect 15714 13640 20116 13696
rect 15653 13638 20116 13640
rect 15653 13635 15719 13638
rect 20110 13636 20116 13638
rect 20180 13636 20186 13700
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 15101 13562 15167 13565
rect 19374 13562 19380 13564
rect 15101 13560 19380 13562
rect 15101 13504 15106 13560
rect 15162 13504 19380 13560
rect 15101 13502 19380 13504
rect 15101 13499 15167 13502
rect 19374 13500 19380 13502
rect 19444 13500 19450 13564
rect 23381 13426 23447 13429
rect 26200 13426 27000 13456
rect 23381 13424 27000 13426
rect 23381 13368 23386 13424
rect 23442 13368 27000 13424
rect 23381 13366 27000 13368
rect 23381 13363 23447 13366
rect 26200 13336 27000 13366
rect 19057 13292 19123 13293
rect 19006 13228 19012 13292
rect 19076 13290 19123 13292
rect 19076 13288 19168 13290
rect 19118 13232 19168 13288
rect 19076 13230 19168 13232
rect 19076 13228 19123 13230
rect 19057 13227 19123 13228
rect 22277 13154 22343 13157
rect 22737 13154 22803 13157
rect 22277 13152 22803 13154
rect 22277 13096 22282 13152
rect 22338 13096 22742 13152
rect 22798 13096 22803 13152
rect 22277 13094 22803 13096
rect 22277 13091 22343 13094
rect 22737 13091 22803 13094
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 26200 13018 27000 13048
rect 22188 12958 27000 13018
rect 22188 12885 22248 12958
rect 26200 12928 27000 12958
rect 4521 12882 4587 12885
rect 18454 12882 18460 12884
rect 4521 12880 18460 12882
rect 4521 12824 4526 12880
rect 4582 12824 18460 12880
rect 4521 12822 18460 12824
rect 4521 12819 4587 12822
rect 18454 12820 18460 12822
rect 18524 12820 18530 12884
rect 22185 12880 22251 12885
rect 22185 12824 22190 12880
rect 22246 12824 22251 12880
rect 22185 12819 22251 12824
rect 22461 12882 22527 12885
rect 23422 12882 23428 12884
rect 22461 12880 23428 12882
rect 22461 12824 22466 12880
rect 22522 12824 23428 12880
rect 22461 12822 23428 12824
rect 22461 12819 22527 12822
rect 23422 12820 23428 12822
rect 23492 12820 23498 12884
rect 12801 12746 12867 12749
rect 24209 12746 24275 12749
rect 12801 12744 24275 12746
rect 12801 12688 12806 12744
rect 12862 12688 24214 12744
rect 24270 12688 24275 12744
rect 12801 12686 24275 12688
rect 12801 12683 12867 12686
rect 24209 12683 24275 12686
rect 18321 12610 18387 12613
rect 20846 12610 20852 12612
rect 18321 12608 20852 12610
rect 18321 12552 18326 12608
rect 18382 12552 20852 12608
rect 18321 12550 20852 12552
rect 18321 12547 18387 12550
rect 20846 12548 20852 12550
rect 20916 12548 20922 12612
rect 24761 12610 24827 12613
rect 26200 12610 27000 12640
rect 24761 12608 27000 12610
rect 24761 12552 24766 12608
rect 24822 12552 27000 12608
rect 24761 12550 27000 12552
rect 24761 12547 24827 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 26200 12520 27000 12550
rect 22946 12479 23262 12480
rect 22277 12338 22343 12341
rect 22502 12338 22508 12340
rect 22277 12336 22508 12338
rect 22277 12280 22282 12336
rect 22338 12280 22508 12336
rect 22277 12278 22508 12280
rect 22277 12275 22343 12278
rect 22502 12276 22508 12278
rect 22572 12276 22578 12340
rect 5533 12202 5599 12205
rect 18689 12202 18755 12205
rect 5533 12200 18755 12202
rect 5533 12144 5538 12200
rect 5594 12144 18694 12200
rect 18750 12144 18755 12200
rect 5533 12142 18755 12144
rect 5533 12139 5599 12142
rect 18689 12139 18755 12142
rect 24669 12202 24735 12205
rect 26200 12202 27000 12232
rect 24669 12200 27000 12202
rect 24669 12144 24674 12200
rect 24730 12144 27000 12200
rect 24669 12142 27000 12144
rect 24669 12139 24735 12142
rect 26200 12112 27000 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 24853 11794 24919 11797
rect 26200 11794 27000 11824
rect 24853 11792 27000 11794
rect 24853 11736 24858 11792
rect 24914 11736 27000 11792
rect 24853 11734 27000 11736
rect 24853 11731 24919 11734
rect 26200 11704 27000 11734
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 20989 11388 21055 11389
rect 20989 11386 21036 11388
rect 20944 11384 21036 11386
rect 20944 11328 20994 11384
rect 20944 11326 21036 11328
rect 20989 11324 21036 11326
rect 21100 11324 21106 11388
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 20989 11323 21055 11324
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 16113 11250 16179 11253
rect 25957 11250 26023 11253
rect 16113 11248 26023 11250
rect 16113 11192 16118 11248
rect 16174 11192 25962 11248
rect 26018 11192 26023 11248
rect 16113 11190 26023 11192
rect 16113 11187 16179 11190
rect 25957 11187 26023 11190
rect 9438 11052 9444 11116
rect 9508 11114 9514 11116
rect 19701 11114 19767 11117
rect 9508 11112 19767 11114
rect 9508 11056 19706 11112
rect 19762 11056 19767 11112
rect 9508 11054 19767 11056
rect 9508 11052 9514 11054
rect 19701 11051 19767 11054
rect 24761 10978 24827 10981
rect 26200 10978 27000 11008
rect 24761 10976 27000 10978
rect 24761 10920 24766 10976
rect 24822 10920 27000 10976
rect 24761 10918 27000 10920
rect 24761 10915 24827 10918
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 26200 10888 27000 10918
rect 17946 10847 18262 10848
rect 24853 10570 24919 10573
rect 26200 10570 27000 10600
rect 24853 10568 27000 10570
rect 24853 10512 24858 10568
rect 24914 10512 27000 10568
rect 24853 10510 27000 10512
rect 24853 10507 24919 10510
rect 26200 10480 27000 10510
rect 16062 10372 16068 10436
rect 16132 10434 16138 10436
rect 20713 10434 20779 10437
rect 16132 10432 20779 10434
rect 16132 10376 20718 10432
rect 20774 10376 20779 10432
rect 16132 10374 20779 10376
rect 16132 10372 16138 10374
rect 20713 10371 20779 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 17534 10236 17540 10300
rect 17604 10298 17610 10300
rect 19425 10298 19491 10301
rect 17604 10296 19491 10298
rect 17604 10240 19430 10296
rect 19486 10240 19491 10296
rect 17604 10238 19491 10240
rect 17604 10236 17610 10238
rect 19425 10235 19491 10238
rect 24669 10162 24735 10165
rect 26200 10162 27000 10192
rect 24669 10160 27000 10162
rect 24669 10104 24674 10160
rect 24730 10104 27000 10160
rect 24669 10102 27000 10104
rect 24669 10099 24735 10102
rect 26200 10072 27000 10102
rect 16614 9964 16620 10028
rect 16684 10026 16690 10028
rect 19241 10026 19307 10029
rect 16684 10024 19307 10026
rect 16684 9968 19246 10024
rect 19302 9968 19307 10024
rect 16684 9966 19307 9968
rect 16684 9964 16690 9966
rect 19241 9963 19307 9966
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 23289 9754 23355 9757
rect 26200 9754 27000 9784
rect 23289 9752 27000 9754
rect 23289 9696 23294 9752
rect 23350 9696 27000 9752
rect 23289 9694 27000 9696
rect 23289 9691 23355 9694
rect 26200 9664 27000 9694
rect 15878 9420 15884 9484
rect 15948 9482 15954 9484
rect 19425 9482 19491 9485
rect 15948 9480 19491 9482
rect 15948 9424 19430 9480
rect 19486 9424 19491 9480
rect 15948 9422 19491 9424
rect 15948 9420 15954 9422
rect 19425 9419 19491 9422
rect 24853 9346 24919 9349
rect 26200 9346 27000 9376
rect 24853 9344 27000 9346
rect 24853 9288 24858 9344
rect 24914 9288 27000 9344
rect 24853 9286 27000 9288
rect 24853 9283 24919 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 26200 9256 27000 9286
rect 22946 9215 23262 9216
rect 25129 8938 25195 8941
rect 26200 8938 27000 8968
rect 25129 8936 27000 8938
rect 25129 8880 25134 8936
rect 25190 8880 27000 8936
rect 25129 8878 27000 8880
rect 25129 8875 25195 8878
rect 26200 8848 27000 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 24945 8530 25011 8533
rect 26200 8530 27000 8560
rect 24945 8528 27000 8530
rect 24945 8472 24950 8528
rect 25006 8472 27000 8528
rect 24945 8470 27000 8472
rect 24945 8467 25011 8470
rect 26200 8440 27000 8470
rect 13670 8332 13676 8396
rect 13740 8394 13746 8396
rect 15101 8394 15167 8397
rect 13740 8392 15167 8394
rect 13740 8336 15106 8392
rect 15162 8336 15167 8392
rect 13740 8334 15167 8336
rect 13740 8332 13746 8334
rect 15101 8331 15167 8334
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 24945 8122 25011 8125
rect 26200 8122 27000 8152
rect 24945 8120 27000 8122
rect 24945 8064 24950 8120
rect 25006 8064 27000 8120
rect 24945 8062 27000 8064
rect 24945 8059 25011 8062
rect 26200 8032 27000 8062
rect 24761 7714 24827 7717
rect 26200 7714 27000 7744
rect 24761 7712 27000 7714
rect 24761 7656 24766 7712
rect 24822 7656 27000 7712
rect 24761 7654 27000 7656
rect 24761 7651 24827 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 26200 7624 27000 7654
rect 17946 7583 18262 7584
rect 24853 7306 24919 7309
rect 26200 7306 27000 7336
rect 24853 7304 27000 7306
rect 24853 7248 24858 7304
rect 24914 7248 27000 7304
rect 24853 7246 27000 7248
rect 24853 7243 24919 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 17718 6972 17724 7036
rect 17788 7034 17794 7036
rect 22001 7034 22067 7037
rect 17788 7032 22067 7034
rect 17788 6976 22006 7032
rect 22062 6976 22067 7032
rect 17788 6974 22067 6976
rect 17788 6972 17794 6974
rect 22001 6971 22067 6974
rect 24853 6898 24919 6901
rect 26200 6898 27000 6928
rect 24853 6896 27000 6898
rect 24853 6840 24858 6896
rect 24914 6840 27000 6896
rect 24853 6838 27000 6840
rect 24853 6835 24919 6838
rect 26200 6808 27000 6838
rect 7946 6560 8262 6561
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 24669 6490 24735 6493
rect 26200 6490 27000 6520
rect 24669 6488 27000 6490
rect 24669 6432 24674 6488
rect 24730 6432 27000 6488
rect 24669 6430 27000 6432
rect 24669 6427 24735 6430
rect 26200 6400 27000 6430
rect 24853 6082 24919 6085
rect 26200 6082 27000 6112
rect 24853 6080 27000 6082
rect 24853 6024 24858 6080
rect 24914 6024 27000 6080
rect 24853 6022 27000 6024
rect 24853 6019 24919 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 26200 5992 27000 6022
rect 22946 5951 23262 5952
rect 24945 5674 25011 5677
rect 26200 5674 27000 5704
rect 24945 5672 27000 5674
rect 24945 5616 24950 5672
rect 25006 5616 27000 5672
rect 24945 5614 27000 5616
rect 24945 5611 25011 5614
rect 26200 5584 27000 5614
rect 22645 5540 22711 5541
rect 22645 5536 22692 5540
rect 22756 5538 22762 5540
rect 22645 5480 22650 5536
rect 22645 5476 22692 5480
rect 22756 5478 22802 5538
rect 22756 5476 22762 5478
rect 22645 5475 22711 5476
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 24761 5266 24827 5269
rect 26200 5266 27000 5296
rect 24761 5264 27000 5266
rect 24761 5208 24766 5264
rect 24822 5208 27000 5264
rect 24761 5206 27000 5208
rect 24761 5203 24827 5206
rect 26200 5176 27000 5206
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 24945 4858 25011 4861
rect 26200 4858 27000 4888
rect 24945 4856 27000 4858
rect 24945 4800 24950 4856
rect 25006 4800 27000 4856
rect 24945 4798 27000 4800
rect 24945 4795 25011 4798
rect 26200 4768 27000 4798
rect 24945 4450 25011 4453
rect 26200 4450 27000 4480
rect 24945 4448 27000 4450
rect 24945 4392 24950 4448
rect 25006 4392 27000 4448
rect 24945 4390 27000 4392
rect 24945 4387 25011 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 26200 4360 27000 4390
rect 17946 4319 18262 4320
rect 25221 4042 25287 4045
rect 26200 4042 27000 4072
rect 25221 4040 27000 4042
rect 25221 3984 25226 4040
rect 25282 3984 27000 4040
rect 25221 3982 27000 3984
rect 25221 3979 25287 3982
rect 26200 3952 27000 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 24945 3634 25011 3637
rect 26200 3634 27000 3664
rect 24945 3632 27000 3634
rect 24945 3576 24950 3632
rect 25006 3576 27000 3632
rect 24945 3574 27000 3576
rect 24945 3571 25011 3574
rect 26200 3544 27000 3574
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 25129 3226 25195 3229
rect 26200 3226 27000 3256
rect 25129 3224 27000 3226
rect 25129 3168 25134 3224
rect 25190 3168 27000 3224
rect 25129 3166 27000 3168
rect 25129 3163 25195 3166
rect 26200 3136 27000 3166
rect 24853 2818 24919 2821
rect 26200 2818 27000 2848
rect 24853 2816 27000 2818
rect 24853 2760 24858 2816
rect 24914 2760 27000 2816
rect 24853 2758 27000 2760
rect 24853 2755 24919 2758
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 26200 2728 27000 2758
rect 22946 2687 23262 2688
rect 24945 2410 25011 2413
rect 26200 2410 27000 2440
rect 24945 2408 27000 2410
rect 24945 2352 24950 2408
rect 25006 2352 27000 2408
rect 24945 2350 27000 2352
rect 24945 2347 25011 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 22185 2002 22251 2005
rect 26200 2002 27000 2032
rect 22185 2000 27000 2002
rect 22185 1944 22190 2000
rect 22246 1944 27000 2000
rect 22185 1942 27000 1944
rect 22185 1939 22251 1942
rect 26200 1912 27000 1942
rect 22093 1594 22159 1597
rect 26200 1594 27000 1624
rect 22093 1592 27000 1594
rect 22093 1536 22098 1592
rect 22154 1536 27000 1592
rect 22093 1534 27000 1536
rect 22093 1531 22159 1534
rect 26200 1504 27000 1534
rect 22093 1186 22159 1189
rect 26200 1186 27000 1216
rect 22093 1184 27000 1186
rect 22093 1128 22098 1184
rect 22154 1128 27000 1184
rect 22093 1126 27000 1128
rect 22093 1123 22159 1126
rect 26200 1096 27000 1126
rect 25037 778 25103 781
rect 26200 778 27000 808
rect 25037 776 27000 778
rect 25037 720 25042 776
rect 25098 720 27000 776
rect 25037 718 27000 720
rect 25037 715 25103 718
rect 26200 688 27000 718
rect 23381 370 23447 373
rect 26200 370 27000 400
rect 23381 368 27000 370
rect 23381 312 23386 368
rect 23442 312 27000 368
rect 23381 310 27000 312
rect 23381 307 23447 310
rect 26200 280 27000 310
<< via3 >>
rect 4844 26148 4908 26212
rect 19380 25060 19444 25124
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 17540 23428 17604 23492
rect 22140 23428 22204 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 20116 22748 20180 22812
rect 16804 22536 16868 22540
rect 16804 22480 16854 22536
rect 16854 22480 16868 22536
rect 16804 22476 16868 22480
rect 18644 22476 18708 22540
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 9444 21796 9508 21860
rect 24532 21856 24596 21860
rect 24532 21800 24582 21856
rect 24582 21800 24596 21856
rect 24532 21796 24596 21800
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 19748 21660 19812 21724
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 13676 20708 13740 20772
rect 16436 20844 16500 20908
rect 22324 20708 22388 20772
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 15884 20632 15948 20636
rect 15884 20576 15898 20632
rect 15898 20576 15948 20632
rect 15884 20572 15948 20576
rect 20852 20436 20916 20500
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 16436 19892 16500 19956
rect 19564 19892 19628 19956
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 20668 19620 20732 19684
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 15148 19348 15212 19412
rect 16068 19348 16132 19412
rect 16436 19348 16500 19412
rect 21036 19076 21100 19140
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 16620 18804 16684 18868
rect 19012 18804 19076 18868
rect 22692 18804 22756 18868
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 4844 17716 4908 17780
rect 19380 17716 19444 17780
rect 15148 17444 15212 17508
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 16804 17308 16868 17372
rect 22508 17368 22572 17372
rect 22508 17312 22522 17368
rect 22522 17312 22572 17368
rect 22508 17308 22572 17312
rect 16436 17036 16500 17100
rect 23428 17036 23492 17100
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 19380 16824 19444 16828
rect 19380 16768 19430 16824
rect 19430 16768 19444 16824
rect 19380 16764 19444 16768
rect 17724 16628 17788 16692
rect 19564 16492 19628 16556
rect 18460 16356 18524 16420
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 24532 16084 24596 16148
rect 22692 15948 22756 16012
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 22140 15540 22204 15604
rect 22324 15268 22388 15332
rect 22692 15268 22756 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 20668 14860 20732 14924
rect 19748 14724 19812 14788
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 18644 14588 18708 14652
rect 18828 14588 18892 14652
rect 18828 14316 18892 14380
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 20116 13636 20180 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 19380 13500 19444 13564
rect 19012 13288 19076 13292
rect 19012 13232 19062 13288
rect 19062 13232 19076 13288
rect 19012 13228 19076 13232
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18460 12820 18524 12884
rect 23428 12820 23492 12884
rect 20852 12548 20916 12612
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 22508 12276 22572 12340
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 21036 11384 21100 11388
rect 21036 11328 21050 11384
rect 21050 11328 21100 11384
rect 21036 11324 21100 11328
rect 9444 11052 9508 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 16068 10372 16132 10436
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 17540 10236 17604 10300
rect 16620 9964 16684 10028
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 15884 9420 15948 9484
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 13676 8332 13740 8396
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 17724 6972 17788 7036
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 22692 5536 22756 5540
rect 22692 5480 22706 5536
rect 22706 5480 22756 5536
rect 22692 5476 22756 5480
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 4843 26212 4909 26213
rect 4843 26148 4844 26212
rect 4908 26148 4909 26212
rect 4843 26147 4909 26148
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 4846 17781 4906 26147
rect 19379 25124 19445 25125
rect 19379 25060 19380 25124
rect 19444 25060 19445 25124
rect 19379 25059 19445 25060
rect 7944 23968 8264 24528
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 17944 23968 18264 24528
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17539 23492 17605 23493
rect 17539 23428 17540 23492
rect 17604 23428 17605 23492
rect 17539 23427 17605 23428
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 16803 22540 16869 22541
rect 16803 22476 16804 22540
rect 16868 22476 16869 22540
rect 16803 22475 16869 22476
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 9443 21860 9509 21861
rect 9443 21796 9444 21860
rect 9508 21796 9509 21860
rect 9443 21795 9509 21796
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 4843 17780 4909 17781
rect 4843 17716 4844 17780
rect 4908 17716 4909 17780
rect 4843 17715 4909 17716
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 9446 11117 9506 21795
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 16435 20908 16501 20909
rect 16435 20844 16436 20908
rect 16500 20844 16501 20908
rect 16435 20843 16501 20844
rect 13675 20772 13741 20773
rect 13675 20708 13676 20772
rect 13740 20708 13741 20772
rect 13675 20707 13741 20708
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 9443 11116 9509 11117
rect 9443 11052 9444 11116
rect 9508 11052 9509 11116
rect 9443 11051 9509 11052
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 13678 8397 13738 20707
rect 15883 20636 15949 20637
rect 15883 20572 15884 20636
rect 15948 20572 15949 20636
rect 15883 20571 15949 20572
rect 15147 19412 15213 19413
rect 15147 19348 15148 19412
rect 15212 19348 15213 19412
rect 15147 19347 15213 19348
rect 15150 17509 15210 19347
rect 15147 17508 15213 17509
rect 15147 17444 15148 17508
rect 15212 17444 15213 17508
rect 15147 17443 15213 17444
rect 15886 9485 15946 20571
rect 16438 19957 16498 20843
rect 16435 19956 16501 19957
rect 16435 19892 16436 19956
rect 16500 19892 16501 19956
rect 16435 19891 16501 19892
rect 16067 19412 16133 19413
rect 16067 19348 16068 19412
rect 16132 19348 16133 19412
rect 16067 19347 16133 19348
rect 16435 19412 16501 19413
rect 16435 19348 16436 19412
rect 16500 19348 16501 19412
rect 16435 19347 16501 19348
rect 16070 10437 16130 19347
rect 16438 17101 16498 19347
rect 16619 18868 16685 18869
rect 16619 18804 16620 18868
rect 16684 18804 16685 18868
rect 16619 18803 16685 18804
rect 16435 17100 16501 17101
rect 16435 17036 16436 17100
rect 16500 17036 16501 17100
rect 16435 17035 16501 17036
rect 16067 10436 16133 10437
rect 16067 10372 16068 10436
rect 16132 10372 16133 10436
rect 16067 10371 16133 10372
rect 16622 10029 16682 18803
rect 16806 17373 16866 22475
rect 16803 17372 16869 17373
rect 16803 17308 16804 17372
rect 16868 17308 16869 17372
rect 16803 17307 16869 17308
rect 17542 10301 17602 23427
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 18643 22540 18709 22541
rect 18643 22476 18644 22540
rect 18708 22476 18709 22540
rect 18643 22475 18709 22476
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17723 16692 17789 16693
rect 17723 16628 17724 16692
rect 17788 16628 17789 16692
rect 17723 16627 17789 16628
rect 17539 10300 17605 10301
rect 17539 10236 17540 10300
rect 17604 10236 17605 10300
rect 17539 10235 17605 10236
rect 16619 10028 16685 10029
rect 16619 9964 16620 10028
rect 16684 9964 16685 10028
rect 16619 9963 16685 9964
rect 15883 9484 15949 9485
rect 15883 9420 15884 9484
rect 15948 9420 15949 9484
rect 15883 9419 15949 9420
rect 13675 8396 13741 8397
rect 13675 8332 13676 8396
rect 13740 8332 13741 8396
rect 13675 8331 13741 8332
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 17726 7037 17786 16627
rect 17944 16352 18264 17376
rect 18459 16420 18525 16421
rect 18459 16356 18460 16420
rect 18524 16356 18525 16420
rect 18459 16355 18525 16356
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 18462 12885 18522 16355
rect 18646 14653 18706 22475
rect 19011 18868 19077 18869
rect 19011 18804 19012 18868
rect 19076 18804 19077 18868
rect 19011 18803 19077 18804
rect 18643 14652 18709 14653
rect 18643 14588 18644 14652
rect 18708 14588 18709 14652
rect 18643 14587 18709 14588
rect 18827 14652 18893 14653
rect 18827 14588 18828 14652
rect 18892 14588 18893 14652
rect 18827 14587 18893 14588
rect 18830 14381 18890 14587
rect 18827 14380 18893 14381
rect 18827 14316 18828 14380
rect 18892 14316 18893 14380
rect 18827 14315 18893 14316
rect 19014 13293 19074 18803
rect 19382 17781 19442 25059
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22139 23492 22205 23493
rect 22139 23428 22140 23492
rect 22204 23428 22205 23492
rect 22139 23427 22205 23428
rect 20115 22812 20181 22813
rect 20115 22748 20116 22812
rect 20180 22748 20181 22812
rect 20115 22747 20181 22748
rect 19747 21724 19813 21725
rect 19747 21660 19748 21724
rect 19812 21660 19813 21724
rect 19747 21659 19813 21660
rect 19563 19956 19629 19957
rect 19563 19892 19564 19956
rect 19628 19892 19629 19956
rect 19563 19891 19629 19892
rect 19379 17780 19445 17781
rect 19379 17716 19380 17780
rect 19444 17716 19445 17780
rect 19379 17715 19445 17716
rect 19379 16828 19445 16829
rect 19379 16764 19380 16828
rect 19444 16764 19445 16828
rect 19379 16763 19445 16764
rect 19382 13565 19442 16763
rect 19566 16557 19626 19891
rect 19563 16556 19629 16557
rect 19563 16492 19564 16556
rect 19628 16492 19629 16556
rect 19563 16491 19629 16492
rect 19750 14789 19810 21659
rect 19747 14788 19813 14789
rect 19747 14724 19748 14788
rect 19812 14724 19813 14788
rect 19747 14723 19813 14724
rect 20118 13701 20178 22747
rect 20851 20500 20917 20501
rect 20851 20436 20852 20500
rect 20916 20436 20917 20500
rect 20851 20435 20917 20436
rect 20667 19684 20733 19685
rect 20667 19620 20668 19684
rect 20732 19620 20733 19684
rect 20667 19619 20733 19620
rect 20670 14925 20730 19619
rect 20667 14924 20733 14925
rect 20667 14860 20668 14924
rect 20732 14860 20733 14924
rect 20667 14859 20733 14860
rect 20115 13700 20181 13701
rect 20115 13636 20116 13700
rect 20180 13636 20181 13700
rect 20115 13635 20181 13636
rect 19379 13564 19445 13565
rect 19379 13500 19380 13564
rect 19444 13500 19445 13564
rect 19379 13499 19445 13500
rect 19011 13292 19077 13293
rect 19011 13228 19012 13292
rect 19076 13228 19077 13292
rect 19011 13227 19077 13228
rect 18459 12884 18525 12885
rect 18459 12820 18460 12884
rect 18524 12820 18525 12884
rect 18459 12819 18525 12820
rect 20854 12613 20914 20435
rect 21035 19140 21101 19141
rect 21035 19076 21036 19140
rect 21100 19076 21101 19140
rect 21035 19075 21101 19076
rect 20851 12612 20917 12613
rect 20851 12548 20852 12612
rect 20916 12548 20917 12612
rect 20851 12547 20917 12548
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 21038 11389 21098 19075
rect 22142 15605 22202 23427
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 24531 21860 24597 21861
rect 24531 21796 24532 21860
rect 24596 21796 24597 21860
rect 24531 21795 24597 21796
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22323 20772 22389 20773
rect 22323 20708 22324 20772
rect 22388 20708 22389 20772
rect 22323 20707 22389 20708
rect 22139 15604 22205 15605
rect 22139 15540 22140 15604
rect 22204 15540 22205 15604
rect 22139 15539 22205 15540
rect 22326 15333 22386 20707
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22691 18868 22757 18869
rect 22691 18804 22692 18868
rect 22756 18804 22757 18868
rect 22691 18803 22757 18804
rect 22507 17372 22573 17373
rect 22507 17308 22508 17372
rect 22572 17308 22573 17372
rect 22507 17307 22573 17308
rect 22323 15332 22389 15333
rect 22323 15268 22324 15332
rect 22388 15268 22389 15332
rect 22323 15267 22389 15268
rect 22510 12341 22570 17307
rect 22694 16013 22754 18803
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 23427 17100 23493 17101
rect 23427 17036 23428 17100
rect 23492 17036 23493 17100
rect 23427 17035 23493 17036
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22691 16012 22757 16013
rect 22691 15948 22692 16012
rect 22756 15948 22757 16012
rect 22691 15947 22757 15948
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22691 15332 22757 15333
rect 22691 15268 22692 15332
rect 22756 15268 22757 15332
rect 22691 15267 22757 15268
rect 22507 12340 22573 12341
rect 22507 12276 22508 12340
rect 22572 12276 22573 12340
rect 22507 12275 22573 12276
rect 21035 11388 21101 11389
rect 21035 11324 21036 11388
rect 21100 11324 21101 11388
rect 21035 11323 21101 11324
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17723 7036 17789 7037
rect 17723 6972 17724 7036
rect 17788 6972 17789 7036
rect 17723 6971 17789 6972
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 22694 5541 22754 15267
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 23430 12885 23490 17035
rect 24534 16149 24594 21795
rect 24531 16148 24597 16149
rect 24531 16084 24532 16148
rect 24596 16084 24597 16148
rect 24531 16083 24597 16084
rect 23427 12884 23493 12885
rect 23427 12820 23428 12884
rect 23492 12820 23493 12884
rect 23427 12819 23493 12820
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22691 5540 22757 5541
rect 22691 5476 22692 5540
rect 22756 5476 22757 5540
rect 22691 5475 22757 5476
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _072_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 18584 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _073_
timestamp 1676037725
transform 1 0 19872 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _074_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _075_
timestamp 1676037725
transform 1 0 25024 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _076_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1676037725
transform 1 0 24656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1676037725
transform 1 0 24656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _079_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _080_
timestamp 1676037725
transform 1 0 24564 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _081_
timestamp 1676037725
transform 1 0 22632 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _082_
timestamp 1676037725
transform 1 0 21988 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _083_
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1676037725
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _085_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _086_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19412 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1676037725
transform 1 0 21344 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _088_
timestamp 1676037725
transform 1 0 24748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _089_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _090_
timestamp 1676037725
transform 1 0 24656 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _091_
timestamp 1676037725
transform 1 0 24564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1676037725
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1676037725
transform 1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _094_
timestamp 1676037725
transform 1 0 18032 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _096_
timestamp 1676037725
transform 1 0 15180 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1676037725
transform 1 0 18032 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1676037725
transform 1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _100_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1676037725
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1676037725
transform 1 0 5152 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 6532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1676037725
transform 1 0 4508 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 13432 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 15824 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 15732 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 13432 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1676037725
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1676037725
transform 1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1676037725
transform 1 0 7728 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 7820 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 12880 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 18400 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 14812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1676037725
transform 1 0 3220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1676037725
transform 1 0 5796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1676037725
transform 1 0 2208 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _125_
timestamp 1676037725
transform 1 0 4508 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _126_
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _127_
timestamp 1676037725
transform 1 0 5152 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _128_
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1676037725
transform 1 0 9200 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _130_
timestamp 1676037725
transform 1 0 5152 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _131_
timestamp 1676037725
transform 1 0 4508 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 24380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 4968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 2024 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 22632 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 3680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 24472 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 23092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 19688 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 8280 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1676037725
transform 1 0 25300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1676037725
transform 1 0 23000 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1676037725
transform 1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1676037725
transform 1 0 21160 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 13708 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 8096 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 7176 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 20608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 17664 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 20424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 11040 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 10304 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 9384 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 22264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 17020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 25300 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 22724 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 2668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 6256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 5152 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 16560 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 14444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 6624 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 6716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 2852 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 4140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 6440 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 4784 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 9568 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 20792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 6808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 7176 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 2392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 17296 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 24012 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 25300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 2116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform 1 0 2116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 2392 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 2116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23000 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20240 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23092 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22908 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20700 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22172 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22816 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25116 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21988 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20240 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21620 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17480 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16100 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13064 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12696 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 9936 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16284 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18860 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16284 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17112 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_prog_clk
timestamp 1676037725
transform 1 0 9568 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_prog_clk
timestamp 1676037725
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_prog_clk
timestamp 1676037725
transform 1 0 10396 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_prog_clk
timestamp 1676037725
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_prog_clk
timestamp 1676037725
transform 1 0 18216 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_prog_clk
timestamp 1676037725
transform 1 0 20792 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_prog_clk
timestamp 1676037725
transform 1 0 18216 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 18496
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1676037725
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1676037725
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1676037725
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1676037725
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1676037725
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1676037725
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_265
timestamp 1676037725
transform 1 0 25484 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 1676037725
transform 1 0 18124 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_202
timestamp 1676037725
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_244
timestamp 1676037725
transform 1 0 23552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_264
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1676037725
transform 1 0 20700 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1676037725
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_258
timestamp 1676037725
transform 1 0 24840 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1676037725
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_244
timestamp 1676037725
transform 1 0 23552 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_264
timestamp 1676037725
transform 1 0 25392 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_229
timestamp 1676037725
transform 1 0 22172 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_232
timestamp 1676037725
transform 1 0 22448 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_250
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_259
timestamp 1676037725
transform 1 0 24932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_244
timestamp 1676037725
transform 1 0 23552 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_264
timestamp 1676037725
transform 1 0 25392 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_217
timestamp 1676037725
transform 1 0 21068 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_223
timestamp 1676037725
transform 1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1676037725
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_244
timestamp 1676037725
transform 1 0 23552 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_217
timestamp 1676037725
transform 1 0 21068 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_223
timestamp 1676037725
transform 1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_259
timestamp 1676037725
transform 1 0 24932 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_211
timestamp 1676037725
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1676037725
transform 1 0 20884 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_216
timestamp 1676037725
transform 1 0 20976 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1676037725
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_230
timestamp 1676037725
transform 1 0 22264 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_250
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_209
timestamp 1676037725
transform 1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_216
timestamp 1676037725
transform 1 0 20976 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_220
timestamp 1676037725
transform 1 0 21344 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_117
timestamp 1676037725
transform 1 0 11868 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_193
timestamp 1676037725
transform 1 0 18860 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_217
timestamp 1676037725
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_222
timestamp 1676037725
transform 1 0 21528 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_229
timestamp 1676037725
transform 1 0 22172 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_259
timestamp 1676037725
transform 1 0 24932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_187
timestamp 1676037725
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_194
timestamp 1676037725
transform 1 0 18952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_201
timestamp 1676037725
transform 1 0 19596 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1676037725
transform 1 0 20240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_212
timestamp 1676037725
transform 1 0 20608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1676037725
transform 1 0 20976 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_244
timestamp 1676037725
transform 1 0 23552 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_264
timestamp 1676037725
transform 1 0 25392 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_182
timestamp 1676037725
transform 1 0 17848 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_202
timestamp 1676037725
transform 1 0 19688 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_216
timestamp 1676037725
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_241
timestamp 1676037725
transform 1 0 23276 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1676037725
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_264
timestamp 1676037725
transform 1 0 25392 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_165
timestamp 1676037725
transform 1 0 16284 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1676037725
transform 1 0 17204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_180
timestamp 1676037725
transform 1 0 17664 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_187
timestamp 1676037725
transform 1 0 18308 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_194
timestamp 1676037725
transform 1 0 18952 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_201
timestamp 1676037725
transform 1 0 19596 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_208
timestamp 1676037725
transform 1 0 20240 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_215
timestamp 1676037725
transform 1 0 20884 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_244
timestamp 1676037725
transform 1 0 23552 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1676037725
transform 1 0 25392 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_149
timestamp 1676037725
transform 1 0 14812 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_155
timestamp 1676037725
transform 1 0 15364 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_159
timestamp 1676037725
transform 1 0 15732 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1676037725
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_173
timestamp 1676037725
transform 1 0 17020 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_180
timestamp 1676037725
transform 1 0 17664 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1676037725
transform 1 0 18308 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_201
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_208
timestamp 1676037725
transform 1 0 20240 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_216
timestamp 1676037725
transform 1 0 20976 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_225
timestamp 1676037725
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_230
timestamp 1676037725
transform 1 0 22264 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_258
timestamp 1676037725
transform 1 0 24840 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1676037725
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_151
timestamp 1676037725
transform 1 0 14996 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1676037725
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1676037725
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_171
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_194
timestamp 1676037725
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_198
timestamp 1676037725
transform 1 0 19320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_219
timestamp 1676037725
transform 1 0 21252 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1676037725
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1676037725
transform 1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1676037725
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1676037725
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1676037725
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1676037725
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_262
timestamp 1676037725
transform 1 0 25208 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_265
timestamp 1676037725
transform 1 0 25484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_121
timestamp 1676037725
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_126
timestamp 1676037725
transform 1 0 12696 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_163
timestamp 1676037725
transform 1 0 16100 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 1676037725
transform 1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_204
timestamp 1676037725
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_247
timestamp 1676037725
transform 1 0 23828 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_254
timestamp 1676037725
transform 1 0 24472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_261
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_265
timestamp 1676037725
transform 1 0 25484 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1676037725
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1676037725
transform 1 0 11408 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_163
timestamp 1676037725
transform 1 0 16100 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_187
timestamp 1676037725
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1676037725
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_199
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_222
timestamp 1676037725
transform 1 0 21528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_246
timestamp 1676037725
transform 1 0 23736 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_264
timestamp 1676037725
transform 1 0 25392 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_119
timestamp 1676037725
transform 1 0 12052 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_126
timestamp 1676037725
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_133
timestamp 1676037725
transform 1 0 13340 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1676037725
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1676037725
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_182
timestamp 1676037725
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1676037725
transform 1 0 20056 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_210
timestamp 1676037725
transform 1 0 20424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_231
timestamp 1676037725
transform 1 0 22356 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_235
timestamp 1676037725
transform 1 0 22724 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_264
timestamp 1676037725
transform 1 0 25392 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1676037725
transform 1 0 10488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_124
timestamp 1676037725
transform 1 0 12512 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1676037725
transform 1 0 13156 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1676037725
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_187
timestamp 1676037725
transform 1 0 18308 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1676037725
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_208
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1676037725
transform 1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp 1676037725
transform 1 0 22632 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_238
timestamp 1676037725
transform 1 0 23000 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_259
timestamp 1676037725
transform 1 0 24932 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1676037725
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_98
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_103
timestamp 1676037725
transform 1 0 10580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_135
timestamp 1676037725
transform 1 0 13524 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_142
timestamp 1676037725
transform 1 0 14168 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_147
timestamp 1676037725
transform 1 0 14628 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_152
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1676037725
transform 1 0 15732 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_191
timestamp 1676037725
transform 1 0 18676 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1676037725
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1676037725
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1676037725
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_231
timestamp 1676037725
transform 1 0 22356 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_235
timestamp 1676037725
transform 1 0 22724 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_256
timestamp 1676037725
transform 1 0 24656 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_263
timestamp 1676037725
transform 1 0 25300 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_81
timestamp 1676037725
transform 1 0 8556 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_91
timestamp 1676037725
transform 1 0 9476 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_98
timestamp 1676037725
transform 1 0 10120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1676037725
transform 1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_135
timestamp 1676037725
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_163
timestamp 1676037725
transform 1 0 16100 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_167
timestamp 1676037725
transform 1 0 16468 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 1676037725
transform 1 0 16744 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1676037725
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1676037725
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_230
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_238
timestamp 1676037725
transform 1 0 23000 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_258
timestamp 1676037725
transform 1 0 24840 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_75
timestamp 1676037725
transform 1 0 8004 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_90
timestamp 1676037725
transform 1 0 9384 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1676037725
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1676037725
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_135
timestamp 1676037725
transform 1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1676037725
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1676037725
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1676037725
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_171
timestamp 1676037725
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1676037725
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1676037725
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_220
timestamp 1676037725
transform 1 0 21344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1676037725
transform 1 0 22816 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1676037725
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_251
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_259
timestamp 1676037725
transform 1 0 24932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_265
timestamp 1676037725
transform 1 0 25484 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_37
timestamp 1676037725
transform 1 0 4508 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_42
timestamp 1676037725
transform 1 0 4968 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_46
timestamp 1676037725
transform 1 0 5336 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_58
timestamp 1676037725
transform 1 0 6440 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1676037725
transform 1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1676037725
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_75
timestamp 1676037725
transform 1 0 8004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_89
timestamp 1676037725
transform 1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_94
timestamp 1676037725
transform 1 0 9752 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_101
timestamp 1676037725
transform 1 0 10396 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_114
timestamp 1676037725
transform 1 0 11592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1676037725
transform 1 0 16100 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1676037725
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1676037725
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_259
timestamp 1676037725
transform 1 0 24932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_33
timestamp 1676037725
transform 1 0 4140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1676037725
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1676037725
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_76
timestamp 1676037725
transform 1 0 8096 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_80
timestamp 1676037725
transform 1 0 8464 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_108
timestamp 1676037725
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_135
timestamp 1676037725
transform 1 0 13524 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1676037725
transform 1 0 14168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_146
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1676037725
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1676037725
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_180
timestamp 1676037725
transform 1 0 17664 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_184
timestamp 1676037725
transform 1 0 18032 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_207
timestamp 1676037725
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_221
timestamp 1676037725
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_231
timestamp 1676037725
transform 1 0 22356 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1676037725
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_261
timestamp 1676037725
transform 1 0 25116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_265
timestamp 1676037725
transform 1 0 25484 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1676037725
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_35
timestamp 1676037725
transform 1 0 4324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1676037725
transform 1 0 4784 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_54
timestamp 1676037725
transform 1 0 6072 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_61
timestamp 1676037725
transform 1 0 6716 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_68
timestamp 1676037725
transform 1 0 7360 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_75
timestamp 1676037725
transform 1 0 8004 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1676037725
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1676037725
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1676037725
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1676037725
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1676037725
transform 1 0 16744 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1676037725
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_187
timestamp 1676037725
transform 1 0 18308 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1676037725
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_212
timestamp 1676037725
transform 1 0 20608 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_233
timestamp 1676037725
transform 1 0 22540 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_239
timestamp 1676037725
transform 1 0 23092 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_260
timestamp 1676037725
transform 1 0 25024 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_8
timestamp 1676037725
transform 1 0 1840 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_26
timestamp 1676037725
transform 1 0 3496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_40
timestamp 1676037725
transform 1 0 4784 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_47
timestamp 1676037725
transform 1 0 5428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1676037725
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1676037725
transform 1 0 6808 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_67
timestamp 1676037725
transform 1 0 7268 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_74
timestamp 1676037725
transform 1 0 7912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_162
timestamp 1676037725
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1676037725
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1676037725
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1676037725
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_219
timestamp 1676037725
transform 1 0 21252 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_247
timestamp 1676037725
transform 1 0 23828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1676037725
transform 1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_12
timestamp 1676037725
transform 1 0 2208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_19
timestamp 1676037725
transform 1 0 2852 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1676037725
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_31
timestamp 1676037725
transform 1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_35
timestamp 1676037725
transform 1 0 4324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp 1676037725
transform 1 0 4784 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_47
timestamp 1676037725
transform 1 0 5428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_54
timestamp 1676037725
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_61
timestamp 1676037725
transform 1 0 6716 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_75
timestamp 1676037725
transform 1 0 8004 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1676037725
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_152
timestamp 1676037725
transform 1 0 15088 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1676037725
transform 1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1676037725
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_202
timestamp 1676037725
transform 1 0 19688 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_208
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_229
timestamp 1676037725
transform 1 0 22172 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_242
timestamp 1676037725
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1676037725
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_23
timestamp 1676037725
transform 1 0 3220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_29
timestamp 1676037725
transform 1 0 3772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_33
timestamp 1676037725
transform 1 0 4140 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_47
timestamp 1676037725
transform 1 0 5428 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1676037725
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1676037725
transform 1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1676037725
transform 1 0 7360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1676037725
transform 1 0 8004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_82
timestamp 1676037725
transform 1 0 8648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 1676037725
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_117
timestamp 1676037725
transform 1 0 11868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1676037725
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_159
timestamp 1676037725
transform 1 0 15732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1676037725
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_219
timestamp 1676037725
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_236
timestamp 1676037725
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_240
timestamp 1676037725
transform 1 0 23184 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_261
timestamp 1676037725
transform 1 0 25116 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_265
timestamp 1676037725
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1676037725
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_40
timestamp 1676037725
transform 1 0 4784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_54
timestamp 1676037725
transform 1 0 6072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_61
timestamp 1676037725
transform 1 0 6716 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_75
timestamp 1676037725
transform 1 0 8004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1676037725
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1676037725
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_110
timestamp 1676037725
transform 1 0 11224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_134
timestamp 1676037725
transform 1 0 13432 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1676037725
transform 1 0 15732 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_167
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_174
timestamp 1676037725
transform 1 0 17112 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_178
timestamp 1676037725
transform 1 0 17480 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_208
timestamp 1676037725
transform 1 0 20240 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_212
timestamp 1676037725
transform 1 0 20608 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1676037725
transform 1 0 20884 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_237
timestamp 1676037725
transform 1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_264
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_8
timestamp 1676037725
transform 1 0 1840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_35
timestamp 1676037725
transform 1 0 4324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_47
timestamp 1676037725
transform 1 0 5428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1676037725
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_68
timestamp 1676037725
transform 1 0 7360 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_75
timestamp 1676037725
transform 1 0 8004 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_82
timestamp 1676037725
transform 1 0 8648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_106
timestamp 1676037725
transform 1 0 10856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_128
timestamp 1676037725
transform 1 0 12880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_132
timestamp 1676037725
transform 1 0 13248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_155
timestamp 1676037725
transform 1 0 15364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_163
timestamp 1676037725
transform 1 0 16100 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1676037725
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1676037725
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_217
timestamp 1676037725
transform 1 0 21068 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_241
timestamp 1676037725
transform 1 0 23276 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_263
timestamp 1676037725
transform 1 0 25300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_9
timestamp 1676037725
transform 1 0 1932 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 1676037725
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_47
timestamp 1676037725
transform 1 0 5428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_54
timestamp 1676037725
transform 1 0 6072 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_58
timestamp 1676037725
transform 1 0 6440 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_62
timestamp 1676037725
transform 1 0 6808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_79
timestamp 1676037725
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_92
timestamp 1676037725
transform 1 0 9568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1676037725
transform 1 0 10764 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1676037725
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1676037725
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_147
timestamp 1676037725
transform 1 0 14628 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_155
timestamp 1676037725
transform 1 0 15364 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_178
timestamp 1676037725
transform 1 0 17480 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_191
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_219
timestamp 1676037725
transform 1 0 21252 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_232
timestamp 1676037725
transform 1 0 22448 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_245
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1676037725
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_9
timestamp 1676037725
transform 1 0 1932 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_13
timestamp 1676037725
transform 1 0 2300 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_17
timestamp 1676037725
transform 1 0 2668 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_34
timestamp 1676037725
transform 1 0 4232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1676037725
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1676037725
transform 1 0 6808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_82
timestamp 1676037725
transform 1 0 8648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_106
timestamp 1676037725
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_130
timestamp 1676037725
transform 1 0 13064 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_147
timestamp 1676037725
transform 1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_160
timestamp 1676037725
transform 1 0 15824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_182
timestamp 1676037725
transform 1 0 17848 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1676037725
transform 1 0 20056 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_219
timestamp 1676037725
transform 1 0 21252 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_262
timestamp 1676037725
transform 1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_9
timestamp 1676037725
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_26
timestamp 1676037725
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_45
timestamp 1676037725
transform 1 0 5244 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_62
timestamp 1676037725
transform 1 0 6808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1676037725
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_87
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_92
timestamp 1676037725
transform 1 0 9568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_96
timestamp 1676037725
transform 1 0 9936 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_100
timestamp 1676037725
transform 1 0 10304 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_124
timestamp 1676037725
transform 1 0 12512 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_128
timestamp 1676037725
transform 1 0 12880 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1676037725
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_163
timestamp 1676037725
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_176
timestamp 1676037725
transform 1 0 17296 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_189
timestamp 1676037725
transform 1 0 18492 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_203
timestamp 1676037725
transform 1 0 19780 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1676037725
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1676037725
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_9
timestamp 1676037725
transform 1 0 1932 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_13
timestamp 1676037725
transform 1 0 2300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_16
timestamp 1676037725
transform 1 0 2576 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_34
timestamp 1676037725
transform 1 0 4232 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1676037725
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_63
timestamp 1676037725
transform 1 0 6900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_68
timestamp 1676037725
transform 1 0 7360 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_86
timestamp 1676037725
transform 1 0 9016 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1676037725
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_124
timestamp 1676037725
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_132
timestamp 1676037725
transform 1 0 13248 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1676037725
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_164
timestamp 1676037725
transform 1 0 16192 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_204
timestamp 1676037725
transform 1 0 19872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_217
timestamp 1676037725
transform 1 0 21068 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_221
timestamp 1676037725
transform 1 0 21436 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_261
timestamp 1676037725
transform 1 0 25116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_265
timestamp 1676037725
transform 1 0 25484 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_9
timestamp 1676037725
transform 1 0 1932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1676037725
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_35
timestamp 1676037725
transform 1 0 4324 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_42
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1676037725
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_91
timestamp 1676037725
transform 1 0 9476 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_111
timestamp 1676037725
transform 1 0 11316 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_131
timestamp 1676037725
transform 1 0 13156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_147
timestamp 1676037725
transform 1 0 14628 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_171
timestamp 1676037725
transform 1 0 16836 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_184
timestamp 1676037725
transform 1 0 18032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1676037725
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_219
timestamp 1676037725
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_243
timestamp 1676037725
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_9
timestamp 1676037725
transform 1 0 1932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_13
timestamp 1676037725
transform 1 0 2300 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_16
timestamp 1676037725
transform 1 0 2576 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1676037725
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1676037725
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_73
timestamp 1676037725
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1676037725
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_115
timestamp 1676037725
transform 1 0 11684 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_135
timestamp 1676037725
transform 1 0 13524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_150
timestamp 1676037725
transform 1 0 14904 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_158
timestamp 1676037725
transform 1 0 15640 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_163
timestamp 1676037725
transform 1 0 16100 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1676037725
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_204
timestamp 1676037725
transform 1 0 19872 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_210
timestamp 1676037725
transform 1 0 20424 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_227
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_250
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_258
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_264
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_9
timestamp 1676037725
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1676037725
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1676037725
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1676037725
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1676037725
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1676037725
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1676037725
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1676037725
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_113
timestamp 1676037725
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1676037725
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_169
timestamp 1676037725
transform 1 0 16652 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1676037725
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1676037725
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_227
timestamp 1676037725
transform 1 0 21988 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 6808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 20056 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 8372 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 12880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 2576 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 13064 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 7176 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1676037725
transform 1 0 18676 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1676037725
transform 1 0 18032 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 15456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 12420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1676037725
transform 1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1676037725
transform 1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 20700 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 18676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 24196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1676037725
transform 1 0 3956 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 4692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 16468 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 7084 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 6440 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1676037725
transform 1 0 7636 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1676037725
transform 1 0 6992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1676037725
transform 1 0 3220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 4508 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 5152 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 9752 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 9108 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1676037725
transform 1 0 9844 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 16100 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 9292 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1676037725
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1676037725
transform 1 0 6532 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1676037725
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 16836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 7728 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input62 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1676037725
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1676037725
transform 1 0 20608 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1676037725
transform 1 0 23184 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1676037725
transform 1 0 21988 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 1564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1676037725
transform 1 0 3956 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1676037725
transform 1 0 20056 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1676037725
transform 1 0 20056 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1676037725
transform 1 0 22080 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1676037725
transform 1 0 23920 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1676037725
transform 1 0 22632 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1676037725
transform 1 0 22080 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1676037725
transform 1 0 23920 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1676037725
transform 1 0 23920 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1676037725
transform 1 0 22632 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 20792 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 22080 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 22080 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 23920 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 23920 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 20056 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 18216 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 22080 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 22632 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 22080 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 23920 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 22632 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 1748 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 5336 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 6900 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 7176 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 7176 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 2024 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 7544 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 9844 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 11684 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 12052 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 2024 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 2852 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 2024 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 2760 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 2760 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 2024 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 4600 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14904 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19228 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21620 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23276 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23276 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22540 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20700 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22816 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21896 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19320 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18308 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16928 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16468 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15732 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__0_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21344 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15456 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16928 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18032 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14996 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13616 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13524 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12696 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11592 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10672 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9016 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9016 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9016 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8924 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9200 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9752 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10488 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10672 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11776 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12788 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17020 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20424 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_0.mux_l1_in_1__159 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23736 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_2.mux_l2_in_0__165
timestamp 1676037725
transform 1 0 2208 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 4508 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_4.mux_l2_in_0__134
timestamp 1676037725
transform 1 0 3864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_6.mux_l1_in_1__139
timestamp 1676037725
transform 1 0 17388 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_8.mux_l2_in_0__140
timestamp 1676037725
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_10.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 16100 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21620 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_12.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 23828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23368 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_14.mux_l2_in_0__162
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_16.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19320 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_18.mux_l2_in_0__164
timestamp 1676037725
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_28.mux_l2_in_0__166
timestamp 1676037725
transform 1 0 25024 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_30.mux_l2_in_0__167
timestamp 1676037725
transform 1 0 23368 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_32.mux_l2_in_0__132
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_34.mux_l2_in_0__133
timestamp 1676037725
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17020 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_44.mux_l2_in_0__135
timestamp 1676037725
transform 1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20700 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_46.mux_l2_in_0__136
timestamp 1676037725
transform 1 0 18032 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20700 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_48.mux_l2_in_0__137
timestamp 1676037725
transform 1 0 21620 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20516 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_right_track_50.mux_l2_in_0__138
timestamp 1676037725
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19412 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_0.mux_l1_in_1__141
timestamp 1676037725
transform 1 0 20516 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17848 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_2.mux_l2_in_0__147
timestamp 1676037725
transform 1 0 19412 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20240 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_4.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_6.mux_l1_in_1__157
timestamp 1676037725
transform 1 0 5152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17204 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_8.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17664 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13800 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_10.mux_l2_in_0__142
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16652 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_12.mux_l2_in_0__143
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12236 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16468 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_14.mux_l2_in_0__144
timestamp 1676037725
transform 1 0 4692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9936 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_16.mux_l2_in_0__145
timestamp 1676037725
transform 1 0 7728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8280 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_18.mux_l2_in_0__146
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_28.mux_l2_in_0__148
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9200 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17664 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12052 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_30.mux_l2_in_0__149
timestamp 1676037725
transform 1 0 9292 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6532 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_32.mux_l2_in_0__150
timestamp 1676037725
transform 1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_34.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 9752 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10764 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 5796 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_44.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 10120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_46.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 13892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19320 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13892 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_48.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17112 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__0_.mux_top_track_50.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 6440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 26200 280 27000 400 0 FreeSans 480 0 0 0 ccff_tail
port 3 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 4 nsew signal input
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 5 nsew signal input
flabel metal3 s 26200 17416 27000 17536 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 6 nsew signal input
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 7 nsew signal input
flabel metal3 s 26200 18232 27000 18352 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 8 nsew signal input
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 9 nsew signal input
flabel metal3 s 26200 19048 27000 19168 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 10 nsew signal input
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 11 nsew signal input
flabel metal3 s 26200 19864 27000 19984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 12 nsew signal input
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 13 nsew signal input
flabel metal3 s 26200 20680 27000 20800 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 14 nsew signal input
flabel metal3 s 26200 13336 27000 13456 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 15 nsew signal input
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 16 nsew signal input
flabel metal3 s 26200 21496 27000 21616 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 17 nsew signal input
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 18 nsew signal input
flabel metal3 s 26200 22312 27000 22432 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 19 nsew signal input
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 20 nsew signal input
flabel metal3 s 26200 23128 27000 23248 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 21 nsew signal input
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 22 nsew signal input
flabel metal3 s 26200 23944 27000 24064 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 23 nsew signal input
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 24 nsew signal input
flabel metal3 s 26200 24760 27000 24880 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 25 nsew signal input
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 26 nsew signal input
flabel metal3 s 26200 14152 27000 14272 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 27 nsew signal input
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 28 nsew signal input
flabel metal3 s 26200 14968 27000 15088 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 29 nsew signal input
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 30 nsew signal input
flabel metal3 s 26200 15784 27000 15904 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 31 nsew signal input
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 32 nsew signal input
flabel metal3 s 26200 16600 27000 16720 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 33 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 34 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 35 nsew signal tristate
flabel metal3 s 26200 5176 27000 5296 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 36 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 37 nsew signal tristate
flabel metal3 s 26200 5992 27000 6112 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 38 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 39 nsew signal tristate
flabel metal3 s 26200 6808 27000 6928 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 40 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 41 nsew signal tristate
flabel metal3 s 26200 7624 27000 7744 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 42 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 43 nsew signal tristate
flabel metal3 s 26200 8440 27000 8560 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 44 nsew signal tristate
flabel metal3 s 26200 1096 27000 1216 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 45 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 46 nsew signal tristate
flabel metal3 s 26200 9256 27000 9376 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 47 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 48 nsew signal tristate
flabel metal3 s 26200 10072 27000 10192 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 49 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 50 nsew signal tristate
flabel metal3 s 26200 10888 27000 11008 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 51 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 52 nsew signal tristate
flabel metal3 s 26200 11704 27000 11824 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 53 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 54 nsew signal tristate
flabel metal3 s 26200 12520 27000 12640 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 55 nsew signal tristate
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 56 nsew signal tristate
flabel metal3 s 26200 1912 27000 2032 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 57 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 58 nsew signal tristate
flabel metal3 s 26200 2728 27000 2848 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 59 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 60 nsew signal tristate
flabel metal3 s 26200 3544 27000 3664 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 61 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 62 nsew signal tristate
flabel metal3 s 26200 4360 27000 4480 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 63 nsew signal tristate
flabel metal2 s 12714 26200 12770 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 64 nsew signal input
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 65 nsew signal input
flabel metal2 s 16762 26200 16818 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 66 nsew signal input
flabel metal2 s 17130 26200 17186 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 67 nsew signal input
flabel metal2 s 17498 26200 17554 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 68 nsew signal input
flabel metal2 s 17866 26200 17922 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 69 nsew signal input
flabel metal2 s 18234 26200 18290 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 70 nsew signal input
flabel metal2 s 18602 26200 18658 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 71 nsew signal input
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 72 nsew signal input
flabel metal2 s 19338 26200 19394 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 73 nsew signal input
flabel metal2 s 19706 26200 19762 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 74 nsew signal input
flabel metal2 s 13082 26200 13138 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 75 nsew signal input
flabel metal2 s 20074 26200 20130 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 76 nsew signal input
flabel metal2 s 20442 26200 20498 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 77 nsew signal input
flabel metal2 s 20810 26200 20866 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 78 nsew signal input
flabel metal2 s 21178 26200 21234 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 79 nsew signal input
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 80 nsew signal input
flabel metal2 s 21914 26200 21970 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 81 nsew signal input
flabel metal2 s 22282 26200 22338 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 82 nsew signal input
flabel metal2 s 22650 26200 22706 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 83 nsew signal input
flabel metal2 s 23018 26200 23074 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 84 nsew signal input
flabel metal2 s 23386 26200 23442 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 85 nsew signal input
flabel metal2 s 13450 26200 13506 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 86 nsew signal input
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 87 nsew signal input
flabel metal2 s 14186 26200 14242 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 88 nsew signal input
flabel metal2 s 14554 26200 14610 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 89 nsew signal input
flabel metal2 s 14922 26200 14978 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 90 nsew signal input
flabel metal2 s 15290 26200 15346 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 91 nsew signal input
flabel metal2 s 15658 26200 15714 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 92 nsew signal input
flabel metal2 s 16026 26200 16082 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 93 nsew signal input
flabel metal2 s 1674 26200 1730 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 94 nsew signal tristate
flabel metal2 s 5354 26200 5410 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 95 nsew signal tristate
flabel metal2 s 5722 26200 5778 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 96 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 97 nsew signal tristate
flabel metal2 s 6458 26200 6514 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 98 nsew signal tristate
flabel metal2 s 6826 26200 6882 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 99 nsew signal tristate
flabel metal2 s 7194 26200 7250 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 100 nsew signal tristate
flabel metal2 s 7562 26200 7618 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 101 nsew signal tristate
flabel metal2 s 7930 26200 7986 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 102 nsew signal tristate
flabel metal2 s 8298 26200 8354 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 103 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 104 nsew signal tristate
flabel metal2 s 2042 26200 2098 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 105 nsew signal tristate
flabel metal2 s 9034 26200 9090 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 106 nsew signal tristate
flabel metal2 s 9402 26200 9458 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 107 nsew signal tristate
flabel metal2 s 9770 26200 9826 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 108 nsew signal tristate
flabel metal2 s 10138 26200 10194 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 109 nsew signal tristate
flabel metal2 s 10506 26200 10562 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 110 nsew signal tristate
flabel metal2 s 10874 26200 10930 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 111 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 112 nsew signal tristate
flabel metal2 s 11610 26200 11666 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 113 nsew signal tristate
flabel metal2 s 11978 26200 12034 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 114 nsew signal tristate
flabel metal2 s 12346 26200 12402 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 115 nsew signal tristate
flabel metal2 s 2410 26200 2466 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 116 nsew signal tristate
flabel metal2 s 2778 26200 2834 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 117 nsew signal tristate
flabel metal2 s 3146 26200 3202 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 118 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 119 nsew signal tristate
flabel metal2 s 3882 26200 3938 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 120 nsew signal tristate
flabel metal2 s 4250 26200 4306 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 121 nsew signal tristate
flabel metal2 s 4618 26200 4674 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 122 nsew signal tristate
flabel metal2 s 4986 26200 5042 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 123 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 prog_clk
port 124 nsew signal input
flabel metal2 s 24490 26200 24546 27000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 125 nsew signal input
flabel metal2 s 24858 26200 24914 27000 0 FreeSans 224 90 0 0 reset_top_in
port 126 nsew signal input
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
port 127 nsew signal input
flabel metal3 s 26200 25576 27000 25696 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
port 128 nsew signal input
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
port 129 nsew signal input
flabel metal3 s 26200 26392 27000 26512 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
port 130 nsew signal input
flabel metal2 s 25226 26200 25282 27000 0 FreeSans 224 90 0 0 test_enable_top_in
port 131 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 132 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 133 nsew signal input
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 134 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 135 nsew signal input
rlabel metal1 13478 23936 13478 23936 0 VGND
rlabel metal1 13478 24480 13478 24480 0 VPWR
rlabel metal2 6762 1571 6762 1571 0 ccff_head
rlabel metal3 24894 340 24894 340 0 ccff_tail
rlabel metal1 21666 8466 21666 8466 0 chanx_right_in[0]
rlabel metal3 22977 12852 22977 12852 0 chanx_right_in[10]
rlabel metal2 12466 18071 12466 18071 0 chanx_right_in[11]
rlabel metal1 13892 15334 13892 15334 0 chanx_right_in[12]
rlabel metal1 20010 18292 20010 18292 0 chanx_right_in[13]
rlabel metal1 20378 17646 20378 17646 0 chanx_right_in[14]
rlabel metal2 21758 20621 21758 20621 0 chanx_right_in[15]
rlabel metal1 13432 13906 13432 13906 0 chanx_right_in[16]
rlabel metal1 12834 14552 12834 14552 0 chanx_right_in[17]
rlabel metal2 12834 17884 12834 17884 0 chanx_right_in[18]
rlabel metal1 7452 17170 7452 17170 0 chanx_right_in[19]
rlabel metal1 18952 12750 18952 12750 0 chanx_right_in[1]
rlabel via3 22517 17340 22517 17340 0 chanx_right_in[20]
rlabel metal2 21344 15436 21344 15436 0 chanx_right_in[21]
rlabel metal3 19619 12580 19619 12580 0 chanx_right_in[22]
rlabel metal2 20516 16116 20516 16116 0 chanx_right_in[23]
rlabel metal3 17917 13668 17917 13668 0 chanx_right_in[24]
rlabel metal2 15686 16014 15686 16014 0 chanx_right_in[25]
rlabel metal2 13754 14535 13754 14535 0 chanx_right_in[26]
rlabel metal3 18492 23800 18492 23800 0 chanx_right_in[27]
rlabel metal2 17066 23732 17066 23732 0 chanx_right_in[28]
rlabel metal2 9522 15300 9522 15300 0 chanx_right_in[29]
rlabel metal1 21712 9690 21712 9690 0 chanx_right_in[2]
rlabel metal3 24848 14212 24848 14212 0 chanx_right_in[3]
rlabel metal2 18906 13090 18906 13090 0 chanx_right_in[4]
rlabel metal2 22770 14637 22770 14637 0 chanx_right_in[5]
rlabel metal2 20194 14064 20194 14064 0 chanx_right_in[6]
rlabel metal2 24840 12852 24840 12852 0 chanx_right_in[7]
rlabel metal1 23184 17578 23184 17578 0 chanx_right_in[8]
rlabel metal1 19412 13430 19412 13430 0 chanx_right_in[9]
rlabel metal3 25722 748 25722 748 0 chanx_right_out[0]
rlabel metal1 23322 5100 23322 5100 0 chanx_right_out[10]
rlabel metal2 24794 4641 24794 4641 0 chanx_right_out[11]
rlabel metal3 25676 5644 25676 5644 0 chanx_right_out[12]
rlabel metal1 24104 6358 24104 6358 0 chanx_right_out[13]
rlabel metal2 24702 5797 24702 5797 0 chanx_right_out[14]
rlabel metal1 24380 6834 24380 6834 0 chanx_right_out[15]
rlabel metal1 24104 7446 24104 7446 0 chanx_right_out[16]
rlabel metal2 24794 6953 24794 6953 0 chanx_right_out[17]
rlabel metal1 24426 7922 24426 7922 0 chanx_right_out[18]
rlabel metal1 24012 8398 24012 8398 0 chanx_right_out[19]
rlabel metal3 24250 1156 24250 1156 0 chanx_right_out[1]
rlabel metal2 25162 8177 25162 8177 0 chanx_right_out[20]
rlabel metal1 24380 9010 24380 9010 0 chanx_right_out[21]
rlabel metal2 23322 9673 23322 9673 0 chanx_right_out[22]
rlabel metal1 24794 8364 24794 8364 0 chanx_right_out[23]
rlabel metal1 24104 10710 24104 10710 0 chanx_right_out[24]
rlabel metal2 24794 10217 24794 10217 0 chanx_right_out[25]
rlabel metal1 24380 11186 24380 11186 0 chanx_right_out[26]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[27]
rlabel metal2 24702 11373 24702 11373 0 chanx_right_out[28]
rlabel metal3 25584 12580 25584 12580 0 chanx_right_out[29]
rlabel metal3 24250 1564 24250 1564 0 chanx_right_out[2]
rlabel metal1 20884 2618 20884 2618 0 chanx_right_out[3]
rlabel metal3 25676 2380 25676 2380 0 chanx_right_out[4]
rlabel metal1 24104 3094 24104 3094 0 chanx_right_out[5]
rlabel metal3 25768 3196 25768 3196 0 chanx_right_out[6]
rlabel metal1 23322 4012 23322 4012 0 chanx_right_out[7]
rlabel metal1 25208 3094 25208 3094 0 chanx_right_out[8]
rlabel metal3 25676 4420 25676 4420 0 chanx_right_out[9]
rlabel metal2 2898 18700 2898 18700 0 chany_top_in[0]
rlabel metal1 13570 23256 13570 23256 0 chany_top_in[10]
rlabel metal1 16376 19346 16376 19346 0 chany_top_in[11]
rlabel metal1 17480 18938 17480 18938 0 chany_top_in[12]
rlabel metal2 17112 21012 17112 21012 0 chany_top_in[13]
rlabel metal1 16698 16524 16698 16524 0 chany_top_in[14]
rlabel metal1 15088 14994 15088 14994 0 chany_top_in[15]
rlabel metal2 18630 24745 18630 24745 0 chany_top_in[16]
rlabel metal2 18998 25493 18998 25493 0 chany_top_in[17]
rlabel metal2 19366 24762 19366 24762 0 chany_top_in[18]
rlabel metal2 19642 22899 19642 22899 0 chany_top_in[19]
rlabel metal2 13386 20111 13386 20111 0 chany_top_in[1]
rlabel metal2 19826 26248 19826 26248 0 chany_top_in[20]
rlabel via1 20194 26299 20194 26299 0 chany_top_in[21]
rlabel metal2 13938 21954 13938 21954 0 chany_top_in[22]
rlabel metal3 16560 22372 16560 22372 0 chany_top_in[23]
rlabel via1 21298 26333 21298 26333 0 chany_top_in[24]
rlabel metal2 21942 25221 21942 25221 0 chany_top_in[25]
rlabel metal2 2162 22457 2162 22457 0 chany_top_in[26]
rlabel metal2 10074 15521 10074 15521 0 chany_top_in[27]
rlabel metal1 20976 11254 20976 11254 0 chany_top_in[28]
rlabel metal1 16376 11118 16376 11118 0 chany_top_in[29]
rlabel metal2 12558 22712 12558 22712 0 chany_top_in[2]
rlabel metal2 13846 25153 13846 25153 0 chany_top_in[3]
rlabel metal1 13294 23120 13294 23120 0 chany_top_in[4]
rlabel metal2 14582 25204 14582 25204 0 chany_top_in[5]
rlabel metal2 13662 23392 13662 23392 0 chany_top_in[6]
rlabel metal1 16330 20026 16330 20026 0 chany_top_in[7]
rlabel metal2 15686 24541 15686 24541 0 chany_top_in[8]
rlabel metal2 16284 21964 16284 21964 0 chany_top_in[9]
rlabel metal1 1978 19278 1978 19278 0 chany_top_out[0]
rlabel metal1 4600 23766 4600 23766 0 chany_top_out[10]
rlabel metal2 5750 24490 5750 24490 0 chany_top_out[11]
rlabel metal2 6118 24184 6118 24184 0 chany_top_out[12]
rlabel metal1 4738 24242 4738 24242 0 chany_top_out[13]
rlabel metal1 7222 20978 7222 20978 0 chany_top_out[14]
rlabel metal2 7268 21454 7268 21454 0 chany_top_out[15]
rlabel metal1 6716 23766 6716 23766 0 chany_top_out[16]
rlabel metal1 6394 22984 6394 22984 0 chany_top_out[17]
rlabel metal2 8326 24184 8326 24184 0 chany_top_out[18]
rlabel metal1 7268 24106 7268 24106 0 chany_top_out[19]
rlabel metal1 2300 19890 2300 19890 0 chany_top_out[1]
rlabel metal2 8786 24497 8786 24497 0 chany_top_out[20]
rlabel metal1 8786 23086 8786 23086 0 chany_top_out[21]
rlabel metal1 8970 24242 8970 24242 0 chany_top_out[22]
rlabel metal1 9660 23766 9660 23766 0 chany_top_out[23]
rlabel metal2 10534 24728 10534 24728 0 chany_top_out[24]
rlabel metal2 10902 25034 10902 25034 0 chany_top_out[25]
rlabel metal1 11132 24242 11132 24242 0 chany_top_out[26]
rlabel metal1 11914 23154 11914 23154 0 chany_top_out[27]
rlabel metal2 12006 24966 12006 24966 0 chany_top_out[28]
rlabel metal1 12834 24276 12834 24276 0 chany_top_out[29]
rlabel metal2 2438 24218 2438 24218 0 chany_top_out[2]
rlabel metal1 3220 26418 3220 26418 0 chany_top_out[3]
rlabel metal2 3029 26316 3029 26316 0 chany_top_out[4]
rlabel metal2 3542 23878 3542 23878 0 chany_top_out[5]
rlabel metal1 4370 20978 4370 20978 0 chany_top_out[6]
rlabel metal1 4140 22678 4140 22678 0 chany_top_out[7]
rlabel metal1 3818 23018 3818 23018 0 chany_top_out[8]
rlabel metal2 5067 26316 5067 26316 0 chany_top_out[9]
rlabel metal1 21436 14382 21436 14382 0 clknet_0_prog_clk
rlabel metal1 10488 13158 10488 13158 0 clknet_3_0__leaf_prog_clk
rlabel metal1 15640 15538 15640 15538 0 clknet_3_1__leaf_prog_clk
rlabel metal2 9062 20978 9062 20978 0 clknet_3_2__leaf_prog_clk
rlabel metal1 12190 19346 12190 19346 0 clknet_3_3__leaf_prog_clk
rlabel metal1 19458 14042 19458 14042 0 clknet_3_4__leaf_prog_clk
rlabel metal1 21896 16626 21896 16626 0 clknet_3_5__leaf_prog_clk
rlabel metal1 19412 20910 19412 20910 0 clknet_3_6__leaf_prog_clk
rlabel metal1 23368 21522 23368 21522 0 clknet_3_7__leaf_prog_clk
rlabel metal2 6854 5746 6854 5746 0 net1
rlabel via2 13478 14773 13478 14773 0 net10
rlabel metal1 24472 14246 24472 14246 0 net100
rlabel metal3 22793 15300 22793 15300 0 net101
rlabel metal2 13202 21539 13202 21539 0 net102
rlabel metal1 14237 23766 14237 23766 0 net103
rlabel metal1 11776 22066 11776 22066 0 net104
rlabel metal1 6440 17850 6440 17850 0 net105
rlabel metal1 3082 24174 3082 24174 0 net106
rlabel metal1 7406 17850 7406 17850 0 net107
rlabel metal1 7636 17306 7636 17306 0 net108
rlabel metal2 12650 23664 12650 23664 0 net109
rlabel metal1 14950 24072 14950 24072 0 net11
rlabel via2 18630 23035 18630 23035 0 net110
rlabel metal2 18998 21913 18998 21913 0 net111
rlabel metal1 5750 24174 5750 24174 0 net112
rlabel via2 16330 19669 16330 19669 0 net113
rlabel metal1 3266 18632 3266 18632 0 net114
rlabel metal1 5888 18938 5888 18938 0 net115
rlabel metal1 3634 20570 3634 20570 0 net116
rlabel metal1 5152 19346 5152 19346 0 net117
rlabel metal1 7452 18802 7452 18802 0 net118
rlabel metal1 6670 19754 6670 19754 0 net119
rlabel metal4 15180 18428 15180 18428 0 net12
rlabel metal1 8464 19822 8464 19822 0 net120
rlabel metal1 11730 23018 11730 23018 0 net121
rlabel metal1 5842 17714 5842 17714 0 net122
rlabel metal2 12650 19108 12650 19108 0 net123
rlabel metal2 2254 21284 2254 21284 0 net124
rlabel metal2 15962 20281 15962 20281 0 net125
rlabel metal1 2254 21964 2254 21964 0 net126
rlabel metal1 3588 21522 3588 21522 0 net127
rlabel metal1 5796 18394 5796 18394 0 net128
rlabel metal1 4186 18394 4186 18394 0 net129
rlabel metal2 14076 16626 14076 16626 0 net13
rlabel metal1 12512 21046 12512 21046 0 net130
rlabel metal1 16100 22610 16100 22610 0 net131
rlabel metal1 20792 15402 20792 15402 0 net132
rlabel metal1 19734 14314 19734 14314 0 net133
rlabel metal1 4784 18190 4784 18190 0 net134
rlabel metal1 17710 12274 17710 12274 0 net135
rlabel metal1 18952 12818 18952 12818 0 net136
rlabel metal1 21160 12818 21160 12818 0 net137
rlabel metal1 24104 9962 24104 9962 0 net138
rlabel metal1 18400 10710 18400 10710 0 net139
rlabel metal1 19412 9418 19412 9418 0 net14
rlabel metal2 22494 14858 22494 14858 0 net140
rlabel metal1 20332 17306 20332 17306 0 net141
rlabel metal1 14260 19822 14260 19822 0 net142
rlabel metal2 10074 21760 10074 21760 0 net143
rlabel metal1 8418 22746 8418 22746 0 net144
rlabel metal1 9062 20570 9062 20570 0 net145
rlabel metal1 9614 19754 9614 19754 0 net146
rlabel metal1 19274 18802 19274 18802 0 net147
rlabel metal1 9384 18734 9384 18734 0 net148
rlabel via2 12466 20587 12466 20587 0 net149
rlabel metal2 17756 13362 17756 13362 0 net15
rlabel metal1 12144 18394 12144 18394 0 net150
rlabel metal1 11040 16558 11040 16558 0 net151
rlabel metal1 15456 15062 15456 15062 0 net152
rlabel metal1 10488 16218 10488 16218 0 net153
rlabel metal1 13478 15470 13478 15470 0 net154
rlabel metal1 13984 15062 13984 15062 0 net155
rlabel metal1 14030 17714 14030 17714 0 net156
rlabel metal1 5152 20570 5152 20570 0 net157
rlabel metal1 14766 23834 14766 23834 0 net158
rlabel metal1 21206 19414 21206 19414 0 net159
rlabel metal1 17572 10506 17572 10506 0 net16
rlabel metal1 20838 14892 20838 14892 0 net160
rlabel metal1 23230 16150 23230 16150 0 net161
rlabel metal1 24196 16082 24196 16082 0 net162
rlabel metal2 24886 13668 24886 13668 0 net163
rlabel metal1 25116 13226 25116 13226 0 net164
rlabel metal2 2254 19159 2254 19159 0 net165
rlabel metal1 21160 14042 21160 14042 0 net166
rlabel metal1 21436 15470 21436 15470 0 net167
rlabel metal1 17940 13702 17940 13702 0 net17
rlabel metal2 19642 21556 19642 21556 0 net18
rlabel metal1 16100 11322 16100 11322 0 net19
rlabel metal3 16445 18836 16445 18836 0 net2
rlabel metal1 12466 13804 12466 13804 0 net20
rlabel metal2 18446 14824 18446 14824 0 net21
rlabel metal2 19642 17136 19642 17136 0 net22
rlabel metal2 14398 22763 14398 22763 0 net23
rlabel metal3 15985 19380 15985 19380 0 net24
rlabel metal3 17641 16660 17641 16660 0 net25
rlabel metal1 19228 13498 19228 13498 0 net26
rlabel metal1 17112 17170 17112 17170 0 net27
rlabel metal1 16054 16082 16054 16082 0 net28
rlabel metal2 12834 14416 12834 14416 0 net29
rlabel metal3 13639 20740 13639 20740 0 net3
rlabel metal1 20930 16966 20930 16966 0 net30
rlabel metal1 16008 23698 16008 23698 0 net31
rlabel metal2 1610 18615 1610 18615 0 net32
rlabel metal2 20102 15215 20102 15215 0 net33
rlabel metal2 16330 18037 16330 18037 0 net34
rlabel metal1 21942 15470 21942 15470 0 net35
rlabel metal2 19734 18105 19734 18105 0 net36
rlabel metal1 16606 16762 16606 16762 0 net37
rlabel metal2 14858 14841 14858 14841 0 net38
rlabel via2 20930 18309 20930 18309 0 net39
rlabel metal2 8418 17408 8418 17408 0 net4
rlabel metal2 9430 17544 9430 17544 0 net40
rlabel metal2 7682 16541 7682 16541 0 net41
rlabel metal2 8878 17867 8878 17867 0 net42
rlabel via2 18722 12155 18722 12155 0 net43
rlabel metal4 18492 14620 18492 14620 0 net44
rlabel metal2 5198 18649 5198 18649 0 net45
rlabel metal4 16468 18224 16468 18224 0 net46
rlabel metal4 19596 18224 19596 18224 0 net47
rlabel metal2 21022 20315 21022 20315 0 net48
rlabel via2 9154 15963 9154 15963 0 net49
rlabel metal1 13294 14586 13294 14586 0 net5
rlabel metal2 1978 21930 1978 21930 0 net50
rlabel metal1 13018 15504 13018 15504 0 net51
rlabel via2 19458 10251 19458 10251 0 net52
rlabel via2 16146 11237 16146 11237 0 net53
rlabel via2 19734 11067 19734 11067 0 net54
rlabel metal2 6578 15623 6578 15623 0 net55
rlabel metal1 25806 14586 25806 14586 0 net56
rlabel metal1 20746 16218 20746 16218 0 net57
rlabel metal1 19872 17714 19872 17714 0 net58
rlabel metal2 18538 19380 18538 19380 0 net59
rlabel metal2 16606 19601 16606 19601 0 net6
rlabel metal3 13478 18428 13478 18428 0 net60
rlabel metal1 23414 21862 23414 21862 0 net61
rlabel metal1 11829 8874 11829 8874 0 net62
rlabel metal2 17480 21522 17480 21522 0 net63
rlabel metal1 20240 18598 20240 18598 0 net64
rlabel metal1 20010 17510 20010 17510 0 net65
rlabel metal1 20976 19414 20976 19414 0 net66
rlabel metal1 14766 18870 14766 18870 0 net67
rlabel via2 7130 23579 7130 23579 0 net68
rlabel metal2 19918 22338 19918 22338 0 net69
rlabel metal1 8694 17034 8694 17034 0 net7
rlabel metal1 14996 18666 14996 18666 0 net70
rlabel metal1 21528 2414 21528 2414 0 net71
rlabel metal1 19872 3026 19872 3026 0 net72
rlabel metal1 22448 14790 22448 14790 0 net73
rlabel metal1 24012 15538 24012 15538 0 net74
rlabel metal1 23184 5678 23184 5678 0 net75
rlabel metal2 22310 7718 22310 7718 0 net76
rlabel metal2 20930 7106 20930 7106 0 net77
rlabel metal1 21390 6664 21390 6664 0 net78
rlabel metal1 25392 17034 25392 17034 0 net79
rlabel metal2 13018 22542 13018 22542 0 net8
rlabel metal1 25254 16626 25254 16626 0 net80
rlabel metal1 25438 17578 25438 17578 0 net81
rlabel metal1 24978 15946 24978 15946 0 net82
rlabel metal1 20700 3502 20700 3502 0 net83
rlabel metal2 20746 7582 20746 7582 0 net84
rlabel metal2 22678 8228 22678 8228 0 net85
rlabel metal2 20746 9826 20746 9826 0 net86
rlabel metal2 20010 8976 20010 8976 0 net87
rlabel metal1 18791 12954 18791 12954 0 net88
rlabel metal2 22494 10030 22494 10030 0 net89
rlabel metal1 13110 13804 13110 13804 0 net9
rlabel metal2 18078 9248 18078 9248 0 net90
rlabel metal1 19688 8602 19688 8602 0 net91
rlabel metal2 21942 10846 21942 10846 0 net92
rlabel metal2 23966 9894 23966 9894 0 net93
rlabel metal1 21114 4114 21114 4114 0 net94
rlabel metal1 18446 3060 18446 3060 0 net95
rlabel metal1 23736 2414 23736 2414 0 net96
rlabel metal1 22954 3026 22954 3026 0 net97
rlabel metal1 23184 3502 23184 3502 0 net98
rlabel metal1 22862 4114 22862 4114 0 net99
rlabel metal1 19596 4046 19596 4046 0 prog_clk
rlabel metal2 24334 25075 24334 25075 0 prog_reset_top_in
rlabel metal2 24794 24497 24794 24497 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 21988 24378 21988 24378 0 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 23230 22100 23230 22100 0 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 21850 22610 21850 22610 0 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 15548 17714 15548 17714 0 sb_0__0_.mem_right_track_0.ccff_head
rlabel metal2 19918 19822 19918 19822 0 sb_0__0_.mem_right_track_0.ccff_tail
rlabel metal2 17342 18530 17342 18530 0 sb_0__0_.mem_right_track_0.mem_out\[0\]
rlabel metal2 25254 19516 25254 19516 0 sb_0__0_.mem_right_track_10.ccff_head
rlabel metal2 21390 19584 21390 19584 0 sb_0__0_.mem_right_track_10.ccff_tail
rlabel metal2 25070 18326 25070 18326 0 sb_0__0_.mem_right_track_10.mem_out\[0\]
rlabel metal2 22402 17442 22402 17442 0 sb_0__0_.mem_right_track_12.ccff_tail
rlabel metal2 21942 19414 21942 19414 0 sb_0__0_.mem_right_track_12.mem_out\[0\]
rlabel metal1 23966 15980 23966 15980 0 sb_0__0_.mem_right_track_14.ccff_tail
rlabel metal1 22586 17850 22586 17850 0 sb_0__0_.mem_right_track_14.mem_out\[0\]
rlabel metal1 24564 13838 24564 13838 0 sb_0__0_.mem_right_track_16.ccff_tail
rlabel metal1 24380 15130 24380 15130 0 sb_0__0_.mem_right_track_16.mem_out\[0\]
rlabel metal1 23138 12954 23138 12954 0 sb_0__0_.mem_right_track_18.ccff_tail
rlabel metal1 22540 12750 22540 12750 0 sb_0__0_.mem_right_track_18.mem_out\[0\]
rlabel metal2 22034 21454 22034 21454 0 sb_0__0_.mem_right_track_2.ccff_tail
rlabel metal1 20930 20570 20930 20570 0 sb_0__0_.mem_right_track_2.mem_out\[0\]
rlabel metal1 21298 13872 21298 13872 0 sb_0__0_.mem_right_track_28.ccff_tail
rlabel metal1 20010 13192 20010 13192 0 sb_0__0_.mem_right_track_28.mem_out\[0\]
rlabel metal2 19274 16762 19274 16762 0 sb_0__0_.mem_right_track_30.ccff_tail
rlabel metal1 21482 14926 21482 14926 0 sb_0__0_.mem_right_track_30.mem_out\[0\]
rlabel metal1 18078 16422 18078 16422 0 sb_0__0_.mem_right_track_32.ccff_tail
rlabel metal1 21206 21454 21206 21454 0 sb_0__0_.mem_right_track_32.mem_out\[0\]
rlabel metal1 19665 14450 19665 14450 0 sb_0__0_.mem_right_track_34.ccff_tail
rlabel metal2 19366 16898 19366 16898 0 sb_0__0_.mem_right_track_34.mem_out\[0\]
rlabel metal1 25392 18190 25392 18190 0 sb_0__0_.mem_right_track_4.ccff_tail
rlabel metal1 17618 24276 17618 24276 0 sb_0__0_.mem_right_track_4.mem_out\[0\]
rlabel metal1 17204 13158 17204 13158 0 sb_0__0_.mem_right_track_44.ccff_tail
rlabel metal1 18492 14518 18492 14518 0 sb_0__0_.mem_right_track_44.mem_out\[0\]
rlabel metal1 19136 12682 19136 12682 0 sb_0__0_.mem_right_track_46.ccff_tail
rlabel metal1 17756 12750 17756 12750 0 sb_0__0_.mem_right_track_46.mem_out\[0\]
rlabel metal1 20746 12682 20746 12682 0 sb_0__0_.mem_right_track_48.ccff_tail
rlabel metal1 20194 17714 20194 17714 0 sb_0__0_.mem_right_track_48.mem_out\[0\]
rlabel metal1 21436 11594 21436 11594 0 sb_0__0_.mem_right_track_50.mem_out\[0\]
rlabel metal1 24426 21454 24426 21454 0 sb_0__0_.mem_right_track_6.ccff_tail
rlabel metal1 17756 23630 17756 23630 0 sb_0__0_.mem_right_track_6.mem_out\[0\]
rlabel metal1 16882 24242 16882 24242 0 sb_0__0_.mem_right_track_8.mem_out\[0\]
rlabel metal1 15916 18666 15916 18666 0 sb_0__0_.mem_top_track_0.ccff_tail
rlabel metal2 14950 19074 14950 19074 0 sb_0__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 15088 22746 15088 22746 0 sb_0__0_.mem_top_track_10.ccff_head
rlabel metal1 15226 20230 15226 20230 0 sb_0__0_.mem_top_track_10.ccff_tail
rlabel metal1 16146 21862 16146 21862 0 sb_0__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 13202 21454 13202 21454 0 sb_0__0_.mem_top_track_12.ccff_tail
rlabel metal2 14490 19771 14490 19771 0 sb_0__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 12374 22066 12374 22066 0 sb_0__0_.mem_top_track_14.ccff_tail
rlabel metal1 13294 21114 13294 21114 0 sb_0__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 10626 21012 10626 21012 0 sb_0__0_.mem_top_track_16.ccff_tail
rlabel metal2 9338 21182 9338 21182 0 sb_0__0_.mem_top_track_16.mem_out\[0\]
rlabel metal2 10810 18666 10810 18666 0 sb_0__0_.mem_top_track_18.ccff_tail
rlabel metal2 10810 19856 10810 19856 0 sb_0__0_.mem_top_track_18.mem_out\[0\]
rlabel metal1 19136 20978 19136 20978 0 sb_0__0_.mem_top_track_2.ccff_tail
rlabel metal1 17480 20366 17480 20366 0 sb_0__0_.mem_top_track_2.mem_out\[0\]
rlabel metal2 10074 17340 10074 17340 0 sb_0__0_.mem_top_track_28.ccff_tail
rlabel metal1 15778 18122 15778 18122 0 sb_0__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 12512 20196 12512 20196 0 sb_0__0_.mem_top_track_30.ccff_tail
rlabel metal2 13478 19448 13478 19448 0 sb_0__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 12880 16422 12880 16422 0 sb_0__0_.mem_top_track_32.ccff_tail
rlabel metal1 15134 17850 15134 17850 0 sb_0__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 11960 15334 11960 15334 0 sb_0__0_.mem_top_track_34.ccff_tail
rlabel metal2 13478 16337 13478 16337 0 sb_0__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 19550 23630 19550 23630 0 sb_0__0_.mem_top_track_4.ccff_tail
rlabel metal1 20838 21114 20838 21114 0 sb_0__0_.mem_top_track_4.mem_out\[0\]
rlabel metal2 12098 15402 12098 15402 0 sb_0__0_.mem_top_track_44.ccff_tail
rlabel metal1 12466 14382 12466 14382 0 sb_0__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 14398 13226 14398 13226 0 sb_0__0_.mem_top_track_46.ccff_tail
rlabel metal1 13984 13430 13984 13430 0 sb_0__0_.mem_top_track_46.mem_out\[0\]
rlabel metal2 14582 15232 14582 15232 0 sb_0__0_.mem_top_track_48.ccff_tail
rlabel metal1 19918 15980 19918 15980 0 sb_0__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 16330 14246 16330 14246 0 sb_0__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 17894 23426 17894 23426 0 sb_0__0_.mem_top_track_6.ccff_tail
rlabel metal2 19826 23766 19826 23766 0 sb_0__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 15732 22950 15732 22950 0 sb_0__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 24058 15334 24058 15334 0 sb_0__0_.mux_right_track_0.out
rlabel metal2 19734 20400 19734 20400 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20056 19482 20056 19482 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19182 18768 19182 18768 0 sb_0__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15916 12818 15916 12818 0 sb_0__0_.mux_right_track_10.out
rlabel metal1 24196 17646 24196 17646 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23460 17510 23460 17510 0 sb_0__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20516 9554 20516 9554 0 sb_0__0_.mux_right_track_12.out
rlabel metal2 21758 16269 21758 16269 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22218 15878 22218 15878 0 sb_0__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19688 10098 19688 10098 0 sb_0__0_.mux_right_track_14.out
rlabel metal1 23782 16218 23782 16218 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21758 10710 21758 10710 0 sb_0__0_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21298 7378 21298 7378 0 sb_0__0_.mux_right_track_16.out
rlabel metal1 23598 14450 23598 14450 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19780 10642 19780 10642 0 sb_0__0_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19826 7854 19826 7854 0 sb_0__0_.mux_right_track_18.out
rlabel metal1 25162 13294 25162 13294 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20608 11186 20608 11186 0 sb_0__0_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9660 12274 9660 12274 0 sb_0__0_.mux_right_track_2.out
rlabel metal1 23368 20842 23368 20842 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 4738 18989 4738 18989 0 sb_0__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21390 6766 21390 6766 0 sb_0__0_.mux_right_track_28.out
rlabel metal1 21114 13838 21114 13838 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20792 10642 20792 10642 0 sb_0__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19458 9044 19458 9044 0 sb_0__0_.mux_right_track_30.out
rlabel metal2 21206 17527 21206 17527 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21068 15334 21068 15334 0 sb_0__0_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24702 8840 24702 8840 0 sb_0__0_.mux_right_track_32.out
rlabel metal2 20010 18394 20010 18394 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20056 15334 20056 15334 0 sb_0__0_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 25070 9554 25070 9554 0 sb_0__0_.mux_right_track_34.out
rlabel metal2 19918 16184 19918 16184 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20194 14518 20194 14518 0 sb_0__0_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14214 17034 14214 17034 0 sb_0__0_.mux_right_track_4.out
rlabel metal2 16974 24480 16974 24480 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20562 17000 20562 17000 0 sb_0__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24656 6766 24656 6766 0 sb_0__0_.mux_right_track_44.out
rlabel metal1 17572 14042 17572 14042 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17112 14042 17112 14042 0 sb_0__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24610 8296 24610 8296 0 sb_0__0_.mux_right_track_46.out
rlabel metal2 19550 12954 19550 12954 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20010 8398 20010 8398 0 sb_0__0_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23414 5916 23414 5916 0 sb_0__0_.mux_right_track_48.out
rlabel metal1 20286 12750 20286 12750 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20562 7378 20562 7378 0 sb_0__0_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 23690 4658 23690 4658 0 sb_0__0_.mux_right_track_50.out
rlabel metal2 20562 15776 20562 15776 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21850 7956 21850 7956 0 sb_0__0_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13386 9554 13386 9554 0 sb_0__0_.mux_right_track_6.out
rlabel metal2 16882 24072 16882 24072 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24656 20026 24656 20026 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 8694 16099 8694 16099 0 sb_0__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20194 10608 20194 10608 0 sb_0__0_.mux_right_track_8.out
rlabel metal3 18584 20332 18584 20332 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24472 17748 24472 17748 0 sb_0__0_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4554 17034 4554 17034 0 sb_0__0_.mux_top_track_0.out
rlabel metal2 14306 19176 14306 19176 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15870 19482 15870 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14904 19482 14904 19482 0 sb_0__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7774 18734 7774 18734 0 sb_0__0_.mux_top_track_10.out
rlabel metal2 17710 21760 17710 21760 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13018 20332 13018 20332 0 sb_0__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3910 17850 3910 17850 0 sb_0__0_.mux_top_track_12.out
rlabel metal1 16698 20978 16698 20978 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 3450 19346 3450 19346 0 sb_0__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2438 20332 2438 20332 0 sb_0__0_.mux_top_track_14.out
rlabel metal1 16606 21862 16606 21862 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11362 19924 11362 19924 0 sb_0__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7176 18394 7176 18394 0 sb_0__0_.mux_top_track_16.out
rlabel metal1 14168 21046 14168 21046 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 8510 19652 8510 19652 0 sb_0__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3818 18734 3818 18734 0 sb_0__0_.mux_top_track_18.out
rlabel metal1 10902 19924 10902 19924 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8832 20026 8832 20026 0 sb_0__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5198 17748 5198 17748 0 sb_0__0_.mux_top_track_2.out
rlabel metal2 18354 21182 18354 21182 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17802 21046 17802 21046 0 sb_0__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 1610 20128 1610 20128 0 sb_0__0_.mux_top_track_28.out
rlabel metal1 13478 18122 13478 18122 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 1794 20468 1794 20468 0 sb_0__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7958 17680 7958 17680 0 sb_0__0_.mux_top_track_30.out
rlabel metal1 17664 20026 17664 20026 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11546 20570 11546 20570 0 sb_0__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8326 18938 8326 18938 0 sb_0__0_.mux_top_track_32.out
rlabel metal1 16376 18122 16376 18122 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10212 18394 10212 18394 0 sb_0__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6256 17646 6256 17646 0 sb_0__0_.mux_top_track_34.out
rlabel metal2 11270 16660 11270 16660 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10810 16150 10810 16150 0 sb_0__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9430 23052 9430 23052 0 sb_0__0_.mux_top_track_4.out
rlabel metal1 19780 22746 19780 22746 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 17986 24259 17986 24259 0 sb_0__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4738 18292 4738 18292 0 sb_0__0_.mux_top_track_44.out
rlabel metal1 14582 15946 14582 15946 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10442 15980 10442 15980 0 sb_0__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6486 18258 6486 18258 0 sb_0__0_.mux_top_track_46.out
rlabel metal1 13202 15572 13202 15572 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12374 15674 12374 15674 0 sb_0__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8418 19278 8418 19278 0 sb_0__0_.mux_top_track_48.out
rlabel metal1 16882 16218 16882 16218 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13938 15776 13938 15776 0 sb_0__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5474 18258 5474 18258 0 sb_0__0_.mux_top_track_50.out
rlabel metal2 17158 18224 17158 18224 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11270 19380 11270 19380 0 sb_0__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 3956 17306 3956 17306 0 sb_0__0_.mux_top_track_6.out
rlabel metal1 16100 21386 16100 21386 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24518 23664 24518 23664 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel via3 16859 22508 16859 22508 0 sb_0__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 5520 19482 5520 19482 0 sb_0__0_.mux_top_track_8.out
rlabel metal1 19090 22644 19090 22644 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13938 23834 13938 23834 0 sb_0__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 1518 22610 1518 22610 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 1518 23698 1518 23698 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 2806 23783 2806 23783 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal1 1932 21590 1932 21590 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 27000 27000
<< end >>
