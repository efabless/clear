//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: FPGA Verilog Testbench for Top-level netlist of Design: top
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Tue Nov 24 18:04:19 2020
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

module top_autocheck_top_tb;
// ----- Local wires for global ports of FPGA fabric -----
wire [0:0] prog_clk;
wire [0:0] Test_en;
wire [0:0] IO_ISOL_N;
wire [0:0] clk;

// ----- Local wires for I/Os of FPGA fabric -----

wire [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_IN;

wire [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_OUT;
wire [0:95] gfpga_pad_EMBEDDED_IO_HD_SOC_DIR;

reg [0:0] config_done;
wire [0:0] prog_clock;
reg [0:0] prog_clock_reg;
wire [0:0] op_clock;
reg [0:0] op_clock_reg;
reg [0:0] prog_reset;
reg [0:0] prog_set;
reg [0:0] greset;
reg [0:0] gset;
// ---- Configuration-chain head -----
reg [0:0] ccff_head;
// ---- Configuration-chain tail -----
wire [0:0] ccff_tail;
// ----- Shared inputs -------
	reg [0:0] a;
	reg [0:0] b;

// ----- FPGA fabric outputs -------
	wire [0:0] out:c_fpga;

`ifdef AUTOCHECKED_SIMULATION

// ----- Benchmark outputs -------
	wire [0:0] out:c_benchmark;

// ----- Output vectors checking flags -------
	reg [0:0] out:c_flag;

`endif

// ----- Error counter: Deposit an error for config_done signal is not raised at the beginning -----
	integer nb_error= 1;
// ----- Number of clock cycles in configuration phase: 29697 -----
// ----- Begin configuration done signal generation -----
initial
	begin
		config_done[0] = 1'b0;
	end

// ----- End configuration done signal generation -----

// ----- Begin raw programming clock signal generation -----
initial
	begin
		prog_clock_reg[0] = 1'b0;
	end
always
	begin
		#5	prog_clock_reg[0] = ~prog_clock_reg[0];
	end

// ----- End raw programming clock signal generation -----

// ----- Actual programming clock is triggered only when config_done and prog_reset are disabled -----
	assign prog_clock[0] = prog_clock_reg[0] & (~config_done[0]) & (~prog_reset[0]);

// ----- Begin raw operating clock signal generation -----
initial
	begin
		op_clock_reg[0] = 1'b0;
	end
always wait(~greset)
	begin
		#0.4159859717	op_clock_reg[0] = ~op_clock_reg[0];
	end

// ----- End raw operating clock signal generation -----
// ----- Actual operating clock is triggered only when config_done is enabled -----
	assign op_clock[0] = op_clock_reg[0] & config_done[0];

// ----- Begin programming reset signal generation -----
initial
	begin
		prog_reset[0] = 1'b1;
	#10	prog_reset[0] = 1'b0;
	end

// ----- End programming reset signal generation -----

// ----- Begin programming set signal generation -----
initial
	begin
		prog_set[0] = 1'b1;
	#10	prog_set[0] = 1'b0;
	end

// ----- End programming set signal generation -----

// ----- Begin operating reset signal generation -----
// ----- Reset signal is enabled until the first clock cycle in operation phase -----
initial
	begin
		greset[0] = 1'b1;
	wait(config_done)
	#0.8319719434	greset[0] = 1'b1;
	#1.663943887	greset[0] = 1'b0;
	end

// ----- End operating reset signal generation -----
// ----- Begin operating set signal generation: always disabled -----
initial
	begin
		gset[0] = 1'b0;
	end

// ----- End operating set signal generation: always disabled -----

// ----- Begin connecting global ports of FPGA fabric to stimuli -----
	assign prog_clk[0] = prog_clock[0];
	assign clk[0] = op_clock[0];
	assign Test_en[0] = 1'b0;
	assign IO_ISOL_N[0] = 1'b1;
// ----- End connecting global ports of FPGA fabric to stimuli -----
// ----- FPGA top-level module to be capsulated -----
	fpga_top FPGA_DUT (
		.prog_clk(prog_clk[0]),
		.Test_en(Test_en[0]),
		.IO_ISOL_N(IO_ISOL_N[0]),
		.clk(clk[0]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_IN(gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0:95]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_OUT(gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0:95]),
		.gfpga_pad_EMBEDDED_IO_HD_SOC_DIR(gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0:95]),
		.ccff_head(ccff_head[0]),
		.ccff_tail(ccff_tail[0]));

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input a is mapped to FPGA IOPAD gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4] -----
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4] = a[0];

// ----- Blif Benchmark input b is mapped to FPGA IOPAD gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3] -----
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3] = b[0];

// ----- Blif Benchmark output out:c is mapped to FPGA IOPAD gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5] -----
	assign out:c_fpga[0] = gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95] = 1'b0;

	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94] = 1'b0;
	assign gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95] = 1'b0;

`ifdef AUTOCHECKED_SIMULATION
// ----- Reference Benchmark Instanication -------
	top REF_DUT(
		.a(a),
		.b(b),
		.c(out:c_benchmark)	);
// ----- End reference Benchmark Instanication -------

`endif


// ----- Task: input values during a programming clock cycle -----
task prog_cycle_task;
input [0:0] ccff_head_val;
	begin
		@(negedge prog_clock[0]);
			ccff_head[0] = ccff_head_val[0];
	end
endtask

// ----- Begin bitstream loading during configuration phase -----
initial
	begin
// ----- Configuration chain default input -----
		ccff_head[0] = 1'b0;
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b1);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		prog_cycle_task(1'b0);
		@(negedge prog_clock[0]);
			config_done[0] <= 1'b1;
	end
// ----- End bitstream loading during configuration phase -----
// ----- Input Initialization -------
	initial begin
		a <= 1'b0;
		b <= 1'b0;

		out:c_flag[0] <= 1'b0;
	end

// ----- Input Stimulus -------
	always@(negedge op_clock[0]) begin
		a <= $random;
		b <= $random;
	end

`ifdef AUTOCHECKED_SIMULATION
// ----- Begin checking output vectors -------
// ----- Skip the first falling edge of clock, it is for initialization -------
	reg [0:0] sim_start;

	always@(negedge op_clock[0]) begin
		if (1'b1 == sim_start[0]) begin
			sim_start[0] <= ~sim_start[0];
		end else begin
			if(!(out:c_fpga === out:c_benchmark) && !(out:c_benchmark === 1'bx)) begin
				out:c_flag <= 1'b1;
			end else begin
				out:c_flag<= 1'b0;
			end
		end
	end

	always@(posedge out:c_flag) begin
		if(out:c_flag) begin
			nb_error = nb_error + 1;
			$display("Mismatch on out:c_fpga at time = %t", $realtime);
		end
	end

`endif

`ifdef AUTOCHECKED_SIMULATION
// ----- Configuration done must be raised in the end -------
	always@(posedge config_done[0]) begin
		nb_error = nb_error - 1;
	end
`endif

`ifdef ICARUS_SIMULATOR
// ----- Begin Icarus requirement -------
	initial begin
		$dumpfile("top_formal.vcd");
		$dumpvars(1, top_autocheck_top_tb);
	end
`endif
// ----- END Icarus requirement -------

initial begin
	sim_start[0] <= 1'b1;
	$timeformat(-9, 2, "ns", 20);
	$display("Simulation start");
// ----- Can be changed by the user for his/her need -------
	#296991
	if(nb_error == 0) begin
		$display("Simulation Succeed");
	end else begin
		$display("Simulation Failed with %d error(s)", nb_error);
	end
	$finish;
end

endmodule
// ----- END Verilog module for top_autocheck_top_tb -----

