magic
tech sky130A
magscale 1 2
timestamp 1625785451
<< viali >>
rect 9137 5117 9171 5151
rect 2697 4165 2731 4199
rect 3893 4165 3927 4199
rect 8677 4029 8711 4063
rect 9597 4029 9631 4063
rect 9781 3961 9815 3995
rect 5181 3417 5215 3451
rect 2697 3349 2731 3383
rect 6745 3349 6779 3383
rect 8217 3349 8251 3383
rect 7389 2941 7423 2975
rect 8493 2941 8527 2975
rect 9597 2941 9631 2975
rect 7205 2873 7239 2907
rect 8309 2873 8343 2907
rect 9689 2805 9723 2839
rect 1593 2533 1627 2567
rect 2697 2533 2731 2567
rect 4813 2533 4847 2567
rect 7481 2533 7515 2567
rect 1409 2329 1443 2363
rect 2513 2329 2547 2363
rect 4629 2329 4663 2363
rect 7297 2329 7331 2363
<< metal1 >>
rect 1104 11450 10856 11472
rect 1104 11398 4246 11450
rect 4298 11398 4310 11450
rect 4362 11398 4374 11450
rect 4426 11398 4438 11450
rect 4490 11398 7510 11450
rect 7562 11398 7574 11450
rect 7626 11398 7638 11450
rect 7690 11398 7702 11450
rect 7754 11398 10856 11450
rect 1104 11376 10856 11398
rect 1104 10906 10856 10928
rect 1104 10854 2614 10906
rect 2666 10854 2678 10906
rect 2730 10854 2742 10906
rect 2794 10854 2806 10906
rect 2858 10854 5878 10906
rect 5930 10854 5942 10906
rect 5994 10854 6006 10906
rect 6058 10854 6070 10906
rect 6122 10854 9142 10906
rect 9194 10854 9206 10906
rect 9258 10854 9270 10906
rect 9322 10854 9334 10906
rect 9386 10854 10856 10906
rect 1104 10832 10856 10854
rect 1104 10362 10856 10384
rect 1104 10310 4246 10362
rect 4298 10310 4310 10362
rect 4362 10310 4374 10362
rect 4426 10310 4438 10362
rect 4490 10310 7510 10362
rect 7562 10310 7574 10362
rect 7626 10310 7638 10362
rect 7690 10310 7702 10362
rect 7754 10310 10856 10362
rect 1104 10288 10856 10310
rect 1104 9818 10856 9840
rect 1104 9766 2614 9818
rect 2666 9766 2678 9818
rect 2730 9766 2742 9818
rect 2794 9766 2806 9818
rect 2858 9766 5878 9818
rect 5930 9766 5942 9818
rect 5994 9766 6006 9818
rect 6058 9766 6070 9818
rect 6122 9766 9142 9818
rect 9194 9766 9206 9818
rect 9258 9766 9270 9818
rect 9322 9766 9334 9818
rect 9386 9766 10856 9818
rect 1104 9744 10856 9766
rect 1104 9274 10856 9296
rect 1104 9222 4246 9274
rect 4298 9222 4310 9274
rect 4362 9222 4374 9274
rect 4426 9222 4438 9274
rect 4490 9222 7510 9274
rect 7562 9222 7574 9274
rect 7626 9222 7638 9274
rect 7690 9222 7702 9274
rect 7754 9222 10856 9274
rect 1104 9200 10856 9222
rect 1104 8730 10856 8752
rect 1104 8678 2614 8730
rect 2666 8678 2678 8730
rect 2730 8678 2742 8730
rect 2794 8678 2806 8730
rect 2858 8678 5878 8730
rect 5930 8678 5942 8730
rect 5994 8678 6006 8730
rect 6058 8678 6070 8730
rect 6122 8678 9142 8730
rect 9194 8678 9206 8730
rect 9258 8678 9270 8730
rect 9322 8678 9334 8730
rect 9386 8678 10856 8730
rect 1104 8656 10856 8678
rect 1104 8186 10856 8208
rect 1104 8134 4246 8186
rect 4298 8134 4310 8186
rect 4362 8134 4374 8186
rect 4426 8134 4438 8186
rect 4490 8134 7510 8186
rect 7562 8134 7574 8186
rect 7626 8134 7638 8186
rect 7690 8134 7702 8186
rect 7754 8134 10856 8186
rect 1104 8112 10856 8134
rect 1104 7642 10856 7664
rect 1104 7590 2614 7642
rect 2666 7590 2678 7642
rect 2730 7590 2742 7642
rect 2794 7590 2806 7642
rect 2858 7590 5878 7642
rect 5930 7590 5942 7642
rect 5994 7590 6006 7642
rect 6058 7590 6070 7642
rect 6122 7590 9142 7642
rect 9194 7590 9206 7642
rect 9258 7590 9270 7642
rect 9322 7590 9334 7642
rect 9386 7590 10856 7642
rect 1104 7568 10856 7590
rect 1104 7098 10856 7120
rect 1104 7046 4246 7098
rect 4298 7046 4310 7098
rect 4362 7046 4374 7098
rect 4426 7046 4438 7098
rect 4490 7046 7510 7098
rect 7562 7046 7574 7098
rect 7626 7046 7638 7098
rect 7690 7046 7702 7098
rect 7754 7046 10856 7098
rect 1104 7024 10856 7046
rect 1104 6554 10856 6576
rect 1104 6502 2614 6554
rect 2666 6502 2678 6554
rect 2730 6502 2742 6554
rect 2794 6502 2806 6554
rect 2858 6502 5878 6554
rect 5930 6502 5942 6554
rect 5994 6502 6006 6554
rect 6058 6502 6070 6554
rect 6122 6502 9142 6554
rect 9194 6502 9206 6554
rect 9258 6502 9270 6554
rect 9322 6502 9334 6554
rect 9386 6502 10856 6554
rect 1104 6480 10856 6502
rect 1104 6010 10856 6032
rect 1104 5958 4246 6010
rect 4298 5958 4310 6010
rect 4362 5958 4374 6010
rect 4426 5958 4438 6010
rect 4490 5958 7510 6010
rect 7562 5958 7574 6010
rect 7626 5958 7638 6010
rect 7690 5958 7702 6010
rect 7754 5958 10856 6010
rect 1104 5936 10856 5958
rect 1104 5466 10856 5488
rect 1104 5414 2614 5466
rect 2666 5414 2678 5466
rect 2730 5414 2742 5466
rect 2794 5414 2806 5466
rect 2858 5414 5878 5466
rect 5930 5414 5942 5466
rect 5994 5414 6006 5466
rect 6058 5414 6070 5466
rect 6122 5414 9142 5466
rect 9194 5414 9206 5466
rect 9258 5414 9270 5466
rect 9322 5414 9334 5466
rect 9386 5414 10856 5466
rect 1104 5392 10856 5414
rect 9125 5151 9183 5157
rect 9125 5117 9137 5151
rect 9171 5148 9183 5151
rect 9582 5148 9588 5160
rect 9171 5120 9588 5148
rect 9171 5117 9183 5120
rect 9125 5111 9183 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 1104 4922 10856 4944
rect 1104 4870 4246 4922
rect 4298 4870 4310 4922
rect 4362 4870 4374 4922
rect 4426 4870 4438 4922
rect 4490 4870 7510 4922
rect 7562 4870 7574 4922
rect 7626 4870 7638 4922
rect 7690 4870 7702 4922
rect 7754 4870 10856 4922
rect 1104 4848 10856 4870
rect 1104 4378 10856 4400
rect 1104 4326 2614 4378
rect 2666 4326 2678 4378
rect 2730 4326 2742 4378
rect 2794 4326 2806 4378
rect 2858 4326 5878 4378
rect 5930 4326 5942 4378
rect 5994 4326 6006 4378
rect 6058 4326 6070 4378
rect 6122 4326 9142 4378
rect 9194 4326 9206 4378
rect 9258 4326 9270 4378
rect 9322 4326 9334 4378
rect 9386 4326 10856 4378
rect 1104 4304 10856 4326
rect 2498 4156 2504 4208
rect 2556 4196 2562 4208
rect 2685 4199 2743 4205
rect 2685 4196 2697 4199
rect 2556 4168 2697 4196
rect 2556 4156 2562 4168
rect 2685 4165 2697 4168
rect 2731 4165 2743 4199
rect 2685 4159 2743 4165
rect 3881 4199 3939 4205
rect 3881 4165 3893 4199
rect 3927 4196 3939 4199
rect 4798 4196 4804 4208
rect 3927 4168 4804 4196
rect 3927 4165 3939 4168
rect 3881 4159 3939 4165
rect 4798 4156 4804 4168
rect 4856 4156 4862 4208
rect 8662 4060 8668 4072
rect 8623 4032 8668 4060
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9582 4060 9588 4072
rect 9543 4032 9588 4060
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 9769 3995 9827 4001
rect 9769 3961 9781 3995
rect 9815 3992 9827 3995
rect 11146 3992 11152 4004
rect 9815 3964 11152 3992
rect 9815 3961 9827 3964
rect 9769 3955 9827 3961
rect 11146 3952 11152 3964
rect 11204 3952 11210 4004
rect 1104 3834 10856 3856
rect 1104 3782 4246 3834
rect 4298 3782 4310 3834
rect 4362 3782 4374 3834
rect 4426 3782 4438 3834
rect 4490 3782 7510 3834
rect 7562 3782 7574 3834
rect 7626 3782 7638 3834
rect 7690 3782 7702 3834
rect 7754 3782 10856 3834
rect 1104 3760 10856 3782
rect 5169 3451 5227 3457
rect 5169 3417 5181 3451
rect 5215 3448 5227 3451
rect 7190 3448 7196 3460
rect 5215 3420 7196 3448
rect 5215 3417 5227 3420
rect 5169 3411 5227 3417
rect 7190 3408 7196 3420
rect 7248 3408 7254 3460
rect 1578 3340 1584 3392
rect 1636 3380 1642 3392
rect 2685 3383 2743 3389
rect 2685 3380 2697 3383
rect 1636 3352 2697 3380
rect 1636 3340 1642 3352
rect 2685 3349 2697 3352
rect 2731 3349 2743 3383
rect 2685 3343 2743 3349
rect 6733 3383 6791 3389
rect 6733 3349 6745 3383
rect 6779 3380 6791 3383
rect 7374 3380 7380 3392
rect 6779 3352 7380 3380
rect 6779 3349 6791 3352
rect 6733 3343 6791 3349
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 8205 3383 8263 3389
rect 8205 3349 8217 3383
rect 8251 3380 8263 3383
rect 8478 3380 8484 3392
rect 8251 3352 8484 3380
rect 8251 3349 8263 3352
rect 8205 3343 8263 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 1104 3290 10856 3312
rect 1104 3238 2614 3290
rect 2666 3238 2678 3290
rect 2730 3238 2742 3290
rect 2794 3238 2806 3290
rect 2858 3238 5878 3290
rect 5930 3238 5942 3290
rect 5994 3238 6006 3290
rect 6058 3238 6070 3290
rect 6122 3238 9142 3290
rect 9194 3238 9206 3290
rect 9258 3238 9270 3290
rect 9322 3238 9334 3290
rect 9386 3238 10856 3290
rect 1104 3216 10856 3238
rect 7374 2972 7380 2984
rect 7335 2944 7380 2972
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 8478 2972 8484 2984
rect 8439 2944 8484 2972
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8662 2932 8668 2984
rect 8720 2972 8726 2984
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 8720 2944 9597 2972
rect 8720 2932 8726 2944
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 7193 2907 7251 2913
rect 7193 2904 7205 2907
rect 6788 2876 7205 2904
rect 6788 2864 6794 2876
rect 7193 2873 7205 2876
rect 7239 2873 7251 2907
rect 7193 2867 7251 2873
rect 8202 2864 8208 2916
rect 8260 2904 8266 2916
rect 8297 2907 8355 2913
rect 8297 2904 8309 2907
rect 8260 2876 8309 2904
rect 8260 2864 8266 2876
rect 8297 2873 8309 2876
rect 8343 2873 8355 2907
rect 8297 2867 8355 2873
rect 9674 2836 9680 2848
rect 9635 2808 9680 2836
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 1104 2746 10856 2768
rect 1104 2694 4246 2746
rect 4298 2694 4310 2746
rect 4362 2694 4374 2746
rect 4426 2694 4438 2746
rect 4490 2694 7510 2746
rect 7562 2694 7574 2746
rect 7626 2694 7638 2746
rect 7690 2694 7702 2746
rect 7754 2694 10856 2746
rect 1104 2672 10856 2694
rect 1578 2564 1584 2576
rect 1539 2536 1584 2564
rect 1578 2524 1584 2536
rect 1636 2524 1642 2576
rect 2498 2524 2504 2576
rect 2556 2564 2562 2576
rect 2685 2567 2743 2573
rect 2685 2564 2697 2567
rect 2556 2536 2697 2564
rect 2556 2524 2562 2536
rect 2685 2533 2697 2536
rect 2731 2533 2743 2567
rect 4798 2564 4804 2576
rect 4759 2536 4804 2564
rect 2685 2527 2743 2533
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 7190 2524 7196 2576
rect 7248 2564 7254 2576
rect 7469 2567 7527 2573
rect 7469 2564 7481 2567
rect 7248 2536 7481 2564
rect 7248 2524 7254 2536
rect 7469 2533 7481 2536
rect 7515 2533 7527 2567
rect 7469 2527 7527 2533
rect 750 2320 756 2372
rect 808 2360 814 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 808 2332 1409 2360
rect 808 2320 814 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 2222 2320 2228 2372
rect 2280 2360 2286 2372
rect 2501 2363 2559 2369
rect 2501 2360 2513 2363
rect 2280 2332 2513 2360
rect 2280 2320 2286 2332
rect 2501 2329 2513 2332
rect 2547 2329 2559 2363
rect 2501 2323 2559 2329
rect 3694 2320 3700 2372
rect 3752 2360 3758 2372
rect 4617 2363 4675 2369
rect 4617 2360 4629 2363
rect 3752 2332 4629 2360
rect 3752 2320 3758 2332
rect 4617 2329 4629 2332
rect 4663 2329 4675 2363
rect 4617 2323 4675 2329
rect 5166 2320 5172 2372
rect 5224 2360 5230 2372
rect 7285 2363 7343 2369
rect 7285 2360 7297 2363
rect 5224 2332 7297 2360
rect 5224 2320 5230 2332
rect 7285 2329 7297 2332
rect 7331 2329 7343 2363
rect 7285 2323 7343 2329
rect 1104 2202 10856 2224
rect 1104 2150 2614 2202
rect 2666 2150 2678 2202
rect 2730 2150 2742 2202
rect 2794 2150 2806 2202
rect 2858 2150 5878 2202
rect 5930 2150 5942 2202
rect 5994 2150 6006 2202
rect 6058 2150 6070 2202
rect 6122 2150 9142 2202
rect 9194 2150 9206 2202
rect 9258 2150 9270 2202
rect 9322 2150 9334 2202
rect 9386 2150 10856 2202
rect 1104 2128 10856 2150
<< via1 >>
rect 4246 11398 4298 11450
rect 4310 11398 4362 11450
rect 4374 11398 4426 11450
rect 4438 11398 4490 11450
rect 7510 11398 7562 11450
rect 7574 11398 7626 11450
rect 7638 11398 7690 11450
rect 7702 11398 7754 11450
rect 2614 10854 2666 10906
rect 2678 10854 2730 10906
rect 2742 10854 2794 10906
rect 2806 10854 2858 10906
rect 5878 10854 5930 10906
rect 5942 10854 5994 10906
rect 6006 10854 6058 10906
rect 6070 10854 6122 10906
rect 9142 10854 9194 10906
rect 9206 10854 9258 10906
rect 9270 10854 9322 10906
rect 9334 10854 9386 10906
rect 4246 10310 4298 10362
rect 4310 10310 4362 10362
rect 4374 10310 4426 10362
rect 4438 10310 4490 10362
rect 7510 10310 7562 10362
rect 7574 10310 7626 10362
rect 7638 10310 7690 10362
rect 7702 10310 7754 10362
rect 2614 9766 2666 9818
rect 2678 9766 2730 9818
rect 2742 9766 2794 9818
rect 2806 9766 2858 9818
rect 5878 9766 5930 9818
rect 5942 9766 5994 9818
rect 6006 9766 6058 9818
rect 6070 9766 6122 9818
rect 9142 9766 9194 9818
rect 9206 9766 9258 9818
rect 9270 9766 9322 9818
rect 9334 9766 9386 9818
rect 4246 9222 4298 9274
rect 4310 9222 4362 9274
rect 4374 9222 4426 9274
rect 4438 9222 4490 9274
rect 7510 9222 7562 9274
rect 7574 9222 7626 9274
rect 7638 9222 7690 9274
rect 7702 9222 7754 9274
rect 2614 8678 2666 8730
rect 2678 8678 2730 8730
rect 2742 8678 2794 8730
rect 2806 8678 2858 8730
rect 5878 8678 5930 8730
rect 5942 8678 5994 8730
rect 6006 8678 6058 8730
rect 6070 8678 6122 8730
rect 9142 8678 9194 8730
rect 9206 8678 9258 8730
rect 9270 8678 9322 8730
rect 9334 8678 9386 8730
rect 4246 8134 4298 8186
rect 4310 8134 4362 8186
rect 4374 8134 4426 8186
rect 4438 8134 4490 8186
rect 7510 8134 7562 8186
rect 7574 8134 7626 8186
rect 7638 8134 7690 8186
rect 7702 8134 7754 8186
rect 2614 7590 2666 7642
rect 2678 7590 2730 7642
rect 2742 7590 2794 7642
rect 2806 7590 2858 7642
rect 5878 7590 5930 7642
rect 5942 7590 5994 7642
rect 6006 7590 6058 7642
rect 6070 7590 6122 7642
rect 9142 7590 9194 7642
rect 9206 7590 9258 7642
rect 9270 7590 9322 7642
rect 9334 7590 9386 7642
rect 4246 7046 4298 7098
rect 4310 7046 4362 7098
rect 4374 7046 4426 7098
rect 4438 7046 4490 7098
rect 7510 7046 7562 7098
rect 7574 7046 7626 7098
rect 7638 7046 7690 7098
rect 7702 7046 7754 7098
rect 2614 6502 2666 6554
rect 2678 6502 2730 6554
rect 2742 6502 2794 6554
rect 2806 6502 2858 6554
rect 5878 6502 5930 6554
rect 5942 6502 5994 6554
rect 6006 6502 6058 6554
rect 6070 6502 6122 6554
rect 9142 6502 9194 6554
rect 9206 6502 9258 6554
rect 9270 6502 9322 6554
rect 9334 6502 9386 6554
rect 4246 5958 4298 6010
rect 4310 5958 4362 6010
rect 4374 5958 4426 6010
rect 4438 5958 4490 6010
rect 7510 5958 7562 6010
rect 7574 5958 7626 6010
rect 7638 5958 7690 6010
rect 7702 5958 7754 6010
rect 2614 5414 2666 5466
rect 2678 5414 2730 5466
rect 2742 5414 2794 5466
rect 2806 5414 2858 5466
rect 5878 5414 5930 5466
rect 5942 5414 5994 5466
rect 6006 5414 6058 5466
rect 6070 5414 6122 5466
rect 9142 5414 9194 5466
rect 9206 5414 9258 5466
rect 9270 5414 9322 5466
rect 9334 5414 9386 5466
rect 9588 5108 9640 5160
rect 4246 4870 4298 4922
rect 4310 4870 4362 4922
rect 4374 4870 4426 4922
rect 4438 4870 4490 4922
rect 7510 4870 7562 4922
rect 7574 4870 7626 4922
rect 7638 4870 7690 4922
rect 7702 4870 7754 4922
rect 2614 4326 2666 4378
rect 2678 4326 2730 4378
rect 2742 4326 2794 4378
rect 2806 4326 2858 4378
rect 5878 4326 5930 4378
rect 5942 4326 5994 4378
rect 6006 4326 6058 4378
rect 6070 4326 6122 4378
rect 9142 4326 9194 4378
rect 9206 4326 9258 4378
rect 9270 4326 9322 4378
rect 9334 4326 9386 4378
rect 2504 4156 2556 4208
rect 4804 4156 4856 4208
rect 8668 4063 8720 4072
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 11152 3952 11204 4004
rect 4246 3782 4298 3834
rect 4310 3782 4362 3834
rect 4374 3782 4426 3834
rect 4438 3782 4490 3834
rect 7510 3782 7562 3834
rect 7574 3782 7626 3834
rect 7638 3782 7690 3834
rect 7702 3782 7754 3834
rect 7196 3408 7248 3460
rect 1584 3340 1636 3392
rect 7380 3340 7432 3392
rect 8484 3340 8536 3392
rect 2614 3238 2666 3290
rect 2678 3238 2730 3290
rect 2742 3238 2794 3290
rect 2806 3238 2858 3290
rect 5878 3238 5930 3290
rect 5942 3238 5994 3290
rect 6006 3238 6058 3290
rect 6070 3238 6122 3290
rect 9142 3238 9194 3290
rect 9206 3238 9258 3290
rect 9270 3238 9322 3290
rect 9334 3238 9386 3290
rect 7380 2975 7432 2984
rect 7380 2941 7389 2975
rect 7389 2941 7423 2975
rect 7423 2941 7432 2975
rect 7380 2932 7432 2941
rect 8484 2975 8536 2984
rect 8484 2941 8493 2975
rect 8493 2941 8527 2975
rect 8527 2941 8536 2975
rect 8484 2932 8536 2941
rect 8668 2932 8720 2984
rect 6736 2864 6788 2916
rect 8208 2864 8260 2916
rect 9680 2839 9732 2848
rect 9680 2805 9689 2839
rect 9689 2805 9723 2839
rect 9723 2805 9732 2839
rect 9680 2796 9732 2805
rect 4246 2694 4298 2746
rect 4310 2694 4362 2746
rect 4374 2694 4426 2746
rect 4438 2694 4490 2746
rect 7510 2694 7562 2746
rect 7574 2694 7626 2746
rect 7638 2694 7690 2746
rect 7702 2694 7754 2746
rect 1584 2567 1636 2576
rect 1584 2533 1593 2567
rect 1593 2533 1627 2567
rect 1627 2533 1636 2567
rect 1584 2524 1636 2533
rect 2504 2524 2556 2576
rect 4804 2567 4856 2576
rect 4804 2533 4813 2567
rect 4813 2533 4847 2567
rect 4847 2533 4856 2567
rect 4804 2524 4856 2533
rect 7196 2524 7248 2576
rect 756 2320 808 2372
rect 2228 2320 2280 2372
rect 3700 2320 3752 2372
rect 5172 2320 5224 2372
rect 2614 2150 2666 2202
rect 2678 2150 2730 2202
rect 2742 2150 2794 2202
rect 2806 2150 2858 2202
rect 5878 2150 5930 2202
rect 5942 2150 5994 2202
rect 6006 2150 6058 2202
rect 6070 2150 6122 2202
rect 9142 2150 9194 2202
rect 9206 2150 9258 2202
rect 9270 2150 9322 2202
rect 9334 2150 9386 2202
<< metal2 >>
rect 4220 11452 4516 11472
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4298 11398 4300 11450
rect 4362 11398 4374 11450
rect 4436 11398 4438 11450
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4220 11376 4516 11396
rect 7484 11452 7780 11472
rect 7540 11450 7564 11452
rect 7620 11450 7644 11452
rect 7700 11450 7724 11452
rect 7562 11398 7564 11450
rect 7626 11398 7638 11450
rect 7700 11398 7702 11450
rect 7540 11396 7564 11398
rect 7620 11396 7644 11398
rect 7700 11396 7724 11398
rect 7484 11376 7780 11396
rect 2588 10908 2884 10928
rect 2644 10906 2668 10908
rect 2724 10906 2748 10908
rect 2804 10906 2828 10908
rect 2666 10854 2668 10906
rect 2730 10854 2742 10906
rect 2804 10854 2806 10906
rect 2644 10852 2668 10854
rect 2724 10852 2748 10854
rect 2804 10852 2828 10854
rect 2588 10832 2884 10852
rect 5852 10908 6148 10928
rect 5908 10906 5932 10908
rect 5988 10906 6012 10908
rect 6068 10906 6092 10908
rect 5930 10854 5932 10906
rect 5994 10854 6006 10906
rect 6068 10854 6070 10906
rect 5908 10852 5932 10854
rect 5988 10852 6012 10854
rect 6068 10852 6092 10854
rect 5852 10832 6148 10852
rect 9116 10908 9412 10928
rect 9172 10906 9196 10908
rect 9252 10906 9276 10908
rect 9332 10906 9356 10908
rect 9194 10854 9196 10906
rect 9258 10854 9270 10906
rect 9332 10854 9334 10906
rect 9172 10852 9196 10854
rect 9252 10852 9276 10854
rect 9332 10852 9356 10854
rect 9116 10832 9412 10852
rect 4220 10364 4516 10384
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4298 10310 4300 10362
rect 4362 10310 4374 10362
rect 4436 10310 4438 10362
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4220 10288 4516 10308
rect 7484 10364 7780 10384
rect 7540 10362 7564 10364
rect 7620 10362 7644 10364
rect 7700 10362 7724 10364
rect 7562 10310 7564 10362
rect 7626 10310 7638 10362
rect 7700 10310 7702 10362
rect 7540 10308 7564 10310
rect 7620 10308 7644 10310
rect 7700 10308 7724 10310
rect 7484 10288 7780 10308
rect 2588 9820 2884 9840
rect 2644 9818 2668 9820
rect 2724 9818 2748 9820
rect 2804 9818 2828 9820
rect 2666 9766 2668 9818
rect 2730 9766 2742 9818
rect 2804 9766 2806 9818
rect 2644 9764 2668 9766
rect 2724 9764 2748 9766
rect 2804 9764 2828 9766
rect 2588 9744 2884 9764
rect 5852 9820 6148 9840
rect 5908 9818 5932 9820
rect 5988 9818 6012 9820
rect 6068 9818 6092 9820
rect 5930 9766 5932 9818
rect 5994 9766 6006 9818
rect 6068 9766 6070 9818
rect 5908 9764 5932 9766
rect 5988 9764 6012 9766
rect 6068 9764 6092 9766
rect 5852 9744 6148 9764
rect 9116 9820 9412 9840
rect 9172 9818 9196 9820
rect 9252 9818 9276 9820
rect 9332 9818 9356 9820
rect 9194 9766 9196 9818
rect 9258 9766 9270 9818
rect 9332 9766 9334 9818
rect 9172 9764 9196 9766
rect 9252 9764 9276 9766
rect 9332 9764 9356 9766
rect 9116 9744 9412 9764
rect 4220 9276 4516 9296
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4298 9222 4300 9274
rect 4362 9222 4374 9274
rect 4436 9222 4438 9274
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4220 9200 4516 9220
rect 7484 9276 7780 9296
rect 7540 9274 7564 9276
rect 7620 9274 7644 9276
rect 7700 9274 7724 9276
rect 7562 9222 7564 9274
rect 7626 9222 7638 9274
rect 7700 9222 7702 9274
rect 7540 9220 7564 9222
rect 7620 9220 7644 9222
rect 7700 9220 7724 9222
rect 7484 9200 7780 9220
rect 2588 8732 2884 8752
rect 2644 8730 2668 8732
rect 2724 8730 2748 8732
rect 2804 8730 2828 8732
rect 2666 8678 2668 8730
rect 2730 8678 2742 8730
rect 2804 8678 2806 8730
rect 2644 8676 2668 8678
rect 2724 8676 2748 8678
rect 2804 8676 2828 8678
rect 2588 8656 2884 8676
rect 5852 8732 6148 8752
rect 5908 8730 5932 8732
rect 5988 8730 6012 8732
rect 6068 8730 6092 8732
rect 5930 8678 5932 8730
rect 5994 8678 6006 8730
rect 6068 8678 6070 8730
rect 5908 8676 5932 8678
rect 5988 8676 6012 8678
rect 6068 8676 6092 8678
rect 5852 8656 6148 8676
rect 9116 8732 9412 8752
rect 9172 8730 9196 8732
rect 9252 8730 9276 8732
rect 9332 8730 9356 8732
rect 9194 8678 9196 8730
rect 9258 8678 9270 8730
rect 9332 8678 9334 8730
rect 9172 8676 9196 8678
rect 9252 8676 9276 8678
rect 9332 8676 9356 8678
rect 9116 8656 9412 8676
rect 4220 8188 4516 8208
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4298 8134 4300 8186
rect 4362 8134 4374 8186
rect 4436 8134 4438 8186
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4220 8112 4516 8132
rect 7484 8188 7780 8208
rect 7540 8186 7564 8188
rect 7620 8186 7644 8188
rect 7700 8186 7724 8188
rect 7562 8134 7564 8186
rect 7626 8134 7638 8186
rect 7700 8134 7702 8186
rect 7540 8132 7564 8134
rect 7620 8132 7644 8134
rect 7700 8132 7724 8134
rect 7484 8112 7780 8132
rect 2588 7644 2884 7664
rect 2644 7642 2668 7644
rect 2724 7642 2748 7644
rect 2804 7642 2828 7644
rect 2666 7590 2668 7642
rect 2730 7590 2742 7642
rect 2804 7590 2806 7642
rect 2644 7588 2668 7590
rect 2724 7588 2748 7590
rect 2804 7588 2828 7590
rect 2588 7568 2884 7588
rect 5852 7644 6148 7664
rect 5908 7642 5932 7644
rect 5988 7642 6012 7644
rect 6068 7642 6092 7644
rect 5930 7590 5932 7642
rect 5994 7590 6006 7642
rect 6068 7590 6070 7642
rect 5908 7588 5932 7590
rect 5988 7588 6012 7590
rect 6068 7588 6092 7590
rect 5852 7568 6148 7588
rect 9116 7644 9412 7664
rect 9172 7642 9196 7644
rect 9252 7642 9276 7644
rect 9332 7642 9356 7644
rect 9194 7590 9196 7642
rect 9258 7590 9270 7642
rect 9332 7590 9334 7642
rect 9172 7588 9196 7590
rect 9252 7588 9276 7590
rect 9332 7588 9356 7590
rect 9116 7568 9412 7588
rect 4220 7100 4516 7120
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4298 7046 4300 7098
rect 4362 7046 4374 7098
rect 4436 7046 4438 7098
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4220 7024 4516 7044
rect 7484 7100 7780 7120
rect 7540 7098 7564 7100
rect 7620 7098 7644 7100
rect 7700 7098 7724 7100
rect 7562 7046 7564 7098
rect 7626 7046 7638 7098
rect 7700 7046 7702 7098
rect 7540 7044 7564 7046
rect 7620 7044 7644 7046
rect 7700 7044 7724 7046
rect 7484 7024 7780 7044
rect 2588 6556 2884 6576
rect 2644 6554 2668 6556
rect 2724 6554 2748 6556
rect 2804 6554 2828 6556
rect 2666 6502 2668 6554
rect 2730 6502 2742 6554
rect 2804 6502 2806 6554
rect 2644 6500 2668 6502
rect 2724 6500 2748 6502
rect 2804 6500 2828 6502
rect 2588 6480 2884 6500
rect 5852 6556 6148 6576
rect 5908 6554 5932 6556
rect 5988 6554 6012 6556
rect 6068 6554 6092 6556
rect 5930 6502 5932 6554
rect 5994 6502 6006 6554
rect 6068 6502 6070 6554
rect 5908 6500 5932 6502
rect 5988 6500 6012 6502
rect 6068 6500 6092 6502
rect 5852 6480 6148 6500
rect 9116 6556 9412 6576
rect 9172 6554 9196 6556
rect 9252 6554 9276 6556
rect 9332 6554 9356 6556
rect 9194 6502 9196 6554
rect 9258 6502 9270 6554
rect 9332 6502 9334 6554
rect 9172 6500 9196 6502
rect 9252 6500 9276 6502
rect 9332 6500 9356 6502
rect 9116 6480 9412 6500
rect 4220 6012 4516 6032
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4298 5958 4300 6010
rect 4362 5958 4374 6010
rect 4436 5958 4438 6010
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4220 5936 4516 5956
rect 7484 6012 7780 6032
rect 7540 6010 7564 6012
rect 7620 6010 7644 6012
rect 7700 6010 7724 6012
rect 7562 5958 7564 6010
rect 7626 5958 7638 6010
rect 7700 5958 7702 6010
rect 7540 5956 7564 5958
rect 7620 5956 7644 5958
rect 7700 5956 7724 5958
rect 7484 5936 7780 5956
rect 2588 5468 2884 5488
rect 2644 5466 2668 5468
rect 2724 5466 2748 5468
rect 2804 5466 2828 5468
rect 2666 5414 2668 5466
rect 2730 5414 2742 5466
rect 2804 5414 2806 5466
rect 2644 5412 2668 5414
rect 2724 5412 2748 5414
rect 2804 5412 2828 5414
rect 2588 5392 2884 5412
rect 5852 5468 6148 5488
rect 5908 5466 5932 5468
rect 5988 5466 6012 5468
rect 6068 5466 6092 5468
rect 5930 5414 5932 5466
rect 5994 5414 6006 5466
rect 6068 5414 6070 5466
rect 5908 5412 5932 5414
rect 5988 5412 6012 5414
rect 6068 5412 6092 5414
rect 5852 5392 6148 5412
rect 9116 5468 9412 5488
rect 9172 5466 9196 5468
rect 9252 5466 9276 5468
rect 9332 5466 9356 5468
rect 9194 5414 9196 5466
rect 9258 5414 9270 5466
rect 9332 5414 9334 5466
rect 9172 5412 9196 5414
rect 9252 5412 9276 5414
rect 9332 5412 9356 5414
rect 9116 5392 9412 5412
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 4220 4924 4516 4944
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4298 4870 4300 4922
rect 4362 4870 4374 4922
rect 4436 4870 4438 4922
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4220 4848 4516 4868
rect 7484 4924 7780 4944
rect 7540 4922 7564 4924
rect 7620 4922 7644 4924
rect 7700 4922 7724 4924
rect 7562 4870 7564 4922
rect 7626 4870 7638 4922
rect 7700 4870 7702 4922
rect 7540 4868 7564 4870
rect 7620 4868 7644 4870
rect 7700 4868 7724 4870
rect 7484 4848 7780 4868
rect 2588 4380 2884 4400
rect 2644 4378 2668 4380
rect 2724 4378 2748 4380
rect 2804 4378 2828 4380
rect 2666 4326 2668 4378
rect 2730 4326 2742 4378
rect 2804 4326 2806 4378
rect 2644 4324 2668 4326
rect 2724 4324 2748 4326
rect 2804 4324 2828 4326
rect 2588 4304 2884 4324
rect 5852 4380 6148 4400
rect 5908 4378 5932 4380
rect 5988 4378 6012 4380
rect 6068 4378 6092 4380
rect 5930 4326 5932 4378
rect 5994 4326 6006 4378
rect 6068 4326 6070 4378
rect 5908 4324 5932 4326
rect 5988 4324 6012 4326
rect 6068 4324 6092 4326
rect 5852 4304 6148 4324
rect 9116 4380 9412 4400
rect 9172 4378 9196 4380
rect 9252 4378 9276 4380
rect 9332 4378 9356 4380
rect 9194 4326 9196 4378
rect 9258 4326 9270 4378
rect 9332 4326 9334 4378
rect 9172 4324 9196 4326
rect 9252 4324 9276 4326
rect 9332 4324 9356 4326
rect 9116 4304 9412 4324
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1596 2582 1624 3334
rect 2516 2582 2544 4150
rect 4220 3836 4516 3856
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4298 3782 4300 3834
rect 4362 3782 4374 3834
rect 4436 3782 4438 3834
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4220 3760 4516 3780
rect 2588 3292 2884 3312
rect 2644 3290 2668 3292
rect 2724 3290 2748 3292
rect 2804 3290 2828 3292
rect 2666 3238 2668 3290
rect 2730 3238 2742 3290
rect 2804 3238 2806 3290
rect 2644 3236 2668 3238
rect 2724 3236 2748 3238
rect 2804 3236 2828 3238
rect 2588 3216 2884 3236
rect 4220 2748 4516 2768
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4298 2694 4300 2746
rect 4362 2694 4374 2746
rect 4436 2694 4438 2746
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4220 2672 4516 2692
rect 4816 2582 4844 4150
rect 9600 4078 9628 5102
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 7484 3836 7780 3856
rect 7540 3834 7564 3836
rect 7620 3834 7644 3836
rect 7700 3834 7724 3836
rect 7562 3782 7564 3834
rect 7626 3782 7638 3834
rect 7700 3782 7702 3834
rect 7540 3780 7564 3782
rect 7620 3780 7644 3782
rect 7700 3780 7724 3782
rect 7484 3760 7780 3780
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 5852 3292 6148 3312
rect 5908 3290 5932 3292
rect 5988 3290 6012 3292
rect 6068 3290 6092 3292
rect 5930 3238 5932 3290
rect 5994 3238 6006 3290
rect 6068 3238 6070 3290
rect 5908 3236 5932 3238
rect 5988 3236 6012 3238
rect 6068 3236 6092 3238
rect 5852 3216 6148 3236
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 1584 2576 1636 2582
rect 1584 2518 1636 2524
rect 2504 2576 2556 2582
rect 2504 2518 2556 2524
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 756 2372 808 2378
rect 756 2314 808 2320
rect 2228 2372 2280 2378
rect 2228 2314 2280 2320
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 768 800 796 2314
rect 2240 800 2268 2314
rect 2588 2204 2884 2224
rect 2644 2202 2668 2204
rect 2724 2202 2748 2204
rect 2804 2202 2828 2204
rect 2666 2150 2668 2202
rect 2730 2150 2742 2202
rect 2804 2150 2806 2202
rect 2644 2148 2668 2150
rect 2724 2148 2748 2150
rect 2804 2148 2828 2150
rect 2588 2128 2884 2148
rect 3712 800 3740 2314
rect 5184 800 5212 2314
rect 5852 2204 6148 2224
rect 5908 2202 5932 2204
rect 5988 2202 6012 2204
rect 6068 2202 6092 2204
rect 5930 2150 5932 2202
rect 5994 2150 6006 2202
rect 6068 2150 6070 2202
rect 5908 2148 5932 2150
rect 5988 2148 6012 2150
rect 6068 2148 6092 2150
rect 5852 2128 6148 2148
rect 6748 800 6776 2858
rect 7208 2582 7236 3402
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 7392 2990 7420 3334
rect 8496 2990 8524 3334
rect 8680 2990 8708 4014
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 9116 3292 9412 3312
rect 9172 3290 9196 3292
rect 9252 3290 9276 3292
rect 9332 3290 9356 3292
rect 9194 3238 9196 3290
rect 9258 3238 9270 3290
rect 9332 3238 9334 3290
rect 9172 3236 9196 3238
rect 9252 3236 9276 3238
rect 9332 3236 9356 3238
rect 9116 3216 9412 3236
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 7484 2748 7780 2768
rect 7540 2746 7564 2748
rect 7620 2746 7644 2748
rect 7700 2746 7724 2748
rect 7562 2694 7564 2746
rect 7626 2694 7638 2746
rect 7700 2694 7702 2746
rect 7540 2692 7564 2694
rect 7620 2692 7644 2694
rect 7700 2692 7724 2694
rect 7484 2672 7780 2692
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 8220 800 8248 2858
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9116 2204 9412 2224
rect 9172 2202 9196 2204
rect 9252 2202 9276 2204
rect 9332 2202 9356 2204
rect 9194 2150 9196 2202
rect 9258 2150 9270 2202
rect 9332 2150 9334 2202
rect 9172 2148 9196 2150
rect 9252 2148 9276 2150
rect 9332 2148 9356 2150
rect 9116 2128 9412 2148
rect 9692 800 9720 2790
rect 11164 800 11192 3946
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6734 0 6790 800
rect 8206 0 8262 800
rect 9678 0 9734 800
rect 11150 0 11206 800
<< via2 >>
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4246 11450
rect 4246 11398 4276 11450
rect 4300 11398 4310 11450
rect 4310 11398 4356 11450
rect 4380 11398 4426 11450
rect 4426 11398 4436 11450
rect 4460 11398 4490 11450
rect 4490 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 7484 11450 7540 11452
rect 7564 11450 7620 11452
rect 7644 11450 7700 11452
rect 7724 11450 7780 11452
rect 7484 11398 7510 11450
rect 7510 11398 7540 11450
rect 7564 11398 7574 11450
rect 7574 11398 7620 11450
rect 7644 11398 7690 11450
rect 7690 11398 7700 11450
rect 7724 11398 7754 11450
rect 7754 11398 7780 11450
rect 7484 11396 7540 11398
rect 7564 11396 7620 11398
rect 7644 11396 7700 11398
rect 7724 11396 7780 11398
rect 2588 10906 2644 10908
rect 2668 10906 2724 10908
rect 2748 10906 2804 10908
rect 2828 10906 2884 10908
rect 2588 10854 2614 10906
rect 2614 10854 2644 10906
rect 2668 10854 2678 10906
rect 2678 10854 2724 10906
rect 2748 10854 2794 10906
rect 2794 10854 2804 10906
rect 2828 10854 2858 10906
rect 2858 10854 2884 10906
rect 2588 10852 2644 10854
rect 2668 10852 2724 10854
rect 2748 10852 2804 10854
rect 2828 10852 2884 10854
rect 5852 10906 5908 10908
rect 5932 10906 5988 10908
rect 6012 10906 6068 10908
rect 6092 10906 6148 10908
rect 5852 10854 5878 10906
rect 5878 10854 5908 10906
rect 5932 10854 5942 10906
rect 5942 10854 5988 10906
rect 6012 10854 6058 10906
rect 6058 10854 6068 10906
rect 6092 10854 6122 10906
rect 6122 10854 6148 10906
rect 5852 10852 5908 10854
rect 5932 10852 5988 10854
rect 6012 10852 6068 10854
rect 6092 10852 6148 10854
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 9276 10906 9332 10908
rect 9356 10906 9412 10908
rect 9116 10854 9142 10906
rect 9142 10854 9172 10906
rect 9196 10854 9206 10906
rect 9206 10854 9252 10906
rect 9276 10854 9322 10906
rect 9322 10854 9332 10906
rect 9356 10854 9386 10906
rect 9386 10854 9412 10906
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 9276 10852 9332 10854
rect 9356 10852 9412 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4246 10362
rect 4246 10310 4276 10362
rect 4300 10310 4310 10362
rect 4310 10310 4356 10362
rect 4380 10310 4426 10362
rect 4426 10310 4436 10362
rect 4460 10310 4490 10362
rect 4490 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 7484 10362 7540 10364
rect 7564 10362 7620 10364
rect 7644 10362 7700 10364
rect 7724 10362 7780 10364
rect 7484 10310 7510 10362
rect 7510 10310 7540 10362
rect 7564 10310 7574 10362
rect 7574 10310 7620 10362
rect 7644 10310 7690 10362
rect 7690 10310 7700 10362
rect 7724 10310 7754 10362
rect 7754 10310 7780 10362
rect 7484 10308 7540 10310
rect 7564 10308 7620 10310
rect 7644 10308 7700 10310
rect 7724 10308 7780 10310
rect 2588 9818 2644 9820
rect 2668 9818 2724 9820
rect 2748 9818 2804 9820
rect 2828 9818 2884 9820
rect 2588 9766 2614 9818
rect 2614 9766 2644 9818
rect 2668 9766 2678 9818
rect 2678 9766 2724 9818
rect 2748 9766 2794 9818
rect 2794 9766 2804 9818
rect 2828 9766 2858 9818
rect 2858 9766 2884 9818
rect 2588 9764 2644 9766
rect 2668 9764 2724 9766
rect 2748 9764 2804 9766
rect 2828 9764 2884 9766
rect 5852 9818 5908 9820
rect 5932 9818 5988 9820
rect 6012 9818 6068 9820
rect 6092 9818 6148 9820
rect 5852 9766 5878 9818
rect 5878 9766 5908 9818
rect 5932 9766 5942 9818
rect 5942 9766 5988 9818
rect 6012 9766 6058 9818
rect 6058 9766 6068 9818
rect 6092 9766 6122 9818
rect 6122 9766 6148 9818
rect 5852 9764 5908 9766
rect 5932 9764 5988 9766
rect 6012 9764 6068 9766
rect 6092 9764 6148 9766
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 9276 9818 9332 9820
rect 9356 9818 9412 9820
rect 9116 9766 9142 9818
rect 9142 9766 9172 9818
rect 9196 9766 9206 9818
rect 9206 9766 9252 9818
rect 9276 9766 9322 9818
rect 9322 9766 9332 9818
rect 9356 9766 9386 9818
rect 9386 9766 9412 9818
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 9276 9764 9332 9766
rect 9356 9764 9412 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4246 9274
rect 4246 9222 4276 9274
rect 4300 9222 4310 9274
rect 4310 9222 4356 9274
rect 4380 9222 4426 9274
rect 4426 9222 4436 9274
rect 4460 9222 4490 9274
rect 4490 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 7484 9274 7540 9276
rect 7564 9274 7620 9276
rect 7644 9274 7700 9276
rect 7724 9274 7780 9276
rect 7484 9222 7510 9274
rect 7510 9222 7540 9274
rect 7564 9222 7574 9274
rect 7574 9222 7620 9274
rect 7644 9222 7690 9274
rect 7690 9222 7700 9274
rect 7724 9222 7754 9274
rect 7754 9222 7780 9274
rect 7484 9220 7540 9222
rect 7564 9220 7620 9222
rect 7644 9220 7700 9222
rect 7724 9220 7780 9222
rect 2588 8730 2644 8732
rect 2668 8730 2724 8732
rect 2748 8730 2804 8732
rect 2828 8730 2884 8732
rect 2588 8678 2614 8730
rect 2614 8678 2644 8730
rect 2668 8678 2678 8730
rect 2678 8678 2724 8730
rect 2748 8678 2794 8730
rect 2794 8678 2804 8730
rect 2828 8678 2858 8730
rect 2858 8678 2884 8730
rect 2588 8676 2644 8678
rect 2668 8676 2724 8678
rect 2748 8676 2804 8678
rect 2828 8676 2884 8678
rect 5852 8730 5908 8732
rect 5932 8730 5988 8732
rect 6012 8730 6068 8732
rect 6092 8730 6148 8732
rect 5852 8678 5878 8730
rect 5878 8678 5908 8730
rect 5932 8678 5942 8730
rect 5942 8678 5988 8730
rect 6012 8678 6058 8730
rect 6058 8678 6068 8730
rect 6092 8678 6122 8730
rect 6122 8678 6148 8730
rect 5852 8676 5908 8678
rect 5932 8676 5988 8678
rect 6012 8676 6068 8678
rect 6092 8676 6148 8678
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 9276 8730 9332 8732
rect 9356 8730 9412 8732
rect 9116 8678 9142 8730
rect 9142 8678 9172 8730
rect 9196 8678 9206 8730
rect 9206 8678 9252 8730
rect 9276 8678 9322 8730
rect 9322 8678 9332 8730
rect 9356 8678 9386 8730
rect 9386 8678 9412 8730
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 9276 8676 9332 8678
rect 9356 8676 9412 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4246 8186
rect 4246 8134 4276 8186
rect 4300 8134 4310 8186
rect 4310 8134 4356 8186
rect 4380 8134 4426 8186
rect 4426 8134 4436 8186
rect 4460 8134 4490 8186
rect 4490 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 7484 8186 7540 8188
rect 7564 8186 7620 8188
rect 7644 8186 7700 8188
rect 7724 8186 7780 8188
rect 7484 8134 7510 8186
rect 7510 8134 7540 8186
rect 7564 8134 7574 8186
rect 7574 8134 7620 8186
rect 7644 8134 7690 8186
rect 7690 8134 7700 8186
rect 7724 8134 7754 8186
rect 7754 8134 7780 8186
rect 7484 8132 7540 8134
rect 7564 8132 7620 8134
rect 7644 8132 7700 8134
rect 7724 8132 7780 8134
rect 2588 7642 2644 7644
rect 2668 7642 2724 7644
rect 2748 7642 2804 7644
rect 2828 7642 2884 7644
rect 2588 7590 2614 7642
rect 2614 7590 2644 7642
rect 2668 7590 2678 7642
rect 2678 7590 2724 7642
rect 2748 7590 2794 7642
rect 2794 7590 2804 7642
rect 2828 7590 2858 7642
rect 2858 7590 2884 7642
rect 2588 7588 2644 7590
rect 2668 7588 2724 7590
rect 2748 7588 2804 7590
rect 2828 7588 2884 7590
rect 5852 7642 5908 7644
rect 5932 7642 5988 7644
rect 6012 7642 6068 7644
rect 6092 7642 6148 7644
rect 5852 7590 5878 7642
rect 5878 7590 5908 7642
rect 5932 7590 5942 7642
rect 5942 7590 5988 7642
rect 6012 7590 6058 7642
rect 6058 7590 6068 7642
rect 6092 7590 6122 7642
rect 6122 7590 6148 7642
rect 5852 7588 5908 7590
rect 5932 7588 5988 7590
rect 6012 7588 6068 7590
rect 6092 7588 6148 7590
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 9276 7642 9332 7644
rect 9356 7642 9412 7644
rect 9116 7590 9142 7642
rect 9142 7590 9172 7642
rect 9196 7590 9206 7642
rect 9206 7590 9252 7642
rect 9276 7590 9322 7642
rect 9322 7590 9332 7642
rect 9356 7590 9386 7642
rect 9386 7590 9412 7642
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 9276 7588 9332 7590
rect 9356 7588 9412 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4246 7098
rect 4246 7046 4276 7098
rect 4300 7046 4310 7098
rect 4310 7046 4356 7098
rect 4380 7046 4426 7098
rect 4426 7046 4436 7098
rect 4460 7046 4490 7098
rect 4490 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 7484 7098 7540 7100
rect 7564 7098 7620 7100
rect 7644 7098 7700 7100
rect 7724 7098 7780 7100
rect 7484 7046 7510 7098
rect 7510 7046 7540 7098
rect 7564 7046 7574 7098
rect 7574 7046 7620 7098
rect 7644 7046 7690 7098
rect 7690 7046 7700 7098
rect 7724 7046 7754 7098
rect 7754 7046 7780 7098
rect 7484 7044 7540 7046
rect 7564 7044 7620 7046
rect 7644 7044 7700 7046
rect 7724 7044 7780 7046
rect 2588 6554 2644 6556
rect 2668 6554 2724 6556
rect 2748 6554 2804 6556
rect 2828 6554 2884 6556
rect 2588 6502 2614 6554
rect 2614 6502 2644 6554
rect 2668 6502 2678 6554
rect 2678 6502 2724 6554
rect 2748 6502 2794 6554
rect 2794 6502 2804 6554
rect 2828 6502 2858 6554
rect 2858 6502 2884 6554
rect 2588 6500 2644 6502
rect 2668 6500 2724 6502
rect 2748 6500 2804 6502
rect 2828 6500 2884 6502
rect 5852 6554 5908 6556
rect 5932 6554 5988 6556
rect 6012 6554 6068 6556
rect 6092 6554 6148 6556
rect 5852 6502 5878 6554
rect 5878 6502 5908 6554
rect 5932 6502 5942 6554
rect 5942 6502 5988 6554
rect 6012 6502 6058 6554
rect 6058 6502 6068 6554
rect 6092 6502 6122 6554
rect 6122 6502 6148 6554
rect 5852 6500 5908 6502
rect 5932 6500 5988 6502
rect 6012 6500 6068 6502
rect 6092 6500 6148 6502
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 9276 6554 9332 6556
rect 9356 6554 9412 6556
rect 9116 6502 9142 6554
rect 9142 6502 9172 6554
rect 9196 6502 9206 6554
rect 9206 6502 9252 6554
rect 9276 6502 9322 6554
rect 9322 6502 9332 6554
rect 9356 6502 9386 6554
rect 9386 6502 9412 6554
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 9276 6500 9332 6502
rect 9356 6500 9412 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4246 6010
rect 4246 5958 4276 6010
rect 4300 5958 4310 6010
rect 4310 5958 4356 6010
rect 4380 5958 4426 6010
rect 4426 5958 4436 6010
rect 4460 5958 4490 6010
rect 4490 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 7484 6010 7540 6012
rect 7564 6010 7620 6012
rect 7644 6010 7700 6012
rect 7724 6010 7780 6012
rect 7484 5958 7510 6010
rect 7510 5958 7540 6010
rect 7564 5958 7574 6010
rect 7574 5958 7620 6010
rect 7644 5958 7690 6010
rect 7690 5958 7700 6010
rect 7724 5958 7754 6010
rect 7754 5958 7780 6010
rect 7484 5956 7540 5958
rect 7564 5956 7620 5958
rect 7644 5956 7700 5958
rect 7724 5956 7780 5958
rect 2588 5466 2644 5468
rect 2668 5466 2724 5468
rect 2748 5466 2804 5468
rect 2828 5466 2884 5468
rect 2588 5414 2614 5466
rect 2614 5414 2644 5466
rect 2668 5414 2678 5466
rect 2678 5414 2724 5466
rect 2748 5414 2794 5466
rect 2794 5414 2804 5466
rect 2828 5414 2858 5466
rect 2858 5414 2884 5466
rect 2588 5412 2644 5414
rect 2668 5412 2724 5414
rect 2748 5412 2804 5414
rect 2828 5412 2884 5414
rect 5852 5466 5908 5468
rect 5932 5466 5988 5468
rect 6012 5466 6068 5468
rect 6092 5466 6148 5468
rect 5852 5414 5878 5466
rect 5878 5414 5908 5466
rect 5932 5414 5942 5466
rect 5942 5414 5988 5466
rect 6012 5414 6058 5466
rect 6058 5414 6068 5466
rect 6092 5414 6122 5466
rect 6122 5414 6148 5466
rect 5852 5412 5908 5414
rect 5932 5412 5988 5414
rect 6012 5412 6068 5414
rect 6092 5412 6148 5414
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 9276 5466 9332 5468
rect 9356 5466 9412 5468
rect 9116 5414 9142 5466
rect 9142 5414 9172 5466
rect 9196 5414 9206 5466
rect 9206 5414 9252 5466
rect 9276 5414 9322 5466
rect 9322 5414 9332 5466
rect 9356 5414 9386 5466
rect 9386 5414 9412 5466
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 9276 5412 9332 5414
rect 9356 5412 9412 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4246 4922
rect 4246 4870 4276 4922
rect 4300 4870 4310 4922
rect 4310 4870 4356 4922
rect 4380 4870 4426 4922
rect 4426 4870 4436 4922
rect 4460 4870 4490 4922
rect 4490 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 7484 4922 7540 4924
rect 7564 4922 7620 4924
rect 7644 4922 7700 4924
rect 7724 4922 7780 4924
rect 7484 4870 7510 4922
rect 7510 4870 7540 4922
rect 7564 4870 7574 4922
rect 7574 4870 7620 4922
rect 7644 4870 7690 4922
rect 7690 4870 7700 4922
rect 7724 4870 7754 4922
rect 7754 4870 7780 4922
rect 7484 4868 7540 4870
rect 7564 4868 7620 4870
rect 7644 4868 7700 4870
rect 7724 4868 7780 4870
rect 2588 4378 2644 4380
rect 2668 4378 2724 4380
rect 2748 4378 2804 4380
rect 2828 4378 2884 4380
rect 2588 4326 2614 4378
rect 2614 4326 2644 4378
rect 2668 4326 2678 4378
rect 2678 4326 2724 4378
rect 2748 4326 2794 4378
rect 2794 4326 2804 4378
rect 2828 4326 2858 4378
rect 2858 4326 2884 4378
rect 2588 4324 2644 4326
rect 2668 4324 2724 4326
rect 2748 4324 2804 4326
rect 2828 4324 2884 4326
rect 5852 4378 5908 4380
rect 5932 4378 5988 4380
rect 6012 4378 6068 4380
rect 6092 4378 6148 4380
rect 5852 4326 5878 4378
rect 5878 4326 5908 4378
rect 5932 4326 5942 4378
rect 5942 4326 5988 4378
rect 6012 4326 6058 4378
rect 6058 4326 6068 4378
rect 6092 4326 6122 4378
rect 6122 4326 6148 4378
rect 5852 4324 5908 4326
rect 5932 4324 5988 4326
rect 6012 4324 6068 4326
rect 6092 4324 6148 4326
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 9276 4378 9332 4380
rect 9356 4378 9412 4380
rect 9116 4326 9142 4378
rect 9142 4326 9172 4378
rect 9196 4326 9206 4378
rect 9206 4326 9252 4378
rect 9276 4326 9322 4378
rect 9322 4326 9332 4378
rect 9356 4326 9386 4378
rect 9386 4326 9412 4378
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 9276 4324 9332 4326
rect 9356 4324 9412 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4246 3834
rect 4246 3782 4276 3834
rect 4300 3782 4310 3834
rect 4310 3782 4356 3834
rect 4380 3782 4426 3834
rect 4426 3782 4436 3834
rect 4460 3782 4490 3834
rect 4490 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 2588 3290 2644 3292
rect 2668 3290 2724 3292
rect 2748 3290 2804 3292
rect 2828 3290 2884 3292
rect 2588 3238 2614 3290
rect 2614 3238 2644 3290
rect 2668 3238 2678 3290
rect 2678 3238 2724 3290
rect 2748 3238 2794 3290
rect 2794 3238 2804 3290
rect 2828 3238 2858 3290
rect 2858 3238 2884 3290
rect 2588 3236 2644 3238
rect 2668 3236 2724 3238
rect 2748 3236 2804 3238
rect 2828 3236 2884 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4246 2746
rect 4246 2694 4276 2746
rect 4300 2694 4310 2746
rect 4310 2694 4356 2746
rect 4380 2694 4426 2746
rect 4426 2694 4436 2746
rect 4460 2694 4490 2746
rect 4490 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 7484 3834 7540 3836
rect 7564 3834 7620 3836
rect 7644 3834 7700 3836
rect 7724 3834 7780 3836
rect 7484 3782 7510 3834
rect 7510 3782 7540 3834
rect 7564 3782 7574 3834
rect 7574 3782 7620 3834
rect 7644 3782 7690 3834
rect 7690 3782 7700 3834
rect 7724 3782 7754 3834
rect 7754 3782 7780 3834
rect 7484 3780 7540 3782
rect 7564 3780 7620 3782
rect 7644 3780 7700 3782
rect 7724 3780 7780 3782
rect 5852 3290 5908 3292
rect 5932 3290 5988 3292
rect 6012 3290 6068 3292
rect 6092 3290 6148 3292
rect 5852 3238 5878 3290
rect 5878 3238 5908 3290
rect 5932 3238 5942 3290
rect 5942 3238 5988 3290
rect 6012 3238 6058 3290
rect 6058 3238 6068 3290
rect 6092 3238 6122 3290
rect 6122 3238 6148 3290
rect 5852 3236 5908 3238
rect 5932 3236 5988 3238
rect 6012 3236 6068 3238
rect 6092 3236 6148 3238
rect 2588 2202 2644 2204
rect 2668 2202 2724 2204
rect 2748 2202 2804 2204
rect 2828 2202 2884 2204
rect 2588 2150 2614 2202
rect 2614 2150 2644 2202
rect 2668 2150 2678 2202
rect 2678 2150 2724 2202
rect 2748 2150 2794 2202
rect 2794 2150 2804 2202
rect 2828 2150 2858 2202
rect 2858 2150 2884 2202
rect 2588 2148 2644 2150
rect 2668 2148 2724 2150
rect 2748 2148 2804 2150
rect 2828 2148 2884 2150
rect 5852 2202 5908 2204
rect 5932 2202 5988 2204
rect 6012 2202 6068 2204
rect 6092 2202 6148 2204
rect 5852 2150 5878 2202
rect 5878 2150 5908 2202
rect 5932 2150 5942 2202
rect 5942 2150 5988 2202
rect 6012 2150 6058 2202
rect 6058 2150 6068 2202
rect 6092 2150 6122 2202
rect 6122 2150 6148 2202
rect 5852 2148 5908 2150
rect 5932 2148 5988 2150
rect 6012 2148 6068 2150
rect 6092 2148 6148 2150
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 9276 3290 9332 3292
rect 9356 3290 9412 3292
rect 9116 3238 9142 3290
rect 9142 3238 9172 3290
rect 9196 3238 9206 3290
rect 9206 3238 9252 3290
rect 9276 3238 9322 3290
rect 9322 3238 9332 3290
rect 9356 3238 9386 3290
rect 9386 3238 9412 3290
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 9276 3236 9332 3238
rect 9356 3236 9412 3238
rect 7484 2746 7540 2748
rect 7564 2746 7620 2748
rect 7644 2746 7700 2748
rect 7724 2746 7780 2748
rect 7484 2694 7510 2746
rect 7510 2694 7540 2746
rect 7564 2694 7574 2746
rect 7574 2694 7620 2746
rect 7644 2694 7690 2746
rect 7690 2694 7700 2746
rect 7724 2694 7754 2746
rect 7754 2694 7780 2746
rect 7484 2692 7540 2694
rect 7564 2692 7620 2694
rect 7644 2692 7700 2694
rect 7724 2692 7780 2694
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 9276 2202 9332 2204
rect 9356 2202 9412 2204
rect 9116 2150 9142 2202
rect 9142 2150 9172 2202
rect 9196 2150 9206 2202
rect 9206 2150 9252 2202
rect 9276 2150 9322 2202
rect 9322 2150 9332 2202
rect 9356 2150 9386 2202
rect 9386 2150 9412 2202
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 9276 2148 9332 2150
rect 9356 2148 9412 2150
<< metal3 >>
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 7472 11456 7792 11457
rect 7472 11392 7480 11456
rect 7544 11392 7560 11456
rect 7624 11392 7640 11456
rect 7704 11392 7720 11456
rect 7784 11392 7792 11456
rect 7472 11391 7792 11392
rect 2576 10912 2896 10913
rect 2576 10848 2584 10912
rect 2648 10848 2664 10912
rect 2728 10848 2744 10912
rect 2808 10848 2824 10912
rect 2888 10848 2896 10912
rect 2576 10847 2896 10848
rect 5840 10912 6160 10913
rect 5840 10848 5848 10912
rect 5912 10848 5928 10912
rect 5992 10848 6008 10912
rect 6072 10848 6088 10912
rect 6152 10848 6160 10912
rect 5840 10847 6160 10848
rect 9104 10912 9424 10913
rect 9104 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9272 10912
rect 9336 10848 9352 10912
rect 9416 10848 9424 10912
rect 9104 10847 9424 10848
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 7472 10368 7792 10369
rect 7472 10304 7480 10368
rect 7544 10304 7560 10368
rect 7624 10304 7640 10368
rect 7704 10304 7720 10368
rect 7784 10304 7792 10368
rect 7472 10303 7792 10304
rect 2576 9824 2896 9825
rect 2576 9760 2584 9824
rect 2648 9760 2664 9824
rect 2728 9760 2744 9824
rect 2808 9760 2824 9824
rect 2888 9760 2896 9824
rect 2576 9759 2896 9760
rect 5840 9824 6160 9825
rect 5840 9760 5848 9824
rect 5912 9760 5928 9824
rect 5992 9760 6008 9824
rect 6072 9760 6088 9824
rect 6152 9760 6160 9824
rect 5840 9759 6160 9760
rect 9104 9824 9424 9825
rect 9104 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9272 9824
rect 9336 9760 9352 9824
rect 9416 9760 9424 9824
rect 9104 9759 9424 9760
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 7472 9280 7792 9281
rect 7472 9216 7480 9280
rect 7544 9216 7560 9280
rect 7624 9216 7640 9280
rect 7704 9216 7720 9280
rect 7784 9216 7792 9280
rect 7472 9215 7792 9216
rect 2576 8736 2896 8737
rect 2576 8672 2584 8736
rect 2648 8672 2664 8736
rect 2728 8672 2744 8736
rect 2808 8672 2824 8736
rect 2888 8672 2896 8736
rect 2576 8671 2896 8672
rect 5840 8736 6160 8737
rect 5840 8672 5848 8736
rect 5912 8672 5928 8736
rect 5992 8672 6008 8736
rect 6072 8672 6088 8736
rect 6152 8672 6160 8736
rect 5840 8671 6160 8672
rect 9104 8736 9424 8737
rect 9104 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9272 8736
rect 9336 8672 9352 8736
rect 9416 8672 9424 8736
rect 9104 8671 9424 8672
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 7472 8192 7792 8193
rect 7472 8128 7480 8192
rect 7544 8128 7560 8192
rect 7624 8128 7640 8192
rect 7704 8128 7720 8192
rect 7784 8128 7792 8192
rect 7472 8127 7792 8128
rect 2576 7648 2896 7649
rect 2576 7584 2584 7648
rect 2648 7584 2664 7648
rect 2728 7584 2744 7648
rect 2808 7584 2824 7648
rect 2888 7584 2896 7648
rect 2576 7583 2896 7584
rect 5840 7648 6160 7649
rect 5840 7584 5848 7648
rect 5912 7584 5928 7648
rect 5992 7584 6008 7648
rect 6072 7584 6088 7648
rect 6152 7584 6160 7648
rect 5840 7583 6160 7584
rect 9104 7648 9424 7649
rect 9104 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9272 7648
rect 9336 7584 9352 7648
rect 9416 7584 9424 7648
rect 9104 7583 9424 7584
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 7472 7104 7792 7105
rect 7472 7040 7480 7104
rect 7544 7040 7560 7104
rect 7624 7040 7640 7104
rect 7704 7040 7720 7104
rect 7784 7040 7792 7104
rect 7472 7039 7792 7040
rect 2576 6560 2896 6561
rect 2576 6496 2584 6560
rect 2648 6496 2664 6560
rect 2728 6496 2744 6560
rect 2808 6496 2824 6560
rect 2888 6496 2896 6560
rect 2576 6495 2896 6496
rect 5840 6560 6160 6561
rect 5840 6496 5848 6560
rect 5912 6496 5928 6560
rect 5992 6496 6008 6560
rect 6072 6496 6088 6560
rect 6152 6496 6160 6560
rect 5840 6495 6160 6496
rect 9104 6560 9424 6561
rect 9104 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9272 6560
rect 9336 6496 9352 6560
rect 9416 6496 9424 6560
rect 9104 6495 9424 6496
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 7472 6016 7792 6017
rect 7472 5952 7480 6016
rect 7544 5952 7560 6016
rect 7624 5952 7640 6016
rect 7704 5952 7720 6016
rect 7784 5952 7792 6016
rect 7472 5951 7792 5952
rect 2576 5472 2896 5473
rect 2576 5408 2584 5472
rect 2648 5408 2664 5472
rect 2728 5408 2744 5472
rect 2808 5408 2824 5472
rect 2888 5408 2896 5472
rect 2576 5407 2896 5408
rect 5840 5472 6160 5473
rect 5840 5408 5848 5472
rect 5912 5408 5928 5472
rect 5992 5408 6008 5472
rect 6072 5408 6088 5472
rect 6152 5408 6160 5472
rect 5840 5407 6160 5408
rect 9104 5472 9424 5473
rect 9104 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9272 5472
rect 9336 5408 9352 5472
rect 9416 5408 9424 5472
rect 9104 5407 9424 5408
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 7472 4928 7792 4929
rect 7472 4864 7480 4928
rect 7544 4864 7560 4928
rect 7624 4864 7640 4928
rect 7704 4864 7720 4928
rect 7784 4864 7792 4928
rect 7472 4863 7792 4864
rect 2576 4384 2896 4385
rect 2576 4320 2584 4384
rect 2648 4320 2664 4384
rect 2728 4320 2744 4384
rect 2808 4320 2824 4384
rect 2888 4320 2896 4384
rect 2576 4319 2896 4320
rect 5840 4384 6160 4385
rect 5840 4320 5848 4384
rect 5912 4320 5928 4384
rect 5992 4320 6008 4384
rect 6072 4320 6088 4384
rect 6152 4320 6160 4384
rect 5840 4319 6160 4320
rect 9104 4384 9424 4385
rect 9104 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9272 4384
rect 9336 4320 9352 4384
rect 9416 4320 9424 4384
rect 9104 4319 9424 4320
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 7472 3840 7792 3841
rect 7472 3776 7480 3840
rect 7544 3776 7560 3840
rect 7624 3776 7640 3840
rect 7704 3776 7720 3840
rect 7784 3776 7792 3840
rect 7472 3775 7792 3776
rect 2576 3296 2896 3297
rect 2576 3232 2584 3296
rect 2648 3232 2664 3296
rect 2728 3232 2744 3296
rect 2808 3232 2824 3296
rect 2888 3232 2896 3296
rect 2576 3231 2896 3232
rect 5840 3296 6160 3297
rect 5840 3232 5848 3296
rect 5912 3232 5928 3296
rect 5992 3232 6008 3296
rect 6072 3232 6088 3296
rect 6152 3232 6160 3296
rect 5840 3231 6160 3232
rect 9104 3296 9424 3297
rect 9104 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9272 3296
rect 9336 3232 9352 3296
rect 9416 3232 9424 3296
rect 9104 3231 9424 3232
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 7472 2752 7792 2753
rect 7472 2688 7480 2752
rect 7544 2688 7560 2752
rect 7624 2688 7640 2752
rect 7704 2688 7720 2752
rect 7784 2688 7792 2752
rect 7472 2687 7792 2688
rect 2576 2208 2896 2209
rect 2576 2144 2584 2208
rect 2648 2144 2664 2208
rect 2728 2144 2744 2208
rect 2808 2144 2824 2208
rect 2888 2144 2896 2208
rect 2576 2143 2896 2144
rect 5840 2208 6160 2209
rect 5840 2144 5848 2208
rect 5912 2144 5928 2208
rect 5992 2144 6008 2208
rect 6072 2144 6088 2208
rect 6152 2144 6160 2208
rect 5840 2143 6160 2144
rect 9104 2208 9424 2209
rect 9104 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9272 2208
rect 9336 2144 9352 2208
rect 9416 2144 9424 2208
rect 9104 2143 9424 2144
<< via3 >>
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 7480 11452 7544 11456
rect 7480 11396 7484 11452
rect 7484 11396 7540 11452
rect 7540 11396 7544 11452
rect 7480 11392 7544 11396
rect 7560 11452 7624 11456
rect 7560 11396 7564 11452
rect 7564 11396 7620 11452
rect 7620 11396 7624 11452
rect 7560 11392 7624 11396
rect 7640 11452 7704 11456
rect 7640 11396 7644 11452
rect 7644 11396 7700 11452
rect 7700 11396 7704 11452
rect 7640 11392 7704 11396
rect 7720 11452 7784 11456
rect 7720 11396 7724 11452
rect 7724 11396 7780 11452
rect 7780 11396 7784 11452
rect 7720 11392 7784 11396
rect 2584 10908 2648 10912
rect 2584 10852 2588 10908
rect 2588 10852 2644 10908
rect 2644 10852 2648 10908
rect 2584 10848 2648 10852
rect 2664 10908 2728 10912
rect 2664 10852 2668 10908
rect 2668 10852 2724 10908
rect 2724 10852 2728 10908
rect 2664 10848 2728 10852
rect 2744 10908 2808 10912
rect 2744 10852 2748 10908
rect 2748 10852 2804 10908
rect 2804 10852 2808 10908
rect 2744 10848 2808 10852
rect 2824 10908 2888 10912
rect 2824 10852 2828 10908
rect 2828 10852 2884 10908
rect 2884 10852 2888 10908
rect 2824 10848 2888 10852
rect 5848 10908 5912 10912
rect 5848 10852 5852 10908
rect 5852 10852 5908 10908
rect 5908 10852 5912 10908
rect 5848 10848 5912 10852
rect 5928 10908 5992 10912
rect 5928 10852 5932 10908
rect 5932 10852 5988 10908
rect 5988 10852 5992 10908
rect 5928 10848 5992 10852
rect 6008 10908 6072 10912
rect 6008 10852 6012 10908
rect 6012 10852 6068 10908
rect 6068 10852 6072 10908
rect 6008 10848 6072 10852
rect 6088 10908 6152 10912
rect 6088 10852 6092 10908
rect 6092 10852 6148 10908
rect 6148 10852 6152 10908
rect 6088 10848 6152 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 9272 10908 9336 10912
rect 9272 10852 9276 10908
rect 9276 10852 9332 10908
rect 9332 10852 9336 10908
rect 9272 10848 9336 10852
rect 9352 10908 9416 10912
rect 9352 10852 9356 10908
rect 9356 10852 9412 10908
rect 9412 10852 9416 10908
rect 9352 10848 9416 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 7480 10364 7544 10368
rect 7480 10308 7484 10364
rect 7484 10308 7540 10364
rect 7540 10308 7544 10364
rect 7480 10304 7544 10308
rect 7560 10364 7624 10368
rect 7560 10308 7564 10364
rect 7564 10308 7620 10364
rect 7620 10308 7624 10364
rect 7560 10304 7624 10308
rect 7640 10364 7704 10368
rect 7640 10308 7644 10364
rect 7644 10308 7700 10364
rect 7700 10308 7704 10364
rect 7640 10304 7704 10308
rect 7720 10364 7784 10368
rect 7720 10308 7724 10364
rect 7724 10308 7780 10364
rect 7780 10308 7784 10364
rect 7720 10304 7784 10308
rect 2584 9820 2648 9824
rect 2584 9764 2588 9820
rect 2588 9764 2644 9820
rect 2644 9764 2648 9820
rect 2584 9760 2648 9764
rect 2664 9820 2728 9824
rect 2664 9764 2668 9820
rect 2668 9764 2724 9820
rect 2724 9764 2728 9820
rect 2664 9760 2728 9764
rect 2744 9820 2808 9824
rect 2744 9764 2748 9820
rect 2748 9764 2804 9820
rect 2804 9764 2808 9820
rect 2744 9760 2808 9764
rect 2824 9820 2888 9824
rect 2824 9764 2828 9820
rect 2828 9764 2884 9820
rect 2884 9764 2888 9820
rect 2824 9760 2888 9764
rect 5848 9820 5912 9824
rect 5848 9764 5852 9820
rect 5852 9764 5908 9820
rect 5908 9764 5912 9820
rect 5848 9760 5912 9764
rect 5928 9820 5992 9824
rect 5928 9764 5932 9820
rect 5932 9764 5988 9820
rect 5988 9764 5992 9820
rect 5928 9760 5992 9764
rect 6008 9820 6072 9824
rect 6008 9764 6012 9820
rect 6012 9764 6068 9820
rect 6068 9764 6072 9820
rect 6008 9760 6072 9764
rect 6088 9820 6152 9824
rect 6088 9764 6092 9820
rect 6092 9764 6148 9820
rect 6148 9764 6152 9820
rect 6088 9760 6152 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 9272 9820 9336 9824
rect 9272 9764 9276 9820
rect 9276 9764 9332 9820
rect 9332 9764 9336 9820
rect 9272 9760 9336 9764
rect 9352 9820 9416 9824
rect 9352 9764 9356 9820
rect 9356 9764 9412 9820
rect 9412 9764 9416 9820
rect 9352 9760 9416 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 7480 9276 7544 9280
rect 7480 9220 7484 9276
rect 7484 9220 7540 9276
rect 7540 9220 7544 9276
rect 7480 9216 7544 9220
rect 7560 9276 7624 9280
rect 7560 9220 7564 9276
rect 7564 9220 7620 9276
rect 7620 9220 7624 9276
rect 7560 9216 7624 9220
rect 7640 9276 7704 9280
rect 7640 9220 7644 9276
rect 7644 9220 7700 9276
rect 7700 9220 7704 9276
rect 7640 9216 7704 9220
rect 7720 9276 7784 9280
rect 7720 9220 7724 9276
rect 7724 9220 7780 9276
rect 7780 9220 7784 9276
rect 7720 9216 7784 9220
rect 2584 8732 2648 8736
rect 2584 8676 2588 8732
rect 2588 8676 2644 8732
rect 2644 8676 2648 8732
rect 2584 8672 2648 8676
rect 2664 8732 2728 8736
rect 2664 8676 2668 8732
rect 2668 8676 2724 8732
rect 2724 8676 2728 8732
rect 2664 8672 2728 8676
rect 2744 8732 2808 8736
rect 2744 8676 2748 8732
rect 2748 8676 2804 8732
rect 2804 8676 2808 8732
rect 2744 8672 2808 8676
rect 2824 8732 2888 8736
rect 2824 8676 2828 8732
rect 2828 8676 2884 8732
rect 2884 8676 2888 8732
rect 2824 8672 2888 8676
rect 5848 8732 5912 8736
rect 5848 8676 5852 8732
rect 5852 8676 5908 8732
rect 5908 8676 5912 8732
rect 5848 8672 5912 8676
rect 5928 8732 5992 8736
rect 5928 8676 5932 8732
rect 5932 8676 5988 8732
rect 5988 8676 5992 8732
rect 5928 8672 5992 8676
rect 6008 8732 6072 8736
rect 6008 8676 6012 8732
rect 6012 8676 6068 8732
rect 6068 8676 6072 8732
rect 6008 8672 6072 8676
rect 6088 8732 6152 8736
rect 6088 8676 6092 8732
rect 6092 8676 6148 8732
rect 6148 8676 6152 8732
rect 6088 8672 6152 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 9272 8732 9336 8736
rect 9272 8676 9276 8732
rect 9276 8676 9332 8732
rect 9332 8676 9336 8732
rect 9272 8672 9336 8676
rect 9352 8732 9416 8736
rect 9352 8676 9356 8732
rect 9356 8676 9412 8732
rect 9412 8676 9416 8732
rect 9352 8672 9416 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 7480 8188 7544 8192
rect 7480 8132 7484 8188
rect 7484 8132 7540 8188
rect 7540 8132 7544 8188
rect 7480 8128 7544 8132
rect 7560 8188 7624 8192
rect 7560 8132 7564 8188
rect 7564 8132 7620 8188
rect 7620 8132 7624 8188
rect 7560 8128 7624 8132
rect 7640 8188 7704 8192
rect 7640 8132 7644 8188
rect 7644 8132 7700 8188
rect 7700 8132 7704 8188
rect 7640 8128 7704 8132
rect 7720 8188 7784 8192
rect 7720 8132 7724 8188
rect 7724 8132 7780 8188
rect 7780 8132 7784 8188
rect 7720 8128 7784 8132
rect 2584 7644 2648 7648
rect 2584 7588 2588 7644
rect 2588 7588 2644 7644
rect 2644 7588 2648 7644
rect 2584 7584 2648 7588
rect 2664 7644 2728 7648
rect 2664 7588 2668 7644
rect 2668 7588 2724 7644
rect 2724 7588 2728 7644
rect 2664 7584 2728 7588
rect 2744 7644 2808 7648
rect 2744 7588 2748 7644
rect 2748 7588 2804 7644
rect 2804 7588 2808 7644
rect 2744 7584 2808 7588
rect 2824 7644 2888 7648
rect 2824 7588 2828 7644
rect 2828 7588 2884 7644
rect 2884 7588 2888 7644
rect 2824 7584 2888 7588
rect 5848 7644 5912 7648
rect 5848 7588 5852 7644
rect 5852 7588 5908 7644
rect 5908 7588 5912 7644
rect 5848 7584 5912 7588
rect 5928 7644 5992 7648
rect 5928 7588 5932 7644
rect 5932 7588 5988 7644
rect 5988 7588 5992 7644
rect 5928 7584 5992 7588
rect 6008 7644 6072 7648
rect 6008 7588 6012 7644
rect 6012 7588 6068 7644
rect 6068 7588 6072 7644
rect 6008 7584 6072 7588
rect 6088 7644 6152 7648
rect 6088 7588 6092 7644
rect 6092 7588 6148 7644
rect 6148 7588 6152 7644
rect 6088 7584 6152 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 9272 7644 9336 7648
rect 9272 7588 9276 7644
rect 9276 7588 9332 7644
rect 9332 7588 9336 7644
rect 9272 7584 9336 7588
rect 9352 7644 9416 7648
rect 9352 7588 9356 7644
rect 9356 7588 9412 7644
rect 9412 7588 9416 7644
rect 9352 7584 9416 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 7480 7100 7544 7104
rect 7480 7044 7484 7100
rect 7484 7044 7540 7100
rect 7540 7044 7544 7100
rect 7480 7040 7544 7044
rect 7560 7100 7624 7104
rect 7560 7044 7564 7100
rect 7564 7044 7620 7100
rect 7620 7044 7624 7100
rect 7560 7040 7624 7044
rect 7640 7100 7704 7104
rect 7640 7044 7644 7100
rect 7644 7044 7700 7100
rect 7700 7044 7704 7100
rect 7640 7040 7704 7044
rect 7720 7100 7784 7104
rect 7720 7044 7724 7100
rect 7724 7044 7780 7100
rect 7780 7044 7784 7100
rect 7720 7040 7784 7044
rect 2584 6556 2648 6560
rect 2584 6500 2588 6556
rect 2588 6500 2644 6556
rect 2644 6500 2648 6556
rect 2584 6496 2648 6500
rect 2664 6556 2728 6560
rect 2664 6500 2668 6556
rect 2668 6500 2724 6556
rect 2724 6500 2728 6556
rect 2664 6496 2728 6500
rect 2744 6556 2808 6560
rect 2744 6500 2748 6556
rect 2748 6500 2804 6556
rect 2804 6500 2808 6556
rect 2744 6496 2808 6500
rect 2824 6556 2888 6560
rect 2824 6500 2828 6556
rect 2828 6500 2884 6556
rect 2884 6500 2888 6556
rect 2824 6496 2888 6500
rect 5848 6556 5912 6560
rect 5848 6500 5852 6556
rect 5852 6500 5908 6556
rect 5908 6500 5912 6556
rect 5848 6496 5912 6500
rect 5928 6556 5992 6560
rect 5928 6500 5932 6556
rect 5932 6500 5988 6556
rect 5988 6500 5992 6556
rect 5928 6496 5992 6500
rect 6008 6556 6072 6560
rect 6008 6500 6012 6556
rect 6012 6500 6068 6556
rect 6068 6500 6072 6556
rect 6008 6496 6072 6500
rect 6088 6556 6152 6560
rect 6088 6500 6092 6556
rect 6092 6500 6148 6556
rect 6148 6500 6152 6556
rect 6088 6496 6152 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 9272 6556 9336 6560
rect 9272 6500 9276 6556
rect 9276 6500 9332 6556
rect 9332 6500 9336 6556
rect 9272 6496 9336 6500
rect 9352 6556 9416 6560
rect 9352 6500 9356 6556
rect 9356 6500 9412 6556
rect 9412 6500 9416 6556
rect 9352 6496 9416 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 7480 6012 7544 6016
rect 7480 5956 7484 6012
rect 7484 5956 7540 6012
rect 7540 5956 7544 6012
rect 7480 5952 7544 5956
rect 7560 6012 7624 6016
rect 7560 5956 7564 6012
rect 7564 5956 7620 6012
rect 7620 5956 7624 6012
rect 7560 5952 7624 5956
rect 7640 6012 7704 6016
rect 7640 5956 7644 6012
rect 7644 5956 7700 6012
rect 7700 5956 7704 6012
rect 7640 5952 7704 5956
rect 7720 6012 7784 6016
rect 7720 5956 7724 6012
rect 7724 5956 7780 6012
rect 7780 5956 7784 6012
rect 7720 5952 7784 5956
rect 2584 5468 2648 5472
rect 2584 5412 2588 5468
rect 2588 5412 2644 5468
rect 2644 5412 2648 5468
rect 2584 5408 2648 5412
rect 2664 5468 2728 5472
rect 2664 5412 2668 5468
rect 2668 5412 2724 5468
rect 2724 5412 2728 5468
rect 2664 5408 2728 5412
rect 2744 5468 2808 5472
rect 2744 5412 2748 5468
rect 2748 5412 2804 5468
rect 2804 5412 2808 5468
rect 2744 5408 2808 5412
rect 2824 5468 2888 5472
rect 2824 5412 2828 5468
rect 2828 5412 2884 5468
rect 2884 5412 2888 5468
rect 2824 5408 2888 5412
rect 5848 5468 5912 5472
rect 5848 5412 5852 5468
rect 5852 5412 5908 5468
rect 5908 5412 5912 5468
rect 5848 5408 5912 5412
rect 5928 5468 5992 5472
rect 5928 5412 5932 5468
rect 5932 5412 5988 5468
rect 5988 5412 5992 5468
rect 5928 5408 5992 5412
rect 6008 5468 6072 5472
rect 6008 5412 6012 5468
rect 6012 5412 6068 5468
rect 6068 5412 6072 5468
rect 6008 5408 6072 5412
rect 6088 5468 6152 5472
rect 6088 5412 6092 5468
rect 6092 5412 6148 5468
rect 6148 5412 6152 5468
rect 6088 5408 6152 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 9272 5468 9336 5472
rect 9272 5412 9276 5468
rect 9276 5412 9332 5468
rect 9332 5412 9336 5468
rect 9272 5408 9336 5412
rect 9352 5468 9416 5472
rect 9352 5412 9356 5468
rect 9356 5412 9412 5468
rect 9412 5412 9416 5468
rect 9352 5408 9416 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 7480 4924 7544 4928
rect 7480 4868 7484 4924
rect 7484 4868 7540 4924
rect 7540 4868 7544 4924
rect 7480 4864 7544 4868
rect 7560 4924 7624 4928
rect 7560 4868 7564 4924
rect 7564 4868 7620 4924
rect 7620 4868 7624 4924
rect 7560 4864 7624 4868
rect 7640 4924 7704 4928
rect 7640 4868 7644 4924
rect 7644 4868 7700 4924
rect 7700 4868 7704 4924
rect 7640 4864 7704 4868
rect 7720 4924 7784 4928
rect 7720 4868 7724 4924
rect 7724 4868 7780 4924
rect 7780 4868 7784 4924
rect 7720 4864 7784 4868
rect 2584 4380 2648 4384
rect 2584 4324 2588 4380
rect 2588 4324 2644 4380
rect 2644 4324 2648 4380
rect 2584 4320 2648 4324
rect 2664 4380 2728 4384
rect 2664 4324 2668 4380
rect 2668 4324 2724 4380
rect 2724 4324 2728 4380
rect 2664 4320 2728 4324
rect 2744 4380 2808 4384
rect 2744 4324 2748 4380
rect 2748 4324 2804 4380
rect 2804 4324 2808 4380
rect 2744 4320 2808 4324
rect 2824 4380 2888 4384
rect 2824 4324 2828 4380
rect 2828 4324 2884 4380
rect 2884 4324 2888 4380
rect 2824 4320 2888 4324
rect 5848 4380 5912 4384
rect 5848 4324 5852 4380
rect 5852 4324 5908 4380
rect 5908 4324 5912 4380
rect 5848 4320 5912 4324
rect 5928 4380 5992 4384
rect 5928 4324 5932 4380
rect 5932 4324 5988 4380
rect 5988 4324 5992 4380
rect 5928 4320 5992 4324
rect 6008 4380 6072 4384
rect 6008 4324 6012 4380
rect 6012 4324 6068 4380
rect 6068 4324 6072 4380
rect 6008 4320 6072 4324
rect 6088 4380 6152 4384
rect 6088 4324 6092 4380
rect 6092 4324 6148 4380
rect 6148 4324 6152 4380
rect 6088 4320 6152 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 9272 4380 9336 4384
rect 9272 4324 9276 4380
rect 9276 4324 9332 4380
rect 9332 4324 9336 4380
rect 9272 4320 9336 4324
rect 9352 4380 9416 4384
rect 9352 4324 9356 4380
rect 9356 4324 9412 4380
rect 9412 4324 9416 4380
rect 9352 4320 9416 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 7480 3836 7544 3840
rect 7480 3780 7484 3836
rect 7484 3780 7540 3836
rect 7540 3780 7544 3836
rect 7480 3776 7544 3780
rect 7560 3836 7624 3840
rect 7560 3780 7564 3836
rect 7564 3780 7620 3836
rect 7620 3780 7624 3836
rect 7560 3776 7624 3780
rect 7640 3836 7704 3840
rect 7640 3780 7644 3836
rect 7644 3780 7700 3836
rect 7700 3780 7704 3836
rect 7640 3776 7704 3780
rect 7720 3836 7784 3840
rect 7720 3780 7724 3836
rect 7724 3780 7780 3836
rect 7780 3780 7784 3836
rect 7720 3776 7784 3780
rect 2584 3292 2648 3296
rect 2584 3236 2588 3292
rect 2588 3236 2644 3292
rect 2644 3236 2648 3292
rect 2584 3232 2648 3236
rect 2664 3292 2728 3296
rect 2664 3236 2668 3292
rect 2668 3236 2724 3292
rect 2724 3236 2728 3292
rect 2664 3232 2728 3236
rect 2744 3292 2808 3296
rect 2744 3236 2748 3292
rect 2748 3236 2804 3292
rect 2804 3236 2808 3292
rect 2744 3232 2808 3236
rect 2824 3292 2888 3296
rect 2824 3236 2828 3292
rect 2828 3236 2884 3292
rect 2884 3236 2888 3292
rect 2824 3232 2888 3236
rect 5848 3292 5912 3296
rect 5848 3236 5852 3292
rect 5852 3236 5908 3292
rect 5908 3236 5912 3292
rect 5848 3232 5912 3236
rect 5928 3292 5992 3296
rect 5928 3236 5932 3292
rect 5932 3236 5988 3292
rect 5988 3236 5992 3292
rect 5928 3232 5992 3236
rect 6008 3292 6072 3296
rect 6008 3236 6012 3292
rect 6012 3236 6068 3292
rect 6068 3236 6072 3292
rect 6008 3232 6072 3236
rect 6088 3292 6152 3296
rect 6088 3236 6092 3292
rect 6092 3236 6148 3292
rect 6148 3236 6152 3292
rect 6088 3232 6152 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 9272 3292 9336 3296
rect 9272 3236 9276 3292
rect 9276 3236 9332 3292
rect 9332 3236 9336 3292
rect 9272 3232 9336 3236
rect 9352 3292 9416 3296
rect 9352 3236 9356 3292
rect 9356 3236 9412 3292
rect 9412 3236 9416 3292
rect 9352 3232 9416 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 7480 2748 7544 2752
rect 7480 2692 7484 2748
rect 7484 2692 7540 2748
rect 7540 2692 7544 2748
rect 7480 2688 7544 2692
rect 7560 2748 7624 2752
rect 7560 2692 7564 2748
rect 7564 2692 7620 2748
rect 7620 2692 7624 2748
rect 7560 2688 7624 2692
rect 7640 2748 7704 2752
rect 7640 2692 7644 2748
rect 7644 2692 7700 2748
rect 7700 2692 7704 2748
rect 7640 2688 7704 2692
rect 7720 2748 7784 2752
rect 7720 2692 7724 2748
rect 7724 2692 7780 2748
rect 7780 2692 7784 2748
rect 7720 2688 7784 2692
rect 2584 2204 2648 2208
rect 2584 2148 2588 2204
rect 2588 2148 2644 2204
rect 2644 2148 2648 2204
rect 2584 2144 2648 2148
rect 2664 2204 2728 2208
rect 2664 2148 2668 2204
rect 2668 2148 2724 2204
rect 2724 2148 2728 2204
rect 2664 2144 2728 2148
rect 2744 2204 2808 2208
rect 2744 2148 2748 2204
rect 2748 2148 2804 2204
rect 2804 2148 2808 2204
rect 2744 2144 2808 2148
rect 2824 2204 2888 2208
rect 2824 2148 2828 2204
rect 2828 2148 2884 2204
rect 2884 2148 2888 2204
rect 2824 2144 2888 2148
rect 5848 2204 5912 2208
rect 5848 2148 5852 2204
rect 5852 2148 5908 2204
rect 5908 2148 5912 2204
rect 5848 2144 5912 2148
rect 5928 2204 5992 2208
rect 5928 2148 5932 2204
rect 5932 2148 5988 2204
rect 5988 2148 5992 2204
rect 5928 2144 5992 2148
rect 6008 2204 6072 2208
rect 6008 2148 6012 2204
rect 6012 2148 6068 2204
rect 6068 2148 6072 2204
rect 6008 2144 6072 2148
rect 6088 2204 6152 2208
rect 6088 2148 6092 2204
rect 6092 2148 6148 2204
rect 6148 2148 6152 2204
rect 6088 2144 6152 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 9272 2204 9336 2208
rect 9272 2148 9276 2204
rect 9276 2148 9332 2204
rect 9332 2148 9336 2204
rect 9272 2144 9336 2148
rect 9352 2204 9416 2208
rect 9352 2148 9356 2204
rect 9356 2148 9412 2204
rect 9412 2148 9416 2204
rect 9352 2144 9416 2148
<< metal4 >>
rect 2576 10912 2896 11472
rect 2576 10848 2584 10912
rect 2648 10848 2664 10912
rect 2728 10848 2744 10912
rect 2808 10848 2824 10912
rect 2888 10848 2896 10912
rect 2576 9824 2896 10848
rect 2576 9760 2584 9824
rect 2648 9760 2664 9824
rect 2728 9760 2744 9824
rect 2808 9760 2824 9824
rect 2888 9760 2896 9824
rect 2576 8736 2896 9760
rect 2576 8672 2584 8736
rect 2648 8672 2664 8736
rect 2728 8672 2744 8736
rect 2808 8672 2824 8736
rect 2888 8672 2896 8736
rect 2576 7648 2896 8672
rect 2576 7584 2584 7648
rect 2648 7584 2664 7648
rect 2728 7584 2744 7648
rect 2808 7584 2824 7648
rect 2888 7584 2896 7648
rect 2576 6560 2896 7584
rect 2576 6496 2584 6560
rect 2648 6496 2664 6560
rect 2728 6496 2744 6560
rect 2808 6496 2824 6560
rect 2888 6496 2896 6560
rect 2576 5472 2896 6496
rect 2576 5408 2584 5472
rect 2648 5408 2664 5472
rect 2728 5408 2744 5472
rect 2808 5408 2824 5472
rect 2888 5408 2896 5472
rect 2576 4384 2896 5408
rect 2576 4320 2584 4384
rect 2648 4320 2664 4384
rect 2728 4320 2744 4384
rect 2808 4320 2824 4384
rect 2888 4320 2896 4384
rect 2576 3296 2896 4320
rect 2576 3232 2584 3296
rect 2648 3232 2664 3296
rect 2728 3232 2744 3296
rect 2808 3232 2824 3296
rect 2888 3232 2896 3296
rect 2576 2208 2896 3232
rect 2576 2144 2584 2208
rect 2648 2144 2664 2208
rect 2728 2144 2744 2208
rect 2808 2144 2824 2208
rect 2888 2144 2896 2208
rect 2576 2128 2896 2144
rect 4208 11456 4528 11472
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 5840 10912 6160 11472
rect 5840 10848 5848 10912
rect 5912 10848 5928 10912
rect 5992 10848 6008 10912
rect 6072 10848 6088 10912
rect 6152 10848 6160 10912
rect 5840 9824 6160 10848
rect 5840 9760 5848 9824
rect 5912 9760 5928 9824
rect 5992 9760 6008 9824
rect 6072 9760 6088 9824
rect 6152 9760 6160 9824
rect 5840 8736 6160 9760
rect 5840 8672 5848 8736
rect 5912 8672 5928 8736
rect 5992 8672 6008 8736
rect 6072 8672 6088 8736
rect 6152 8672 6160 8736
rect 5840 7648 6160 8672
rect 5840 7584 5848 7648
rect 5912 7584 5928 7648
rect 5992 7584 6008 7648
rect 6072 7584 6088 7648
rect 6152 7584 6160 7648
rect 5840 6560 6160 7584
rect 5840 6496 5848 6560
rect 5912 6496 5928 6560
rect 5992 6496 6008 6560
rect 6072 6496 6088 6560
rect 6152 6496 6160 6560
rect 5840 5472 6160 6496
rect 5840 5408 5848 5472
rect 5912 5408 5928 5472
rect 5992 5408 6008 5472
rect 6072 5408 6088 5472
rect 6152 5408 6160 5472
rect 5840 4384 6160 5408
rect 5840 4320 5848 4384
rect 5912 4320 5928 4384
rect 5992 4320 6008 4384
rect 6072 4320 6088 4384
rect 6152 4320 6160 4384
rect 5840 3296 6160 4320
rect 5840 3232 5848 3296
rect 5912 3232 5928 3296
rect 5992 3232 6008 3296
rect 6072 3232 6088 3296
rect 6152 3232 6160 3296
rect 5840 2208 6160 3232
rect 5840 2144 5848 2208
rect 5912 2144 5928 2208
rect 5992 2144 6008 2208
rect 6072 2144 6088 2208
rect 6152 2144 6160 2208
rect 5840 2128 6160 2144
rect 7472 11456 7792 11472
rect 7472 11392 7480 11456
rect 7544 11392 7560 11456
rect 7624 11392 7640 11456
rect 7704 11392 7720 11456
rect 7784 11392 7792 11456
rect 7472 10368 7792 11392
rect 7472 10304 7480 10368
rect 7544 10304 7560 10368
rect 7624 10304 7640 10368
rect 7704 10304 7720 10368
rect 7784 10304 7792 10368
rect 7472 9280 7792 10304
rect 7472 9216 7480 9280
rect 7544 9216 7560 9280
rect 7624 9216 7640 9280
rect 7704 9216 7720 9280
rect 7784 9216 7792 9280
rect 7472 8192 7792 9216
rect 7472 8128 7480 8192
rect 7544 8128 7560 8192
rect 7624 8128 7640 8192
rect 7704 8128 7720 8192
rect 7784 8128 7792 8192
rect 7472 7104 7792 8128
rect 7472 7040 7480 7104
rect 7544 7040 7560 7104
rect 7624 7040 7640 7104
rect 7704 7040 7720 7104
rect 7784 7040 7792 7104
rect 7472 6016 7792 7040
rect 7472 5952 7480 6016
rect 7544 5952 7560 6016
rect 7624 5952 7640 6016
rect 7704 5952 7720 6016
rect 7784 5952 7792 6016
rect 7472 4928 7792 5952
rect 7472 4864 7480 4928
rect 7544 4864 7560 4928
rect 7624 4864 7640 4928
rect 7704 4864 7720 4928
rect 7784 4864 7792 4928
rect 7472 3840 7792 4864
rect 7472 3776 7480 3840
rect 7544 3776 7560 3840
rect 7624 3776 7640 3840
rect 7704 3776 7720 3840
rect 7784 3776 7792 3840
rect 7472 2752 7792 3776
rect 7472 2688 7480 2752
rect 7544 2688 7560 2752
rect 7624 2688 7640 2752
rect 7704 2688 7720 2752
rect 7784 2688 7792 2752
rect 7472 2128 7792 2688
rect 9104 10912 9424 11472
rect 9104 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9272 10912
rect 9336 10848 9352 10912
rect 9416 10848 9424 10912
rect 9104 9824 9424 10848
rect 9104 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9272 9824
rect 9336 9760 9352 9824
rect 9416 9760 9424 9824
rect 9104 8736 9424 9760
rect 9104 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9272 8736
rect 9336 8672 9352 8736
rect 9416 8672 9424 8736
rect 9104 7648 9424 8672
rect 9104 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9272 7648
rect 9336 7584 9352 7648
rect 9416 7584 9424 7648
rect 9104 6560 9424 7584
rect 9104 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9272 6560
rect 9336 6496 9352 6560
rect 9416 6496 9424 6560
rect 9104 5472 9424 6496
rect 9104 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9272 5472
rect 9336 5408 9352 5472
rect 9416 5408 9424 5472
rect 9104 4384 9424 5408
rect 9104 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9272 4384
rect 9336 4320 9352 4384
rect 9416 4320 9424 4384
rect 9104 3296 9424 4320
rect 9104 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9272 3296
rect 9336 3232 9352 3296
rect 9416 3232 9424 3296
rect 9104 2208 9424 3232
rect 9104 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9272 2208
rect 9336 2144 9352 2208
rect 9416 2144 9424 2208
rect 9104 2128 9424 2144
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1748 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output2
timestamp 1624635492
transform -1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19
timestamp 1624635492
transform 1 0 2852 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1624635492
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output3
timestamp 1624635492
transform -1 0 4968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30
timestamp 1624635492
transform 1 0 3864 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1624635492
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1624635492
transform 1 0 4968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1624635492
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_58
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output4
timestamp 1624635492
transform -1 0 7636 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output5
timestamp 1624635492
transform -1 0 7544 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1624635492
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_70
timestamp 1624635492
transform 1 0 7544 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output6
timestamp 1624635492
transform -1 0 8648 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1624635492
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_82
timestamp 1624635492
transform 1 0 8648 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output7
timestamp 1624635492
transform 1 0 9476 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_100
timestamp 1624635492
transform 1 0 10304 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_90 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 9384 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_95
timestamp 1624635492
transform 1 0 9844 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 10856 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 10856 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1624635492
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  conb_1\[0\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_15
timestamp 1624635492
transform 1 0 2484 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1624635492
transform 1 0 2944 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_28
timestamp 1624635492
transform 1 0 3680 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  conb_1\[3\]
timestamp 1624635492
transform 1 0 4968 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_45
timestamp 1624635492
transform 1 0 5244 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  conb_1\[4\]
timestamp 1624635492
transform 1 0 6532 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_57
timestamp 1624635492
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1624635492
transform 1 0 6808 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  conb_1\[5\]
timestamp 1624635492
transform 1 0 8004 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_74
timestamp 1624635492
transform 1 0 7912 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1624635492
transform 1 0 8280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1624635492
transform 1 0 10212 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 10856 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  conb_1\[1\]
timestamp 1624635492
transform -1 0 2944 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1624635492
transform 1 0 2484 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_20
timestamp 1624635492
transform 1 0 2944 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  conb_1\[2\]
timestamp 1624635492
transform 1 0 3680 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_31
timestamp 1624635492
transform 1 0 3956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_43
timestamp 1624635492
transform 1 0 5060 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1624635492
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_70
timestamp 1624635492
transform 1 0 7544 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  conb_1\[6\]
timestamp 1624635492
transform 1 0 8464 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1624635492
transform 1 0 8280 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_83
timestamp 1624635492
transform 1 0 8740 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output8
timestamp 1624635492
transform 1 0 9476 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_95
timestamp 1624635492
transform 1 0 9844 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 10856 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1624635492
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1624635492
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1624635492
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1624635492
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1624635492
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1624635492
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_99
timestamp 1624635492
transform 1 0 10212 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 10856 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1624635492
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1624635492
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1624635492
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_51
timestamp 1624635492
transform 1 0 5796 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1624635492
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  conb_1\[7\]
timestamp 1624635492
transform 1 0 8924 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_82
timestamp 1624635492
transform 1 0 8648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_88
timestamp 1624635492
transform 1 0 9200 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_100
timestamp 1624635492
transform 1 0 10304 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 10856 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1624635492
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1624635492
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1624635492
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1624635492
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1624635492
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1624635492
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1624635492
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1624635492
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1624635492
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1624635492
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1624635492
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1624635492
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1624635492
transform 1 0 10212 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_94
timestamp 1624635492
transform 1 0 9752 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_102
timestamp 1624635492
transform 1 0 10488 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 10856 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 10856 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1624635492
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1624635492
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1624635492
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1624635492
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1624635492
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1624635492
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1624635492
transform 1 0 10212 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 10856 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1624635492
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1624635492
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1624635492
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1624635492
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1624635492
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1624635492
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_94
timestamp 1624635492
transform 1 0 9752 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1624635492
transform 1 0 10488 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 10856 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1624635492
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624635492
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1624635492
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1624635492
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1624635492
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1624635492
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_99
timestamp 1624635492
transform 1 0 10212 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 10856 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1624635492
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1624635492
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1624635492
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1624635492
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1624635492
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_82
timestamp 1624635492
transform 1 0 8648 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_94
timestamp 1624635492
transform 1 0 9752 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_102
timestamp 1624635492
transform 1 0 10488 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 10856 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1624635492
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1624635492
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1624635492
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1624635492
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_66
timestamp 1624635492
transform 1 0 7176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1624635492
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_87
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_99
timestamp 1624635492
transform 1 0 10212 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 10856 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1624635492
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1624635492
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1624635492
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1624635492
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1624635492
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1624635492
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1624635492
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1624635492
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1624635492
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1624635492
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1624635492
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1624635492
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_87
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_94
timestamp 1624635492
transform 1 0 9752 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_102
timestamp 1624635492
transform 1 0 10488 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_99
timestamp 1624635492
transform 1 0 10212 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 10856 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 10856 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1624635492
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1624635492
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1624635492
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1624635492
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1624635492
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1624635492
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_94
timestamp 1624635492
transform 1 0 9752 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_102
timestamp 1624635492
transform 1 0 10488 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 10856 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1624635492
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1624635492
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1624635492
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1624635492
transform 1 0 6440 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_54
timestamp 1624635492
transform 1 0 6072 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_59
timestamp 1624635492
transform 1 0 6532 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_71
timestamp 1624635492
transform 1 0 7636 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_83
timestamp 1624635492
transform 1 0 8740 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_88
timestamp 1624635492
transform 1 0 9200 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_100
timestamp 1624635492
transform 1 0 10304 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 10856 0 -1 11424
box -38 -48 314 592
<< labels >>
rlabel metal2 s 754 0 810 800 6 x[0]
port 0 nsew signal tristate
rlabel metal2 s 2226 0 2282 800 6 x[1]
port 1 nsew signal tristate
rlabel metal2 s 3698 0 3754 800 6 x[2]
port 2 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 x[3]
port 3 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 x[4]
port 4 nsew signal tristate
rlabel metal2 s 8206 0 8262 800 6 x[5]
port 5 nsew signal tristate
rlabel metal2 s 9678 0 9734 800 6 x[6]
port 6 nsew signal tristate
rlabel metal2 s 11150 0 11206 800 6 x[7]
port 7 nsew signal tristate
rlabel metal4 s 9104 2128 9424 11472 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 5840 2128 6160 11472 6 VPWR
port 9 nsew power bidirectional
rlabel metal4 s 2576 2128 2896 11472 6 VPWR
port 10 nsew power bidirectional
rlabel metal4 s 7472 2128 7792 11472 6 VGND
port 11 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 11472 6 VGND
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 12000 14000
<< end >>
