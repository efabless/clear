* NGSPICE file created from bottom_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt bottom_tile VGND VPWR ccff_head ccff_head_1 ccff_tail ccff_tail_0 chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23]
+ chanx_left_in[24] chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28]
+ chanx_left_in[29] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23]
+ chanx_left_out[24] chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28]
+ chanx_left_out[29] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in_0[0]
+ chanx_right_in_0[10] chanx_right_in_0[11] chanx_right_in_0[12] chanx_right_in_0[13]
+ chanx_right_in_0[14] chanx_right_in_0[15] chanx_right_in_0[16] chanx_right_in_0[17]
+ chanx_right_in_0[18] chanx_right_in_0[19] chanx_right_in_0[1] chanx_right_in_0[20]
+ chanx_right_in_0[21] chanx_right_in_0[22] chanx_right_in_0[23] chanx_right_in_0[24]
+ chanx_right_in_0[25] chanx_right_in_0[26] chanx_right_in_0[27] chanx_right_in_0[28]
+ chanx_right_in_0[29] chanx_right_in_0[2] chanx_right_in_0[3] chanx_right_in_0[4]
+ chanx_right_in_0[5] chanx_right_in_0[6] chanx_right_in_0[7] chanx_right_in_0[8]
+ chanx_right_in_0[9] chanx_right_out_0[0] chanx_right_out_0[10] chanx_right_out_0[11]
+ chanx_right_out_0[12] chanx_right_out_0[13] chanx_right_out_0[14] chanx_right_out_0[15]
+ chanx_right_out_0[16] chanx_right_out_0[17] chanx_right_out_0[18] chanx_right_out_0[19]
+ chanx_right_out_0[1] chanx_right_out_0[20] chanx_right_out_0[21] chanx_right_out_0[22]
+ chanx_right_out_0[23] chanx_right_out_0[24] chanx_right_out_0[25] chanx_right_out_0[26]
+ chanx_right_out_0[27] chanx_right_out_0[28] chanx_right_out_0[29] chanx_right_out_0[2]
+ chanx_right_out_0[3] chanx_right_out_0[4] chanx_right_out_0[5] chanx_right_out_0[6]
+ chanx_right_out_0[7] chanx_right_out_0[8] chanx_right_out_0[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1]
+ chany_top_in[20] chany_top_in[21] chany_top_in[22] chany_top_in[23] chany_top_in[24]
+ chany_top_in[25] chany_top_in[26] chany_top_in[27] chany_top_in[28] chany_top_in[29]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10]
+ chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15]
+ chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1]
+ chany_top_out[20] chany_top_out[21] chany_top_out[22] chany_top_out[23] chany_top_out[24]
+ chany_top_out[25] chany_top_out[26] chany_top_out[27] chany_top_out[28] chany_top_out[29]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] gfpga_pad_io_soc_dir[0] gfpga_pad_io_soc_dir[1]
+ gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0] gfpga_pad_io_soc_in[1]
+ gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0] gfpga_pad_io_soc_out[1]
+ gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] isol_n prog_clk prog_reset_top_in
+ reset_top_in right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_ right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ test_enable_top_in top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
+ top_width_0_height_0_subtile_0__pin_inpad_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ top_width_0_height_0_subtile_2__pin_inpad_0_ top_width_0_height_0_subtile_3__pin_inpad_0_
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_1__0_.mem_right_track_12.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input92_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net96 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_42.mux_l2_in_0__246 VGND VGND VPWR VPWR net246 sb_1__0_.mux_top_track_42.mux_l2_in_0__246/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mux_left_track_29.mux_l1_in_1_ net39 net86 sb_1__0_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_0.mux_l1_in_0_ net91 net73 sb_1__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_1__0_.mem_right_track_36.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_4.mux_l2_in_1_ net244 net17 sb_1__0_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_1__0_.mem_top_track_14.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_14.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__124__A net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_ net255 net58 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_left_track_53.mux_l2_in_1__215 VGND VGND VPWR VPWR net215 sb_1__0_.mux_left_track_53.mux_l2_in_1__215/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_32_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_14.mux_l2_in_1__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_1__0_.mem_top_track_4.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
X_200_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
X_131_ sb_1__0_.mux_left_track_5.out VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_1__0_.mem_left_track_11.ccff_head
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_7_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_1__0_.mem_top_track_44.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_46.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input55_A chanx_right_in_0[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_28.mux_l1_in_0_ net29 net59 sb_1__0_.mem_top_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_30.mux_l1_in_0_ net28 net58 sb_1__0_.mem_top_track_30.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_28_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_ net35 net4 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
X_114_ net35 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_42.mux_l2_in_0_ net246 sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_42.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A0 net39 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_1__0_.mem_right_track_2.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input18_A chanx_left_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0 net25 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__0_.mux_right_track_36.mux_l2_in_1__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_1__0_.mem_right_track_10.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_input85_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_29.mux_l1_in_0_ net68 net80 sb_1__0_.mem_left_track_29.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_12.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_4.mux_l2_in_0_ sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__140__A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_ net27 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_24.mux_l1_in_1__237 VGND VGND VPWR VPWR net237 sb_1__0_.mux_top_track_24.mux_l1_in_1__237/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.out sky130_fd_sc_hd__clkbuf_1
XFILLER_9_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput210 net210 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__buf_12
XFILLER_28_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_130_ sb_1__0_.mux_left_track_7.out VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
XFILLER_23_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input48_A chanx_right_in_0[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__135__A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_top_track_32.mux_l1_in_0__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_4.mux_l1_in_1_ net47 net50 sb_1__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input102_A right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_113_ net34 VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_ net41 net10 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1 net8 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk sb_1__0_.mem_right_track_0.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_30.out sky130_fd_sc_hd__clkbuf_1
XFILLER_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_42.mux_l1_in_0_ net27 net104 sb_1__0_.mem_top_track_42.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput110 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND VGND VPWR
+ VPWR net110 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input30_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__143__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_24.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input78_A chany_top_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_29.mux_l2_in_1__262 VGND VGND VPWR VPWR net262 sb_1__0_.mux_left_track_29.mux_l2_in_1__262/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__138__A net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A0 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_40.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_18.out sky130_fd_sc_hd__clkbuf_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
Xoutput200 net200 VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_189_ sb_1__0_.mux_top_track_8.out VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__151__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_4.mux_l1_in_0_ net106 net103 sb_1__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_28_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_5.mux_l2_in_1__A1 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_28.mux_l3_in_0_ sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_28.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_112_ net62 VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_ net48 net17 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input60_A chanx_right_in_0[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__146__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_0_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mux_top_track_16.mux_l2_in_1__232 VGND VGND VPWR VPWR net232 sb_1__0_.mux_top_track_16.mux_l2_in_1__232/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mux_right_track_28.mux_l2_in_1_ net222 sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_28.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_4.mux_l2_in_1__244 VGND VGND VPWR VPWR net244 sb_1__0_.mux_top_track_4.mux_l2_in_1__244/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_21_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput100 right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_ VGND VGND
+ VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input23_A chanx_left_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_1__0_.mem_top_track_32.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_32.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_36.mux_l1_in_1__243 VGND VGND VPWR VPWR net243 sb_1__0_.mux_top_track_36.mux_l1_in_1__243/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_28.mux_l1_in_2_ net14 net9 sb_1__0_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_1__0_.mem_right_track_36.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA__154__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_46.out sky130_fd_sc_hd__clkbuf_1
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_12.mux_l3_in_0_ sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sb_1__0_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input90_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput201 net201 VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_1__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_188_ sb_1__0_.mux_top_track_10.out VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_4_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\] net98 VGND VGND VPWR VPWR net112
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_12.mux_l2_in_1_ net230 net11 sb_1__0_.mem_top_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_16_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_ net51 net20 cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_111_ sb_1__0_.mux_left_track_45.out VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input53_A chanx_right_in_0[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_28.mux_l2_in_0_ sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_28.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_38_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput101 right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_ VGND VGND
+ VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_1__0_.mem_top_track_30.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_32.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input16_A chanx_left_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_13.mux_l3_in_0_ sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_8_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_9_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input8_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_28.mux_l1_in_1_ net101 net74 sb_1__0_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_29_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_1__0_.mem_right_track_36.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_36.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_45.out sky130_fd_sc_hd__clkbuf_1
XFILLER_23_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_13.mux_l2_in_1_ net260 sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_left_track_13.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input83_A chany_top_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_0__A0 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput202 net202 VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_12
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_187_ sb_1__0_.mux_top_track_12.out VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_2
XFILLER_37_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_4_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_12.mux_l2_in_0_ net36 sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_left_track_13.mux_l1_in_2_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net56 sb_1__0_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A0 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_110_ net60 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_ sb_1__0_.mux_left_track_3.out net23
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input46_A chanx_right_in_0[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input100_A right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__0_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_52.out sky130_fd_sc_hd__clkbuf_1
XFILLER_34_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A0 net47 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput102 right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_ VGND VGND
+ VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_31_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_28.mux_l1_in_0_ net66 net78 sb_1__0_.mem_right_track_28.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk sb_1__0_.mem_right_track_28.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_40_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_1__0_.mem_left_track_53.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_6.mux_l1_in_3_ net227 net29 sb_1__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_37_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_13.mux_l2_in_0_ sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_13.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input76_A chany_top_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput203 net203 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_186_ sb_1__0_.mux_top_track_14.out VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_0_0_prog_clk net1 net98 VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
Xsb_1__0_.mux_left_track_13.mux_l1_in_1_ net42 net74 sb_1__0_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_2__A1 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_1__0_.mem_top_track_50.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_50.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input39_A chanx_right_in_0[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_6.mux_l3_in_0_ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sb_1__0_.mem_right_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
X_169_ sb_1__0_.mux_top_track_48.out VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_12.mux_l1_in_0_ net41 net109 sb_1__0_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk
+ cbx_1__0_.cbx_8__0_.ccff_head net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_24.mux_l2_in_0_ sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_24.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_3__A1 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput103 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND VGND VPWR
+ VPWR net103 sky130_fd_sc_hd__buf_2
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mux_right_track_6.mux_l2_in_1_ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_6_0_prog_clk sb_1__0_.mem_left_track_21.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_21.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.out sky130_fd_sc_hd__clkbuf_2
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_4_0_prog_clk sb_1__0_.mem_left_track_5.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_input21_A chanx_left_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_1__0_.mem_left_track_53.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_53.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_24.mux_l1_in_1_ net237 net32 sb_1__0_.mem_top_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_40.mux_l2_in_0__245 VGND VGND VPWR VPWR net245 sb_1__0_.mux_top_track_40.mux_l2_in_0__245/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mux_right_track_6.mux_l1_in_2_ net16 net101 sb_1__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_0.mux_l1_in_3_ net228 net21 sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_26_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input69_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__A1 net59 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput204 net204 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A0 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_185_ sb_1__0_.mux_top_track_16.out VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_13.mux_l1_in_0_ net66 net78 sb_1__0_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_1__0_.mem_top_track_48.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_50.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_168_ sb_1__0_.mux_top_track_50.out VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_left_track_37.mux_l3_in_0_ sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_left_track_37.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_0.mux_l3_in_0_ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sb_1__0_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_37_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input51_A chanx_right_in_0[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput104 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND VGND VPWR
+ VPWR net104 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_right_track_6.mux_l2_in_0_ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_37.mux_l2_in_1_ net212 top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__0_.mem_left_track_37.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input99_A right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_top_track_0.mux_l2_in_1_ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_1__0_.mem_left_track_21.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_21.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_1__A0 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_1__0_.mem_left_track_5.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_5.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input14_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_1__0_.mem_left_track_45.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_53.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_24.mux_l1_in_0_ net62 net107 sb_1__0_.mem_top_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_35_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_6.mux_l1_in_1_ net99 net88 sb_1__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_36.mux_l2_in_0_ sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_input6_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_0.mux_l1_in_2_ net24 net51 sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_14_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_22.mux_l1_in_1__236 VGND VGND VPWR VPWR net236 sb_1__0_.mux_top_track_22.mux_l1_in_1__236/LO
+ sky130_fd_sc_hd__conb_1
Xoutput205 net205 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
XFILLER_28_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_46.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_13.mux_l2_in_1__260 VGND VGND VPWR VPWR net260 sb_1__0_.mux_left_track_13.mux_l2_in_1__260/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input81_A chany_top_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_1__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_184_ sb_1__0_.mux_top_track_18.out VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A0 net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_36.mux_l1_in_1_ net243 net14 sb_1__0_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_28.mux_l2_in_1__222 VGND VGND VPWR VPWR net222 sb_1__0_.mux_right_track_28.mux_l2_in_1__222/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_36_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_ net256 sb_1__0_.mux_left_track_53.out
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
X_167_ net19 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_3__A1 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input44_A chanx_right_in_0[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_1__0_.mem_top_track_24.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_24.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_38_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mux_right_track_12.mux_l3_in_0_ sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xinput105 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND VGND VPWR
+ VPWR net105 sky130_fd_sc_hd__clkbuf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_ net34 net32 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_37.mux_l2_in_0_ sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_37.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_12_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_top_track_0.mux_l2_in_0_ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_1__0_.mem_left_track_13.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_21.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk sb_1__0_.mem_right_track_28.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_38_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_1__0_.mem_left_track_3.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_12.mux_l2_in_1_ net219 sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_12.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_6.mux_l1_in_0_ net70 net82 sb_1__0_.mem_right_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_left_track_37.mux_l1_in_1_ net38 net87 sb_1__0_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_0.mux_l1_in_1_ net53 net107 sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_1__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A0 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput206 net206 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input109_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_183_ sb_1__0_.mux_top_track_20.out VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input74_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_12.mux_l1_in_2_ net26 net12 sb_1__0_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_38_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_12.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_36.mux_l1_in_0_ net44 net109 sb_1__0_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_9_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_20.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_48.mux_l2_in_0_ net249 sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_48.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_ net26 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
X_166_ net20 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_50.mux_l2_in_0_ net250 sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_50.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input37_A chanx_right_in_0[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_14.out sky130_fd_sc_hd__clkbuf_1
XFILLER_19_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_1__0_.mem_top_track_22.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_24.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_149_ sb_1__0_.mux_right_track_28.out VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_14.mux_l2_in_1__231 VGND VGND VPWR VPWR net231 sb_1__0_.mux_top_track_14.mux_l2_in_1__231/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput106 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND VGND VPWR
+ VPWR net106 sky130_fd_sc_hd__buf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_ sb_1__0_.mux_left_track_29.out net9
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_10.mux_l2_in_1__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_1__0_.mem_right_track_28.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_28.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_12.mux_l2_in_0_ sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_12.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_left_track_37.mux_l1_in_0_ net69 net81 sb_1__0_.mem_left_track_37.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_0.mux_l1_in_0_ net104 net109 sb_1__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_14_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xoutput207 net207 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__buf_12
XFILLER_36_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_182_ sb_1__0_.mux_top_track_22.out VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_top_track_0.mux_l1_in_3__228 VGND VGND VPWR VPWR net228 sb_1__0_.mux_top_track_0.mux_l1_in_3__228/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_0__A0 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input67_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_12.mux_l1_in_1_ net99 net86 sb_1__0_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_2.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
X_165_ net22 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_42.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_13.out sky130_fd_sc_hd__clkbuf_1
XFILLER_24_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_148_ net9 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_48.mux_l1_in_0_ net10 net107 sb_1__0_.mem_top_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A0 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput107 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND VGND VPWR
+ VPWR net107 sky130_fd_sc_hd__buf_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_ net47 net16 cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_50.mux_l1_in_0_ net15 net108 sb_1__0_.mem_top_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_1__0_.mem_right_track_20.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_1__0_.mem_left_track_45.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_38_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_0_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input97_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input12_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_1__0_.mem_top_track_10.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput208 net208 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__buf_12
Xsb_1__0_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.out sky130_fd_sc_hd__clkbuf_1
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_181_ sb_1__0_.mux_top_track_24.out VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_2.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_right_track_12.mux_l1_in_0_ net68 net80 sb_1__0_.mem_right_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_1__0_.mem_top_track_42.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_42.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_9_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_52.mux_l1_in_1__226 VGND VGND VPWR VPWR net226 sb_1__0_.mux_right_track_52.mux_l1_in_1__226/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_36.mux_l3_in_0_ sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_right_track_36.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_164_ sb_1__0_.mux_top_track_58.out VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
XFILLER_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_2__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net111 net97 VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_5_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XANTENNA__106__A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_147_ net8 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A0 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_8.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk sb_1__0_.mem_left_track_13.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_21_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_2__A1 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_36.mux_l2_in_1_ net223 net8 sb_1__0_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xinput108 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND VGND VPWR
+ VPWR net108 sky130_fd_sc_hd__buf_2
Xsb_1__0_.mux_top_track_2.mux_l2_in_1__234 VGND VGND VPWR VPWR net234 sb_1__0_.mux_top_track_2.mux_l2_in_1__234/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_ sb_1__0_.mux_left_track_11.out net19
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_11.mux_l1_in_3__259 VGND VGND VPWR VPWR net259 sb_1__0_.mux_left_track_11.mux_l1_in_3__259/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_37_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input42_A chanx_right_in_0[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_1__0_.mem_left_track_45.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_45.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_1__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput90 chany_top_in[7] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mux_top_track_18.mux_l3_in_0_ sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X sb_1__0_.mem_top_track_18.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__256 VGND VGND VPWR VPWR net256 cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__256/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_58.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_58.out sky130_fd_sc_hd__clkbuf_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net94 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_37_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_10.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__114__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput209 net209 VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__buf_12
XFILLER_36_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_34.mux_l2_in_0__242 VGND VGND VPWR VPWR net242 sb_1__0_.mux_top_track_34.mux_l2_in_0__242/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_180_ sb_1__0_.mux_top_track_26.out VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_1__0_.mem_top_track_0.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__0_.mux_top_track_18.mux_l2_in_1_ net233 net7 sb_1__0_.mem_top_track_18.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA__109__A net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk sb_1__0_.mem_top_track_40.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_42.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input107_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input72_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_163_ sb_1__0_.mux_right_track_0.out VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0 net46 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_1__0_.mem_top_track_16.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_16.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_5.mux_l3_in_0_ sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__122__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_146_ net7 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_2__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_8.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_1__0_.mem_left_track_13.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_13.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_36.mux_l2_in_0_ sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_36.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0 net35 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput109 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND VGND VPWR
+ VPWR net109 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_1__0_.mem_top_track_48.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_48.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_ sb_1__0_.mux_left_track_5.out net22
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail net97
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_12_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_1__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input35_A chanx_right_in_0[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_21.mux_l3_in_0_ sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_left_track_21.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA__117__A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_129_ net51 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_1__0_.mem_left_track_37.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput91 chany_top_in[8] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
Xinput80 chany_top_in[25] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_left_track_5.mux_l2_in_1_ net214 top_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_1__0_.mem_left_track_5.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_right_track_36.mux_l1_in_1_ net102 net63 sb_1__0_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_1__0_.mem_right_track_4.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_8_0_prog_clk cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
+ net98 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfrtp_2
Xsb_1__0_.mux_left_track_21.mux_l2_in_1_ net261 sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_left_track_21.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_10.ccff_head
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_right_track_2.mux_l3_in_0_ sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A0 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.out sky130_fd_sc_hd__clkbuf_1
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_top_track_18.mux_l2_in_0_ net33 sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_18.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__125__A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_21.mux_l1_in_2_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net55 sb_1__0_.mem_left_track_21.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_20.mux_l2_in_0_ sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A0 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_2.mux_l2_in_1_ net220 sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
X_162_ sb_1__0_.mux_right_track_2.out VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input65_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_44.mux_l1_in_1__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_1__0_.mem_top_track_16.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_16.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xinput1 ccff_head VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_1__A0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_145_ sb_1__0_.mux_right_track_36.out VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_6.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
Xsb_1__0_.mux_top_track_20.mux_l1_in_1_ net235 net5 sb_1__0_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_1__0_.mem_left_track_11.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_21_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1 net4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_1__0_.mem_top_track_46.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_48.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_right_track_2.mux_l1_in_2_ net32 net18 sb_1__0_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput190 net190 VGND VGND VPWR VPWR chany_top_out[25] sky130_fd_sc_hd__buf_12
XANTENNA_input28_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ sb_1__0_.mux_left_track_11.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_5.mux_l2_in_0_ sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_5.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_21_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput70 chany_top_in[16] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
Xinput92 chany_top_in[9] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
Xinput81 chany_top_in[26] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__A1 net58 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_35_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_36.mux_l1_in_0_ net65 net77 sb_1__0_.mem_right_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_31_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_1__0_.mem_right_track_4.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_21.mux_l2_in_0_ sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_21.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_right_track_4.mux_l1_in_1__A0 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_5.mux_l1_in_1__A1 net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input95_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_20.mux_l1_in_1__235 VGND VGND VPWR VPWR net235 sb_1__0_.mux_top_track_20.mux_l1_in_1__235/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_5.mux_l1_in_1_ net60 net47 sb_1__0_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A0 net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_right_track_52.mux_l1_in_1__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_14_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input10_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_left_track_21.mux_l1_in_1_ net41 net85 sb_1__0_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_input2_A ccff_head_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_45.mux_l2_in_1__213 VGND VGND VPWR VPWR net213 sb_1__0_.mux_left_track_45.mux_l2_in_1__213/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__0_.mux_top_track_18.mux_l1_in_0__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_2.mux_l2_in_0_ sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_161_ sb_1__0_.mux_right_track_4.out VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input58_A chanx_right_in_0[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__136__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_1__0_.mem_top_track_14.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_16.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 ccff_head_1 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_18.mux_l1_in_0_ net37 net104 sb_1__0_.mem_top_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_144_ net5 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_20.mux_l1_in_0_ net35 net105 sb_1__0_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_2.mux_l1_in_1_ net100 net90 sb_1__0_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_32.mux_l2_in_0_ net241 sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_32.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_50.mux_l2_in_0__250 VGND VGND VPWR VPWR net250 sb_1__0_.mux_top_track_50.mux_l2_in_0__250/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_24_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput180 net180 VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_12
Xoutput191 net191 VGND VGND VPWR VPWR chany_top_out[26] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_127_ sb_1__0_.mux_left_track_13.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput82 chany_top_in[27] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_1
Xinput71 chany_top_in[17] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_1
Xinput60 chanx_right_in_0[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_top_track_16.mux_l2_in_1__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput93 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input40_A chanx_right_in_0[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_1__0_.mem_right_track_2.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__144__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input88_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_left_track_5.mux_l1_in_0_ net92 net75 sb_1__0_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__139__A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_26.mux_l1_in_0__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_7.mux_l2_in_1__216 VGND VGND VPWR VPWR net216 sb_1__0_.mux_left_track_7.mux_l2_in_1__216/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mux_left_track_21.mux_l1_in_0_ net67 net79 sb_1__0_.mem_left_track_21.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_160_ sb_1__0_.mux_right_track_6.out VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_6.mux_l3_in_0_ sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_top_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_45.mux_l3_in_0_ sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X sb_1__0_.mem_left_track_45.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA__152__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 chanx_left_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input105_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input70_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_143_ net4 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_top_track_12.mux_l2_in_1__230 VGND VGND VPWR VPWR net230 sb_1__0_.mux_top_track_12.mux_l2_in_1__230/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__147__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_2.mux_l1_in_0_ net72 net84 sb_1__0_.mem_right_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_6.mux_l2_in_1_ net252 sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_top_track_6.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_12_0_prog_clk sb_1__0_.mem_left_track_37.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_37.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput192 net192 VGND VGND VPWR VPWR chany_top_out[27] sky130_fd_sc_hd__buf_12
Xoutput181 net181 VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_12
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_ net257 net56 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
Xoutput170 net170 VGND VGND VPWR VPWR chanx_right_out_0[7] sky130_fd_sc_hd__buf_12
XFILLER_28_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A0 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A0 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_45.mux_l2_in_1_ net213 net37 sb_1__0_.mem_left_track_45.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_126_ net48 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A0 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput50 chanx_right_in_0[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
Xinput72 chany_top_in[18] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
Xinput61 chanx_right_in_0[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
Xinput83 chany_top_in[28] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_1
Xinput94 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input33_A chanx_right_in_0[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_34.mux_l1_in_0__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_6.mux_l1_in_2_ net16 net46 sb_1__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_109_ net59 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_32.mux_l1_in_0_ net26 net56 sb_1__0_.mem_top_track_32.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_ net62 net31 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_44.mux_l2_in_0_ net247 sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_44.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_27_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_right_track_10.mux_l1_in_3__218 VGND VGND VPWR VPWR net218 sb_1__0_.mux_right_track_10.mux_l1_in_3__218/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__155__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X net112 VGND VGND
+ VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_1__0_.mem_top_track_34.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_34.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A0 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput4 chanx_left_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
XFILLER_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_142_ net32 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input63_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_6.mux_l2_in_0_ sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_1__0_.mem_left_track_37.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_37.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A0 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_20.mux_l3_in_0_ sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_20.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_ net25 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
Xoutput193 net193 VGND VGND VPWR VPWR chany_top_out[28] sky130_fd_sc_hd__buf_12
Xoutput182 net182 VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_12
Xoutput171 net171 VGND VGND VPWR VPWR chanx_right_out_0[8] sky130_fd_sc_hd__buf_12
Xoutput160 net160 VGND VGND VPWR VPWR chanx_right_out_0[25] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_2__A1 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_45.mux_l2_in_0_ net88 sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_left_track_45.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_42.mux_l1_in_0__A1 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_125_ net47 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_2__A1 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput73 chany_top_in[19] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput51 chanx_right_in_0[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
Xinput84 chany_top_in[29] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_1
Xinput40 chanx_right_in_0[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput62 chanx_right_in_0[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0 net42 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput95 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_right_track_4.mux_l2_in_1__224 VGND VGND VPWR VPWR net224 sb_1__0_.mux_right_track_4.mux_l2_in_1__224/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input26_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_108_ net58 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A0 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_6.mux_l1_in_1_ net49 net107 sb_1__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__254 VGND VGND VPWR VPWR net254 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__254/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mux_right_track_20.mux_l2_in_1_ net221 sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_20.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_ net39 net8 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_1_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_27_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk sb_1__0_.mem_top_track_32.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_34.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_2__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input93_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_32.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_right_track_20.mux_l1_in_2_ net25 net11 sb_1__0_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_36_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_44.mux_l1_in_0_ net31 net105 sb_1__0_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_1__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XFILLER_32_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_50.mux_l1_in_0__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_26.out sky130_fd_sc_hd__clkbuf_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_141_ sb_1__0_.mux_right_track_44.out VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input56_A chanx_right_in_0[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_1__0_.mem_left_track_29.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_37.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_2__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput161 net161 VGND VGND VPWR VPWR chanx_right_out_0[26] sky130_fd_sc_hd__buf_12
Xoutput150 net150 VGND VGND VPWR VPWR chanx_right_out_0[16] sky130_fd_sc_hd__buf_12
Xoutput194 net194 VGND VGND VPWR VPWR chany_top_out[29] sky130_fd_sc_hd__buf_12
Xoutput183 net183 VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_12
Xoutput172 net172 VGND VGND VPWR VPWR chanx_right_out_0[9] sky130_fd_sc_hd__buf_12
XANTENNA_input110_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_124_ net46 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput85 chany_top_in[2] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 chanx_right_in_0[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
Xinput74 chany_top_in[1] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 chanx_right_in_0[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
Xinput63 chany_top_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_left_track_37.mux_l2_in_1__A1 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2
Xinput96 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_40_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.out sky130_fd_sc_hd__clkbuf_1
XFILLER_28_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input19_A chanx_left_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_1__0_.mem_left_track_1.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
X_107_ sb_1__0_.mux_left_track_53.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_2__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_top_track_6.mux_l1_in_0_ net104 net109 sb_1__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_ net46 net15 cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_20.mux_l2_in_0_ sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_20.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_45.mux_l1_in_0_ net70 net82 sb_1__0_.mem_left_track_45.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_32.mux_l2_in_0__241 VGND VGND VPWR VPWR net241 sb_1__0_.mux_top_track_32.mux_l2_in_0__241/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input86_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_20.mux_l1_in_1_ net100 net85 sb_1__0_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A0 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 chanx_left_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_140_ net30 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input49_A chanx_right_in_0[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_1__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_45.mux_l2_in_1__A1 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_14.mux_l3_in_0_ sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X sb_1__0_.mem_top_track_14.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_37_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput195 net195 VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_12
Xoutput184 net184 VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_12
Xoutput173 net173 VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_12
Xoutput140 net140 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xoutput162 net162 VGND VGND VPWR VPWR chanx_right_out_0[27] sky130_fd_sc_hd__buf_12
Xoutput151 net151 VGND VGND VPWR VPWR chanx_right_out_0[17] sky130_fd_sc_hd__buf_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input103_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_48.out sky130_fd_sc_hd__clkbuf_1
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_123_ sb_1__0_.mux_left_track_21.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_6_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_1.mux_l1_in_3_ net258 top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput75 chany_top_in[20] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput64 chany_top_in[10] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
Xinput86 chany_top_in[3] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput53 chanx_right_in_0[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput42 chanx_right_in_0[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
Xinput97 isol_n VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_48.mux_l2_in_0__249 VGND VGND VPWR VPWR net249 sb_1__0_.mux_top_track_48.mux_l2_in_0__249/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_16_446 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_14.mux_l2_in_1_ net231 net9 sb_1__0_.mem_top_track_14.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_1__0_.mem_left_track_1.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_1.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_106_ net56 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_ sb_1__0_.mux_left_track_7.out net21
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A0 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input31_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_1.mux_l3_in_0_ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sb_1__0_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input79_A chany_top_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_20.mux_l1_in_0_ net67 net79 sb_1__0_.mem_right_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_1_0_prog_clk sb_1__0_.mem_left_track_7.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_53.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_53.out sky130_fd_sc_hd__clkbuf_1
XFILLER_1_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_left_track_53.mux_l2_in_1__A1 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_2__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0 net34 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 chanx_left_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_1.mux_l2_in_1_ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_19_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_199_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk sb_1__0_.mem_top_track_20.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput174 net174 VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_12
Xoutput196 net196 VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_12
Xoutput185 net185 VGND VGND VPWR VPWR chany_top_out[20] sky130_fd_sc_hd__buf_12
Xoutput130 net130 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
Xoutput163 net163 VGND VGND VPWR VPWR chanx_right_out_0[28] sky130_fd_sc_hd__buf_12
Xoutput152 net152 VGND VGND VPWR VPWR chanx_right_out_0[18] sky130_fd_sc_hd__buf_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_122_ net43 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input61_A chanx_right_in_0[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput54 chanx_right_in_0[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 chanx_right_in_0[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_top_track_4.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_1.mux_l1_in_2_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net34 sb_1__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_2
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
Xinput98 prog_reset_top_in VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_16
Xinput76 chany_top_in[21] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput65 chany_top_in[11] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
Xinput87 chany_top_in[4] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_2.mux_l2_in_1__220 VGND VGND VPWR VPWR net220 sb_1__0_.mux_right_track_2.mux_l2_in_1__220/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_top_track_14.mux_l2_in_0_ net61 sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_14.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
X_105_ net55 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_1__0_.mem_left_track_1.ccff_head
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_ sb_1__0_.mux_left_track_1.out net24
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_2__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input24_A chanx_left_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk sb_1__0_.mem_top_track_58.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_0.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_5.mux_l2_in_1__214 VGND VGND VPWR VPWR net214 sb_1__0_.mux_left_track_5.mux_l2_in_1__214/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_1__0_.mem_left_track_7.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_7.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_39_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input91_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_1__A1 net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_1.mux_l2_in_0_ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_1.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_7_0_prog_clk sb_1__0_.mem_left_track_29.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_198_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_1__0_.mem_top_track_18.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_44.mux_l2_in_0_ sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput175 net175 VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_12
Xoutput186 net186 VGND VGND VPWR VPWR chany_top_out[21] sky130_fd_sc_hd__buf_12
Xoutput197 net197 VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_12
Xoutput120 net120 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
Xoutput142 net142 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
Xoutput164 net164 VGND VGND VPWR VPWR chanx_right_out_0[29] sky130_fd_sc_hd__buf_12
Xoutput153 net153 VGND VGND VPWR VPWR chanx_right_out_0[19] sky130_fd_sc_hd__buf_12
XFILLER_28_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_121_ net42 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input54_A chanx_right_in_0[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput77 chany_top_in[22] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput66 chany_top_in[12] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xinput88 chany_top_in[5] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_left_track_1.mux_l1_in_1_ net51 net90 sb_1__0_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xinput55 chanx_right_in_0[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
Xinput44 chanx_right_in_0[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
Xinput33 chanx_right_in_0[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
XFILLER_14_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput99 right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_ VGND VGND
+ VPWR VPWR net99 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_left_track_1.mux_l1_in_3__258 VGND VGND VPWR VPWR net258 sb_1__0_.mux_left_track_1.mux_l1_in_3__258/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_10_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_104_ net44 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_right_track_44.mux_l1_in_1_ net225 net7 sb_1__0_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_22_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_1__0_.mem_top_track_26.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_26.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_13_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input17_A chanx_left_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_1__0_.mem_top_track_50.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_58.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_14.mux_l1_in_0_ net39 net110 sb_1__0_.mem_top_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input9_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_26.mux_l2_in_0_ sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_26.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_12_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk sb_1__0_.mem_left_track_5.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_input84_A chany_top_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_15_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_26.mux_l1_in_1_ net238 net30 sb_1__0_.mem_top_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_1__0_.mem_left_track_29.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_29.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_197_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_1__A0 net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput121 net121 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xoutput143 net143 VGND VGND VPWR VPWR chanx_right_out_0[0] sky130_fd_sc_hd__buf_12
Xoutput187 net187 VGND VGND VPWR VPWR chany_top_out[22] sky130_fd_sc_hd__buf_12
Xoutput198 net198 VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_12
Xoutput176 net176 VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_12
Xoutput165 net165 VGND VGND VPWR VPWR chanx_right_out_0[2] sky130_fd_sc_hd__buf_12
Xoutput154 net154 VGND VGND VPWR VPWR chanx_right_out_0[1] sky130_fd_sc_hd__buf_12
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_120_ net41 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input47_A chanx_right_in_0[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_1.mux_l1_in_0_ net72 net84 sb_1__0_.mem_left_track_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_34_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput78 chany_top_in[23] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput67 chany_top_in[13] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
Xinput89 chany_top_in[6] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_1
Xinput45 chanx_right_in_0[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput34 chanx_right_in_0[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput56 chanx_right_in_0[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_top_track_48.mux_l1_in_0__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input101_A right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_14.mux_l1_in_0__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_right_track_44.mux_l1_in_0_ net64 net76 sb_1__0_.mem_right_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_1__0_.mem_top_track_24.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_26.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_2.mux_l3_in_0_ sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_31_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_2.mux_l2_in_1_ net234 sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_top_track_2.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input77_A chany_top_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_1__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_26.mux_l1_in_0_ net60 net108 sb_1__0_.mem_top_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_1__0_.mem_left_track_21.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_196_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mux_top_track_2.mux_l1_in_2_ net18 net48 sb_1__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput177 net177 VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_12
Xoutput122 net122 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
Xsb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_1__0_.mem_top_track_4.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xoutput166 net166 VGND VGND VPWR VPWR chanx_right_out_0[3] sky130_fd_sc_hd__buf_12
Xoutput111 net111 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xoutput144 net144 VGND VGND VPWR VPWR chanx_right_out_0[10] sky130_fd_sc_hd__buf_12
Xoutput155 net155 VGND VGND VPWR VPWR chanx_right_out_0[20] sky130_fd_sc_hd__buf_12
Xoutput199 net199 VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR chany_top_out[23] sky130_fd_sc_hd__buf_12
XFILLER_23_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_40.mux_l2_in_0_ net245 sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_40.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A0 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
+ net98 VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput79 chany_top_in[24] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
Xinput68 chany_top_in[14] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
Xinput46 chanx_right_in_0[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
X_179_ sb_1__0_.mux_top_track_28.out VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_2
Xinput35 chanx_right_in_0[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_2
Xinput57 chanx_right_in_0[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
Xinput24 chanx_left_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__104__A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input22_A chanx_left_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_1__0_.mem_right_track_10.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_2.mux_l2_in_0_ sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_12.mux_l2_in_1__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_left_track_53.mux_l3_in_0_ sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X cbx_1__0_.cbx_8__0_.ccff_head
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_12.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_right_track_12.mux_l2_in_1__219 VGND VGND VPWR VPWR net219 sb_1__0_.mux_right_track_12.mux_l2_in_1__219/LO
+ sky130_fd_sc_hd__conb_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_195_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_8.mux_l2_in_1__253 VGND VGND VPWR VPWR net253 sb_1__0_.mux_top_track_8.mux_l2_in_1__253/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__112__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_right_track_0.mux_l1_in_1__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_2.mux_l1_in_1_ net52 net108 sb_1__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_58.mux_l2_in_0__251 VGND VGND VPWR VPWR net251 sb_1__0_.mux_top_track_58.mux_l2_in_0__251/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_4.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0 net41 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_9_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput189 net189 VGND VGND VPWR VPWR chany_top_out[24] sky130_fd_sc_hd__buf_12
Xoutput178 net178 VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
Xoutput134 net134 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
Xoutput112 net112 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xoutput167 net167 VGND VGND VPWR VPWR chanx_right_out_0[4] sky130_fd_sc_hd__buf_12
Xoutput145 net145 VGND VGND VPWR VPWR chanx_right_out_0[11] sky130_fd_sc_hd__buf_12
Xoutput156 net156 VGND VGND VPWR VPWR chanx_right_out_0[21] sky130_fd_sc_hd__buf_12
XFILLER_28_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_1__0_.mem_top_track_44.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mux_top_track_22.mux_l1_in_0__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_53.mux_l2_in_1_ net215 net35 sb_1__0_.mem_left_track_53.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_19_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 chanx_right_in_0[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_2
Xinput14 chanx_left_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput47 chanx_right_in_0[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_2
Xinput69 chany_top_in[15] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
X_178_ sb_1__0_.mux_top_track_30.out VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
Xinput58 chanx_right_in_0[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_2
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input52_A chanx_right_in_0[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2__A0 net27 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_1__0_.mem_right_track_0.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_top_track_40.mux_l1_in_0_ net3 net103 sb_1__0_.mem_top_track_40.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_22.out sky130_fd_sc_hd__clkbuf_1
XFILLER_25_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__120__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_30.mux_l2_in_0__240 VGND VGND VPWR VPWR net240 sb_1__0_.mux_top_track_30.mux_l2_in_0__240/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input15_A chanx_left_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_16.out sky130_fd_sc_hd__clkbuf_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_3.mux_l2_in_1__211 VGND VGND VPWR VPWR net211 sb_1__0_.mux_left_track_3.mux_l2_in_1__211/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk sb_1__0_.mem_right_track_10.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net95 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XANTENNA_input7_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_12.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_12.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mux_top_track_30.mux_l1_in_0__A1 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input82_A chany_top_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_194_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_top_track_2.mux_l1_in_0_ net105 net110 sb_1__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_2.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1 net10 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xoutput179 net179 VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
Xoutput124 net124 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
Xoutput168 net168 VGND VGND VPWR VPWR chanx_right_out_0[5] sky130_fd_sc_hd__buf_12
Xoutput146 net146 VGND VGND VPWR VPWR chanx_right_out_0[12] sky130_fd_sc_hd__buf_12
Xoutput157 net157 VGND VGND VPWR VPWR chanx_right_out_0[22] sky130_fd_sc_hd__buf_12
XFILLER_36_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk sb_1__0_.mem_top_track_42.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_53.mux_l2_in_0_ net89 sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_left_track_53.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput48 chanx_right_in_0[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_2
X_177_ sb_1__0_.mux_top_track_32.out VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_2
Xinput37 chanx_right_in_0[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
Xinput59 chanx_right_in_0[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_2
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mux_top_track_46.mux_l2_in_0__248 VGND VGND VPWR VPWR net248 sb_1__0_.mux_top_track_46.mux_l2_in_0__248/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input45_A chanx_right_in_0[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_1__0_.mem_top_track_18.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_18.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_50.out sky130_fd_sc_hd__clkbuf_1
XFILLER_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_21.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_21.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_21.out sky130_fd_sc_hd__clkbuf_1
XANTENNA__118__A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_1__0_.mem_right_track_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_18_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_2__A1 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A0 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_10.mux_l3_in_0_ sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_1__0_.mem_right_track_10.ccff_head
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_11_0_prog_clk sb_1__0_.mem_right_track_6.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_2_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__126__A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xsb_1__0_.mux_right_track_44.mux_l1_in_1__225 VGND VGND VPWR VPWR net225 sb_1__0_.mux_right_track_44.mux_l1_in_1__225/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk sb_1__0_.mem_top_track_10.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_23_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_3.mux_l2_in_1__A1 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ sb_1__0_.mux_top_track_0.out VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input75_A chany_top_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_10.mux_l2_in_1_ net229 net12 sb_1__0_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_left_track_11.mux_l1_in_3_ net259 top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_1__0_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput125 net125 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput114 net114 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
XFILLER_13_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput136 net136 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
Xoutput169 net169 VGND VGND VPWR VPWR chanx_right_out_0[6] sky130_fd_sc_hd__buf_12
Xoutput147 net147 VGND VGND VPWR VPWR chanx_right_out_0[13] sky130_fd_sc_hd__buf_12
Xoutput158 net158 VGND VGND VPWR VPWR chanx_right_out_0[23] sky130_fd_sc_hd__buf_12
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_176_ sb_1__0_.mux_top_track_34.out VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xinput49 chanx_right_in_0[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput38 chanx_right_in_0[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_2
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 chanx_left_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input38_A chanx_right_in_0[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk sb_1__0_.mem_top_track_18.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_18.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_37.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk sb_1__0_.mem_right_track_0.ccff_head
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
X_159_ net21 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_2
XANTENNA__134__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_53.mux_l1_in_0_ net71 net83 sb_1__0_.mem_left_track_53.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_53.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_left_track_11.mux_l3_in_0_ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sb_1__0_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_7_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__129__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0 net62 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_35_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_11.mux_l2_in_1_ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_1__A1 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk sb_1__0_.mem_right_track_6.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_37.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_37.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_37.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_input20_A chanx_left_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__142__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_35_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_192_ sb_1__0_.mux_top_track_2.out VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input68_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_10.mux_l2_in_0_ sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_left_track_11.mux_l1_in_2_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net58 sb_1__0_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput126 net126 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
Xoutput115 net115 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
Xoutput137 net137 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
Xoutput148 net148 VGND VGND VPWR VPWR chanx_right_out_0[14] sky130_fd_sc_hd__buf_12
XFILLER_9_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput159 net159 VGND VGND VPWR VPWR chanx_right_out_0[24] sky130_fd_sc_hd__buf_12
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A0 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_175_ sb_1__0_.mux_top_track_36.out VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
Xinput39 chanx_right_in_0[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
XANTENNA_sb_1__0_.mux_left_track_29.mux_l1_in_1__A0 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
XFILLER_6_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_10.mux_l1_in_1_ net40 net42 sb_1__0_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_24_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk sb_1__0_.mem_top_track_16.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_18.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_158_ sb_1__0_.mux_right_track_10.out VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__150__A net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_44.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input50_A chanx_right_in_0[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_7.mux_l3_in_0_ sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_right_track_12.mux_l1_in_1__A0 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_1__0_.mem_top_track_30.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_30.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_5_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input98_A prog_reset_top_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1 net31 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_11.mux_l2_in_0_ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_11.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_23_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_21.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_1__0_.mem_right_track_4.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__257 VGND VGND VPWR VPWR net257 cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__257/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input13_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_7.mux_l2_in_1_ net216 sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_left_track_7.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input5_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_left_track_37.mux_l1_in_1__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1 net56 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_191_ sb_1__0_.mux_top_track_4.out VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
Xsb_1__0_.mux_left_track_11.mux_l1_in_1_ net43 net63 sb_1__0_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput127 net127 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
Xoutput116 net116 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput138 net138 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
Xoutput149 net149 VGND VGND VPWR VPWR chanx_right_out_0[15] sky130_fd_sc_hd__buf_12
Xsb_1__0_.mux_right_track_4.mux_l3_in_0_ sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_3_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_6.mux_l1_in_1__A0 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_left_track_7.mux_l1_in_2_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ top_width_0_height_0_subtile_0__pin_inpad_0_ sb_1__0_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_left_track_7.mux_l1_in_1__A1 net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input80_A chany_top_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ sky130_fd_sc_hd__ebufn_1
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_1__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
X_174_ net110 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xinput29 chanx_left_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A0 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__148__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mux_top_track_10.mux_l1_in_0_ net106 net103 sb_1__0_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_5.out sky130_fd_sc_hd__clkbuf_1
XFILLER_30_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_22.mux_l2_in_0_ sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_22.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
X_157_ sb_1__0_.mux_right_track_12.out VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_4.mux_l2_in_1_ net224 sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_4.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input43_A chanx_right_in_0[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_1__0_.mem_top_track_28.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_30.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_1__0_.mux_top_track_22.mux_l1_in_1_ net236 net4 sb_1__0_.mem_top_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_4.mux_l1_in_2_ net30 net17 sb_1__0_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_35_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__156__A net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_10.mux_l1_in_3__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_28.mux_l2_in_0__239 VGND VGND VPWR VPWR net239 sb_1__0_.mux_top_track_28.mux_l2_in_0__239/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_left_track_7.mux_l2_in_0_ sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_7.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_top_track_18.mux_l2_in_1__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ sb_1__0_.mux_top_track_6.out VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_37.mux_l2_in_1__212 VGND VGND VPWR VPWR net212 sb_1__0_.mux_left_track_37.mux_l2_in_1__212/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_1__0_.mem_top_track_36.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mux_left_track_11.mux_l1_in_0_ net65 net77 sb_1__0_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A0 net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput128 net128 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
Xoutput117 net117 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_52.mux_l2_in_0_ sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_7.mux_l1_in_1_ net59 net46 sb_1__0_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input108_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_173_ sb_1__0_.mux_top_track_40.out VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput19 chanx_left_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XANTENNA_input73_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_28.mux_l1_in_0__A1 net59 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_156_ net18 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_right_track_20.mux_l1_in_1__A1 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_52.mux_l1_in_1_ net226 net5 sb_1__0_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_4.mux_l2_in_0_ sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA__159__A net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input36_A chanx_right_in_0[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_139_ net29 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_2
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_22.mux_l1_in_0_ net34 net106 sb_1__0_.mem_top_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_8_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_4.mux_l1_in_1_ net101 net89 sb_1__0_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_34.mux_l2_in_0_ net242 sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_34.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A0 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_11.mux_l1_in_1__A0 net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_right_track_10.mux_l1_in_3_ net218 net28 sb_1__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_39_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk sb_1__0_.mem_top_track_34.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mux_top_track_36.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_6.mux_l2_in_1__252 VGND VGND VPWR VPWR net252 sb_1__0_.mux_top_track_6.mux_l2_in_1__252/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput129 net129 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
Xoutput118 net118 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
XANTENNA_sb_1__0_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_ net254 net59 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_7.mux_l1_in_0_ net64 net76 sb_1__0_.mem_left_track_7.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_172_ sb_1__0_.mux_top_track_42.out VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input66_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_21.mux_l2_in_1__261 VGND VGND VPWR VPWR net261 sb_1__0_.mux_left_track_21.mux_l2_in_1__261/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_155_ net17 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_52.mux_l1_in_0_ net92 net75 sb_1__0_.mem_right_track_52.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_10.mux_l3_in_0_ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X
+ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sb_1__0_.mem_right_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_6_X sky130_fd_sc_hd__mux2_1
XFILLER_33_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_ sb_1__0_.mux_left_track_37.out net5
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_8.mux_l3_in_0_ sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_36.mux_l2_in_1__223 VGND VGND VPWR VPWR net223 sb_1__0_.mux_right_track_36.mux_l2_in_1__223/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail net97
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XANTENNA_sb_1__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input29_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_138_ net28 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_10.mux_l2_in_1_ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_right_track_4.mux_l1_in_0_ net71 net83 sb_1__0_.mem_right_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_20_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_8.mux_l2_in_1_ net253 sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_top_track_8.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_5_0_prog_clk sb_1__0_.mem_left_track_3.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_47 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_44.mux_l1_in_0__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input96_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A0 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_right_track_10.mux_l1_in_2_ net13 net102 sb_1__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_34.mux_l1_in_0_ net25 net55 sb_1__0_.mem_top_track_34.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_8.mux_l1_in_2_ net13 net43 sb_1__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input11_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput119 net119 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xsb_1__0_.mux_top_track_46.mux_l2_in_0_ net248 sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_46.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_ net28 cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input3_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail net98 VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_171_ sb_1__0_.mux_top_track_44.out VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_22_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input59_A chanx_right_in_0[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_44.mux_l2_in_0__247 VGND VGND VPWR VPWR net247 sb_1__0_.mux_top_track_44.mux_l2_in_0__247/LO
+ sky130_fd_sc_hd__conb_1
Xsb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk sb_1__0_.mem_right_track_20.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_27_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_154_ net16 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_ net42 net11 cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_top_track_2.mux_l1_in_1__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_1__0_.mem_right_track_52.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_137_ sb_1__0_.mux_right_track_52.out VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_top_track_0.mux_l1_in_3__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_10.mux_l2_in_0_ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input41_A chanx_right_in_0[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_top_track_8.mux_l2_in_0_ sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_top_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail net97
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_1
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk sb_1__0_.mem_left_track_3.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_3.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input89_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_top_track_10.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_right_track_10.mux_l1_in_1_ net100 net87 sb_1__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_8.mux_l1_in_1_ net45 net108 sb_1__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_1_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_11.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_40.out sky130_fd_sc_hd__clkbuf_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_170_ sb_1__0_.mux_top_track_46.out VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk sb_1__0_.mem_right_track_20.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_20.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input106_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_46.mux_l1_in_0_ net6 net106 sb_1__0_.mem_top_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_153_ sb_1__0_.mux_right_track_20.out VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input71_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_34.out sky130_fd_sc_hd__clkbuf_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_ sb_1__0_.mux_left_track_13.out net18
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_top_track_58.mux_l2_in_0_ net251 sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_right_track_0.ccff_head VGND VGND VPWR VPWR sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_26.mux_l1_in_1__238 VGND VGND VPWR VPWR net238 sb_1__0_.mux_top_track_26.mux_l1_in_1__238/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk sb_1__0_.mem_top_track_22.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_22.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk sb_1__0_.mem_right_track_44.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_52.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A0 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_136_ net26 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
XFILLER_2_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_12_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input34_A chanx_right_in_0[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_119_ sb_1__0_.mux_left_track_29.out VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk sb_1__0_.mem_left_track_1.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__255 VGND VGND VPWR VPWR net255 cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__255/LO
+ sky130_fd_sc_hd__conb_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
+ net98 VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A0 net104 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mux_right_track_10.mux_l1_in_0_ net69 net81 sb_1__0_.mem_right_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_10.mux_l2_in_1__229 VGND VGND VPWR VPWR net229 sb_1__0_.mux_top_track_10.mux_l2_in_1__229/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_8.mux_l1_in_0_ net105 net110 sb_1__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_22_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_12.out sky130_fd_sc_hd__clkbuf_1
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_3_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk sb_1__0_.mem_right_track_12.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A0 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_152_ net13 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input64_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_ sb_1__0_.mux_left_track_7.out net21
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk sb_1__0_.mem_top_track_20.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_22.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_13.mux_l1_in_2__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_135_ net25 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_58.mux_l1_in_0_ net23 net54 sb_1__0_.mem_top_track_58.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_58.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_16.mux_l3_in_0_ sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X sb_1__0_.mem_top_track_16.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_input27_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_118_ net39 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_8_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mux_top_track_6.mux_l1_in_0__A1 net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk sb_1__0_.mem_top_track_28.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_18.mux_l2_in_1__233 VGND VGND VPWR VPWR net233 sb_1__0_.mux_top_track_18.mux_l2_in_1__233/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_top_track_16.mux_l2_in_1_ net232 net8 sb_1__0_.mem_top_track_16.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_1_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input94_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_13_0_prog_clk sb_1__0_.mem_top_track_0.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_3.mux_l3_in_0_ sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_32_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_1__0_.mux_left_track_21.mux_l1_in_2__A1 net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_1__0_.mux_top_track_4.mux_l2_in_1__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_151_ net12 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_1__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ sb_1__0_.mux_left_track_1.out net24
+ cbx_1__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_1__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input57_A chanx_right_in_0[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_28.out sky130_fd_sc_hd__clkbuf_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_3.mux_l2_in_1_ net211 top_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_1__0_.mem_left_track_3.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
X_134_ net14 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_117_ net38 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_0.mux_l3_in_0_ sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_right_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_1.out sky130_fd_sc_hd__clkbuf_2
XFILLER_35_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk sb_1__0_.mem_top_track_26.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_16.mux_l2_in_0_ net57 sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_16.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input87_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A0 net48 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_0.mux_l2_in_1_ net217 sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_right_track_0.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk sb_1__0_.mem_top_track_0.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk sb_1__0_.mem_top_track_40.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_40.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_10_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_0.mux_l2_in_1__217 VGND VGND VPWR VPWR net217 sb_1__0_.mux_right_track_0.mux_l2_in_1__217/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_150_ net11 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_1__0_.mux_top_track_20.mux_l1_in_1__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_0.mux_l1_in_2_ net4 net21 sb_1__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input104_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_6.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
X_133_ sb_1__0_.mux_left_track_1.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_6_0_prog_clk sb_1__0_.mem_left_track_11.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_7_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mux_left_track_3.mux_l2_in_0_ sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__110__A net60 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_20.mux_l2_in_1__221 VGND VGND VPWR VPWR net221 sb_1__0_.mux_right_track_20.mux_l2_in_1__221/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_1__0_.mux_top_track_58.mux_l1_in_0__A0 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_116_ net37 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_1__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B net98
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__105__A net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_left_track_29.mux_l3_in_0_ sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X sb_1__0_.mem_left_track_29.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_5_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_6.mux_l1_in_3__227 VGND VGND VPWR VPWR net227 sb_1__0_.mux_right_track_6.mux_l1_in_3__227/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_3.mux_l1_in_1_ net62 net48 sb_1__0_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_25_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_1__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input32_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net93 cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_12_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_29.mux_l2_in_1_ net262 sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sb_1__0_.mem_left_track_29.mem_out\[1\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A0 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_right_track_0.mux_l2_in_0_ sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_right_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_1__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_1__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net2
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_28.mux_l1_in_2__A0 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_1__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk sb_1__0_.mem_top_track_36.ccff_tail
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_40.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_1__0_.mem_left_track_53.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_10_0_prog_clk sb_1__0_.mem_right_track_12.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__113__A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_top_track_16.mux_l1_in_0_ net38 net103 sb_1__0_.mem_top_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_ sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.out sky130_fd_sc_hd__clkbuf_1
Xsb_1__0_.mux_left_track_29.mux_l1_in_2_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net44 sb_1__0_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mux_top_track_28.mux_l2_in_0_ net239 sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_28.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mux_right_track_0.mux_l1_in_1_ net102 net99 sb_1__0_.mem_right_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_18_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk sb_1__0_.mem_right_track_44.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_1__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_1__0_.mem_top_track_14.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_26_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_30.mux_l2_in_0_ net240 sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
+ sb_1__0_.mem_top_track_30.ccff_tail VGND VGND VPWR VPWR sb_1__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__108__A net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_1__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk sb_1__0_.mem_top_track_6.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_132_ sb_1__0_.mux_left_track_3.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_1__0_.mux_top_track_8.mux_l1_in_1__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_1__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk sb_1__0_.mem_left_track_11.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_left_track_11.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
X_201_ cbx_1__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
+ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input62_A chanx_right_in_0[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk sb_1__0_.mem_top_track_46.mem_out\[0\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_top_track_46.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_37_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mux_right_track_2.mux_l1_in_1__A0 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_115_ sb_1__0_.mux_left_track_37.out VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__121__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_1__0_.mux_left_track_3.mux_l1_in_1__A1 net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_1__0_.mux_top_track_24.mux_l1_in_0__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_1__0_.mux_left_track_3.mux_l1_in_0_ net91 net73 sb_1__0_.mem_left_track_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_1__0_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk sb_1__0_.mem_right_track_2.mem_out\[1\]
+ net98 VGND VGND VPWR VPWR sb_1__0_.mem_right_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input25_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__116__A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_1__0_.mux_left_track_1.mux_l1_in_3__A1 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_left_track_29.mux_l2_in_0_ sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X sb_1__0_.mem_left_track_29.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_1__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_1__0_.mux_top_track_16.mux_l1_in_0__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_1__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net98 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_1__0_.mux_top_track_4.mux_l3_in_0_ sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
+ sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sb_1__0_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_1__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

