magic
tech sky130A
magscale 1 2
timestamp 1625783622
<< locali >>
rect 7021 20315 7055 20417
rect 8861 15351 8895 15589
rect 12817 14263 12851 14433
rect 21097 11543 21131 11645
rect 10057 10523 10091 10693
rect 11897 10523 11931 10761
rect 17693 10523 17727 10693
rect 22017 8619 22051 9605
rect 20913 2907 20947 3009
rect 22017 1411 22051 2533
<< viali >>
rect 2789 20553 2823 20587
rect 11437 20553 11471 20587
rect 16221 20553 16255 20587
rect 4997 20485 5031 20519
rect 7849 20485 7883 20519
rect 10057 20485 10091 20519
rect 12081 20485 12115 20519
rect 12633 20485 12667 20519
rect 13185 20485 13219 20519
rect 13737 20485 13771 20519
rect 16865 20485 16899 20519
rect 17877 20485 17911 20519
rect 18429 20485 18463 20519
rect 18981 20485 19015 20519
rect 19533 20485 19567 20519
rect 7021 20417 7055 20451
rect 15761 20417 15795 20451
rect 1685 20349 1719 20383
rect 2145 20349 2179 20383
rect 2605 20349 2639 20383
rect 3065 20349 3099 20383
rect 4077 20349 4111 20383
rect 4537 20349 4571 20383
rect 5181 20349 5215 20383
rect 5641 20349 5675 20383
rect 5917 20349 5951 20383
rect 6745 20349 6779 20383
rect 7205 20349 7239 20383
rect 7665 20349 7699 20383
rect 8309 20349 8343 20383
rect 8861 20349 8895 20383
rect 9413 20349 9447 20383
rect 9873 20349 9907 20383
rect 10333 20349 10367 20383
rect 10793 20349 10827 20383
rect 15025 20349 15059 20383
rect 16129 20349 16163 20383
rect 18797 20349 18831 20383
rect 20269 20349 20303 20383
rect 21189 20349 21223 20383
rect 7021 20281 7055 20315
rect 11345 20281 11379 20315
rect 12265 20281 12299 20315
rect 12817 20281 12851 20315
rect 13369 20281 13403 20315
rect 13921 20281 13955 20315
rect 15209 20281 15243 20315
rect 15577 20281 15611 20315
rect 16681 20281 16715 20315
rect 17693 20281 17727 20315
rect 18245 20281 18279 20315
rect 19349 20281 19383 20315
rect 20637 20281 20671 20315
rect 20821 20281 20855 20315
rect 21373 20281 21407 20315
rect 1777 20213 1811 20247
rect 2329 20213 2363 20247
rect 3249 20213 3283 20247
rect 4261 20213 4295 20247
rect 4721 20213 4755 20247
rect 5457 20213 5491 20247
rect 6101 20213 6135 20247
rect 6929 20213 6963 20247
rect 7389 20213 7423 20247
rect 8125 20213 8159 20247
rect 8677 20213 8711 20247
rect 9597 20213 9631 20247
rect 10517 20213 10551 20247
rect 10977 20213 11011 20247
rect 14565 20213 14599 20247
rect 20085 20213 20119 20247
rect 1409 20009 1443 20043
rect 2053 20009 2087 20043
rect 2513 20009 2547 20043
rect 2881 20009 2915 20043
rect 3801 20009 3835 20043
rect 4445 20009 4479 20043
rect 6837 20009 6871 20043
rect 9689 20009 9723 20043
rect 11161 20009 11195 20043
rect 12081 20009 12115 20043
rect 17785 20009 17819 20043
rect 19901 20009 19935 20043
rect 3525 19941 3559 19975
rect 5181 19941 5215 19975
rect 5549 19941 5583 19975
rect 7113 19941 7147 19975
rect 10793 19941 10827 19975
rect 14565 19941 14599 19975
rect 15301 19941 15335 19975
rect 15853 19941 15887 19975
rect 17141 19941 17175 19975
rect 20545 19941 20579 19975
rect 4537 19873 4571 19907
rect 5917 19873 5951 19907
rect 6653 19873 6687 19907
rect 7840 19873 7874 19907
rect 10425 19873 10459 19907
rect 11897 19873 11931 19907
rect 12725 19873 12759 19907
rect 14657 19873 14691 19907
rect 15485 19873 15519 19907
rect 16037 19873 16071 19907
rect 17325 19873 17359 19907
rect 17877 19873 17911 19907
rect 19533 19873 19567 19907
rect 19993 19873 20027 19907
rect 21189 19873 21223 19907
rect 4261 19805 4295 19839
rect 7573 19805 7607 19839
rect 9413 19805 9447 19839
rect 12449 19805 12483 19839
rect 14473 19805 14507 19839
rect 16589 19805 16623 19839
rect 18705 19805 18739 19839
rect 20361 19805 20395 19839
rect 6101 19737 6135 19771
rect 10057 19737 10091 19771
rect 15025 19737 15059 19771
rect 21373 19737 21407 19771
rect 4905 19669 4939 19703
rect 8953 19669 8987 19703
rect 13093 19669 13127 19703
rect 7573 19465 7607 19499
rect 18613 19465 18647 19499
rect 19257 19465 19291 19499
rect 7297 19397 7331 19431
rect 18337 19397 18371 19431
rect 8125 19329 8159 19363
rect 8309 19329 8343 19363
rect 9413 19329 9447 19363
rect 16313 19329 16347 19363
rect 16497 19329 16531 19363
rect 4077 19261 4111 19295
rect 5917 19261 5951 19295
rect 9689 19261 9723 19295
rect 10793 19261 10827 19295
rect 12449 19261 12483 19295
rect 14565 19261 14599 19295
rect 14832 19261 14866 19295
rect 16589 19261 16623 19295
rect 17233 19261 17267 19295
rect 18153 19261 18187 19295
rect 18797 19261 18831 19295
rect 19073 19261 19107 19295
rect 19993 19261 20027 19295
rect 20453 19261 20487 19295
rect 3525 19193 3559 19227
rect 4322 19193 4356 19227
rect 6184 19193 6218 19227
rect 8401 19193 8435 19227
rect 11060 19193 11094 19227
rect 12694 19193 12728 19227
rect 17417 19193 17451 19227
rect 20637 19193 20671 19227
rect 21189 19193 21223 19227
rect 21373 19193 21407 19227
rect 5457 19125 5491 19159
rect 8769 19125 8803 19159
rect 9597 19125 9631 19159
rect 10057 19125 10091 19159
rect 12173 19125 12207 19159
rect 13829 19125 13863 19159
rect 15945 19125 15979 19159
rect 16957 19125 16991 19159
rect 20085 19125 20119 19159
rect 3709 18921 3743 18955
rect 4721 18921 4755 18955
rect 5733 18921 5767 18955
rect 7665 18921 7699 18955
rect 11345 18921 11379 18955
rect 14749 18921 14783 18955
rect 16589 18921 16623 18955
rect 17509 18921 17543 18955
rect 19073 18921 19107 18955
rect 19533 18921 19567 18955
rect 20177 18921 20211 18955
rect 8033 18853 8067 18887
rect 13636 18853 13670 18887
rect 20821 18853 20855 18887
rect 2585 18785 2619 18819
rect 4629 18785 4663 18819
rect 5273 18785 5307 18819
rect 7205 18785 7239 18819
rect 10232 18785 10266 18819
rect 12173 18785 12207 18819
rect 12265 18785 12299 18819
rect 13369 18785 13403 18819
rect 16405 18785 16439 18819
rect 17325 18785 17359 18819
rect 18061 18785 18095 18819
rect 19257 18785 19291 18819
rect 19717 18785 19751 18819
rect 20085 18785 20119 18819
rect 20637 18785 20671 18819
rect 21189 18785 21223 18819
rect 2329 18717 2363 18751
rect 4813 18717 4847 18751
rect 6929 18717 6963 18751
rect 9965 18717 9999 18751
rect 12081 18717 12115 18751
rect 13093 18717 13127 18751
rect 18521 18717 18555 18751
rect 7389 18649 7423 18683
rect 18245 18649 18279 18683
rect 21373 18649 21407 18683
rect 4261 18581 4295 18615
rect 8953 18581 8987 18615
rect 12633 18581 12667 18615
rect 15209 18581 15243 18615
rect 6653 18377 6687 18411
rect 6929 18377 6963 18411
rect 11713 18377 11747 18411
rect 19717 18377 19751 18411
rect 20361 18377 20395 18411
rect 20821 18377 20855 18411
rect 16957 18309 16991 18343
rect 7481 18241 7515 18275
rect 11161 18241 11195 18275
rect 13185 18241 13219 18275
rect 13369 18241 13403 18275
rect 15577 18241 15611 18275
rect 17325 18241 17359 18275
rect 18337 18241 18371 18275
rect 5273 18173 5307 18207
rect 7297 18173 7331 18207
rect 9321 18173 9355 18207
rect 9577 18173 9611 18207
rect 13461 18173 13495 18207
rect 15844 18173 15878 18207
rect 18613 18173 18647 18207
rect 20177 18173 20211 18207
rect 20637 18173 20671 18207
rect 5540 18105 5574 18139
rect 11345 18105 11379 18139
rect 11989 18105 12023 18139
rect 17509 18105 17543 18139
rect 21189 18105 21223 18139
rect 21373 18105 21407 18139
rect 7389 18037 7423 18071
rect 10701 18037 10735 18071
rect 11253 18037 11287 18071
rect 12725 18037 12759 18071
rect 13829 18037 13863 18071
rect 17601 18037 17635 18071
rect 17969 18037 18003 18071
rect 18521 18037 18555 18071
rect 18981 18037 19015 18071
rect 3617 17833 3651 17867
rect 5733 17833 5767 17867
rect 7573 17833 7607 17867
rect 9873 17833 9907 17867
rect 10333 17833 10367 17867
rect 18521 17833 18555 17867
rect 19349 17833 19383 17867
rect 20269 17833 20303 17867
rect 1777 17765 1811 17799
rect 17386 17765 17420 17799
rect 18797 17765 18831 17799
rect 3525 17697 3559 17731
rect 4261 17697 4295 17731
rect 7205 17697 7239 17731
rect 9965 17697 9999 17731
rect 10609 17697 10643 17731
rect 19165 17697 19199 17731
rect 19625 17697 19659 17731
rect 20085 17697 20119 17731
rect 20637 17697 20671 17731
rect 21189 17697 21223 17731
rect 3709 17629 3743 17663
rect 6929 17629 6963 17663
rect 7113 17629 7147 17663
rect 9781 17629 9815 17663
rect 17141 17629 17175 17663
rect 12173 17561 12207 17595
rect 19809 17561 19843 17595
rect 20821 17561 20855 17595
rect 21373 17561 21407 17595
rect 1685 17493 1719 17527
rect 3157 17493 3191 17527
rect 7849 17493 7883 17527
rect 1777 17289 1811 17323
rect 15485 17289 15519 17323
rect 19257 17289 19291 17323
rect 20637 17289 20671 17323
rect 4721 17221 4755 17255
rect 13001 17221 13035 17255
rect 7481 17153 7515 17187
rect 8493 17153 8527 17187
rect 11345 17153 11379 17187
rect 12449 17153 12483 17187
rect 14933 17153 14967 17187
rect 3157 17085 3191 17119
rect 4537 17085 4571 17119
rect 7665 17085 7699 17119
rect 7757 17085 7791 17119
rect 11529 17085 11563 17119
rect 11621 17085 11655 17119
rect 15117 17085 15151 17119
rect 19073 17085 19107 17119
rect 19809 17085 19843 17119
rect 20821 17085 20855 17119
rect 2912 17017 2946 17051
rect 15761 17017 15795 17051
rect 21189 17017 21223 17051
rect 21373 17017 21407 17051
rect 8125 16949 8159 16983
rect 11989 16949 12023 16983
rect 12541 16949 12575 16983
rect 12633 16949 12667 16983
rect 15025 16949 15059 16983
rect 19993 16949 20027 16983
rect 3065 16745 3099 16779
rect 3525 16745 3559 16779
rect 5917 16745 5951 16779
rect 9229 16745 9263 16779
rect 9689 16745 9723 16779
rect 10609 16745 10643 16779
rect 12173 16745 12207 16779
rect 14381 16745 14415 16779
rect 14841 16745 14875 16779
rect 18889 16745 18923 16779
rect 20361 16745 20395 16779
rect 20821 16745 20855 16779
rect 4804 16677 4838 16711
rect 7542 16677 7576 16711
rect 3157 16609 3191 16643
rect 3801 16609 3835 16643
rect 4537 16609 4571 16643
rect 7297 16609 7331 16643
rect 9321 16609 9355 16643
rect 9965 16609 9999 16643
rect 10425 16609 10459 16643
rect 12449 16609 12483 16643
rect 12705 16609 12739 16643
rect 14473 16609 14507 16643
rect 15209 16609 15243 16643
rect 15476 16609 15510 16643
rect 18705 16609 18739 16643
rect 19717 16609 19751 16643
rect 20177 16609 20211 16643
rect 20637 16609 20671 16643
rect 21189 16609 21223 16643
rect 21373 16609 21407 16643
rect 2881 16541 2915 16575
rect 9137 16541 9171 16575
rect 14289 16541 14323 16575
rect 8677 16473 8711 16507
rect 13829 16473 13863 16507
rect 16589 16405 16623 16439
rect 19901 16405 19935 16439
rect 4905 16201 4939 16235
rect 10701 16201 10735 16235
rect 12357 16201 12391 16235
rect 15945 16201 15979 16235
rect 17417 16201 17451 16235
rect 18521 16201 18555 16235
rect 20085 16201 20119 16235
rect 20821 16201 20855 16235
rect 6285 16065 6319 16099
rect 10977 16065 11011 16099
rect 14565 16065 14599 16099
rect 16497 16065 16531 16099
rect 17969 16065 18003 16099
rect 9321 15997 9355 16031
rect 9577 15997 9611 16031
rect 11244 15997 11278 16031
rect 19901 15997 19935 16031
rect 20637 15997 20671 16031
rect 6040 15929 6074 15963
rect 14810 15929 14844 15963
rect 16589 15929 16623 15963
rect 18061 15929 18095 15963
rect 21189 15929 21223 15963
rect 21373 15929 21407 15963
rect 16681 15861 16715 15895
rect 17049 15861 17083 15895
rect 18153 15861 18187 15895
rect 18797 15861 18831 15895
rect 3249 15657 3283 15691
rect 7849 15657 7883 15691
rect 18521 15657 18555 15691
rect 20821 15657 20855 15691
rect 8861 15589 8895 15623
rect 21189 15589 21223 15623
rect 1869 15521 1903 15555
rect 2136 15521 2170 15555
rect 7481 15521 7515 15555
rect 8125 15521 8159 15555
rect 8769 15521 8803 15555
rect 7205 15453 7239 15487
rect 7389 15453 7423 15487
rect 17397 15521 17431 15555
rect 19993 15521 20027 15555
rect 20637 15521 20671 15555
rect 17141 15453 17175 15487
rect 20177 15385 20211 15419
rect 21373 15385 21407 15419
rect 8585 15317 8619 15351
rect 8861 15317 8895 15351
rect 9137 15317 9171 15351
rect 14933 15317 14967 15351
rect 4813 15113 4847 15147
rect 6101 15113 6135 15147
rect 7757 15113 7791 15147
rect 14749 15113 14783 15147
rect 20361 15113 20395 15147
rect 4169 14977 4203 15011
rect 8217 14977 8251 15011
rect 8309 14977 8343 15011
rect 12541 14977 12575 15011
rect 17785 14977 17819 15011
rect 7481 14909 7515 14943
rect 9505 14909 9539 14943
rect 14565 14909 14599 14943
rect 20177 14909 20211 14943
rect 20637 14909 20671 14943
rect 4445 14841 4479 14875
rect 5089 14841 5123 14875
rect 7214 14841 7248 14875
rect 18030 14841 18064 14875
rect 21189 14841 21223 14875
rect 21373 14841 21407 14875
rect 4353 14773 4387 14807
rect 8125 14773 8159 14807
rect 9321 14773 9355 14807
rect 12633 14773 12667 14807
rect 12725 14773 12759 14807
rect 13093 14773 13127 14807
rect 19165 14773 19199 14807
rect 20821 14773 20855 14807
rect 2513 14569 2547 14603
rect 4261 14569 4295 14603
rect 4721 14569 4755 14603
rect 8585 14569 8619 14603
rect 9689 14569 9723 14603
rect 12173 14569 12207 14603
rect 12633 14569 12667 14603
rect 15577 14569 15611 14603
rect 17969 14569 18003 14603
rect 18429 14569 18463 14603
rect 18981 14569 19015 14603
rect 20821 14569 20855 14603
rect 4629 14501 4663 14535
rect 5365 14501 5399 14535
rect 3637 14433 3671 14467
rect 8677 14433 8711 14467
rect 9505 14433 9539 14467
rect 12265 14433 12299 14467
rect 12817 14433 12851 14467
rect 14758 14433 14792 14467
rect 15025 14433 15059 14467
rect 15669 14433 15703 14467
rect 18061 14433 18095 14467
rect 19073 14433 19107 14467
rect 19993 14433 20027 14467
rect 20637 14433 20671 14467
rect 21097 14433 21131 14467
rect 3893 14365 3927 14399
rect 4813 14365 4847 14399
rect 8493 14365 8527 14399
rect 9965 14365 9999 14399
rect 12081 14365 12115 14399
rect 15393 14365 15427 14399
rect 17877 14365 17911 14399
rect 18797 14365 18831 14399
rect 19441 14297 19475 14331
rect 20177 14297 20211 14331
rect 21281 14297 21315 14331
rect 9045 14229 9079 14263
rect 12817 14229 12851 14263
rect 13001 14229 13035 14263
rect 13645 14229 13679 14263
rect 16037 14229 16071 14263
rect 4169 14025 4203 14059
rect 7297 14025 7331 14059
rect 11069 14025 11103 14059
rect 14013 14025 14047 14059
rect 15669 14025 15703 14059
rect 16589 14025 16623 14059
rect 15025 13889 15059 13923
rect 17325 13889 17359 13923
rect 21373 13889 21407 13923
rect 5293 13821 5327 13855
rect 5549 13821 5583 13855
rect 8677 13821 8711 13855
rect 12357 13821 12391 13855
rect 12633 13821 12667 13855
rect 12889 13821 12923 13855
rect 16405 13821 16439 13855
rect 17592 13821 17626 13855
rect 19625 13821 19659 13855
rect 20361 13821 20395 13855
rect 20821 13821 20855 13855
rect 8432 13753 8466 13787
rect 18981 13753 19015 13787
rect 21189 13753 21223 13787
rect 15209 13685 15243 13719
rect 15301 13685 15335 13719
rect 15945 13685 15979 13719
rect 18705 13685 18739 13719
rect 20637 13685 20671 13719
rect 6653 13481 6687 13515
rect 8861 13481 8895 13515
rect 9321 13481 9355 13515
rect 12541 13481 12575 13515
rect 13001 13481 13035 13515
rect 13461 13481 13495 13515
rect 15853 13481 15887 13515
rect 18889 13481 18923 13515
rect 19349 13481 19383 13515
rect 20361 13481 20395 13515
rect 7788 13413 7822 13447
rect 21373 13413 21407 13447
rect 8953 13345 8987 13379
rect 10721 13345 10755 13379
rect 12633 13345 12667 13379
rect 13277 13345 13311 13379
rect 18981 13345 19015 13379
rect 19625 13345 19659 13379
rect 20177 13345 20211 13379
rect 20821 13345 20855 13379
rect 21189 13345 21223 13379
rect 8033 13277 8067 13311
rect 8677 13277 8711 13311
rect 10977 13277 11011 13311
rect 12357 13277 12391 13311
rect 14105 13277 14139 13311
rect 18705 13277 18739 13311
rect 20637 13209 20671 13243
rect 9597 13141 9631 13175
rect 13737 13141 13771 13175
rect 17049 13141 17083 13175
rect 9781 12937 9815 12971
rect 12173 12937 12207 12971
rect 13829 12937 13863 12971
rect 19993 12937 20027 12971
rect 20913 12937 20947 12971
rect 21189 12937 21223 12971
rect 20453 12869 20487 12903
rect 10333 12801 10367 12835
rect 16405 12801 16439 12835
rect 16589 12801 16623 12835
rect 17049 12801 17083 12835
rect 17233 12801 17267 12835
rect 10793 12733 10827 12767
rect 13645 12733 13679 12767
rect 16313 12733 16347 12767
rect 19257 12733 19291 12767
rect 19809 12733 19843 12767
rect 20269 12733 20303 12767
rect 20729 12733 20763 12767
rect 21373 12733 21407 12767
rect 10149 12665 10183 12699
rect 11060 12665 11094 12699
rect 10241 12597 10275 12631
rect 15945 12597 15979 12631
rect 17325 12597 17359 12631
rect 17693 12597 17727 12631
rect 10701 12393 10735 12427
rect 11069 12393 11103 12427
rect 12081 12393 12115 12427
rect 16129 12393 16163 12427
rect 16589 12393 16623 12427
rect 17141 12393 17175 12427
rect 19533 12393 19567 12427
rect 20361 12393 20395 12427
rect 20821 12393 20855 12427
rect 14228 12325 14262 12359
rect 16221 12325 16255 12359
rect 8677 12257 8711 12291
rect 11897 12257 11931 12291
rect 14473 12257 14507 12291
rect 17509 12257 17543 12291
rect 19073 12257 19107 12291
rect 19349 12257 19383 12291
rect 19809 12257 19843 12291
rect 20545 12257 20579 12291
rect 21005 12257 21039 12291
rect 15945 12189 15979 12223
rect 17601 12189 17635 12223
rect 17785 12189 17819 12223
rect 18153 12121 18187 12155
rect 19993 12121 20027 12155
rect 8493 12053 8527 12087
rect 13093 12053 13127 12087
rect 18613 12053 18647 12087
rect 21373 12053 21407 12087
rect 11713 11849 11747 11883
rect 14841 11849 14875 11883
rect 17417 11849 17451 11883
rect 19073 11849 19107 11883
rect 20085 11849 20119 11883
rect 20821 11849 20855 11883
rect 10701 11781 10735 11815
rect 20545 11781 20579 11815
rect 11069 11713 11103 11747
rect 13737 11713 13771 11747
rect 17969 11713 18003 11747
rect 9321 11645 9355 11679
rect 15965 11645 15999 11679
rect 16221 11645 16255 11679
rect 19257 11645 19291 11679
rect 19901 11645 19935 11679
rect 20361 11645 20395 11679
rect 21005 11645 21039 11679
rect 21097 11645 21131 11679
rect 9566 11577 9600 11611
rect 12909 11577 12943 11611
rect 13645 11577 13679 11611
rect 17785 11577 17819 11611
rect 18429 11577 18463 11611
rect 11253 11509 11287 11543
rect 11345 11509 11379 11543
rect 13185 11509 13219 11543
rect 13553 11509 13587 11543
rect 14473 11509 14507 11543
rect 17877 11509 17911 11543
rect 21097 11509 21131 11543
rect 21373 11509 21407 11543
rect 8769 11305 8803 11339
rect 9321 11305 9355 11339
rect 9781 11305 9815 11339
rect 11161 11305 11195 11339
rect 13921 11305 13955 11339
rect 18061 11305 18095 11339
rect 19073 11305 19107 11339
rect 20085 11305 20119 11339
rect 20821 11305 20855 11339
rect 8309 11237 8343 11271
rect 10149 11237 10183 11271
rect 18521 11237 18555 11271
rect 8401 11169 8435 11203
rect 9413 11169 9447 11203
rect 10793 11169 10827 11203
rect 13553 11169 13587 11203
rect 14565 11169 14599 11203
rect 17785 11169 17819 11203
rect 18429 11169 18463 11203
rect 19257 11169 19291 11203
rect 19901 11169 19935 11203
rect 20545 11169 20579 11203
rect 21005 11169 21039 11203
rect 8217 11101 8251 11135
rect 9229 11101 9263 11135
rect 10517 11101 10551 11135
rect 10701 11101 10735 11135
rect 13277 11101 13311 11135
rect 13461 11101 13495 11135
rect 18613 11101 18647 11135
rect 19625 11101 19659 11135
rect 20361 11033 20395 11067
rect 21373 11033 21407 11067
rect 14749 10965 14783 10999
rect 8769 10761 8803 10795
rect 11069 10761 11103 10795
rect 11897 10761 11931 10795
rect 13737 10761 13771 10795
rect 16129 10761 16163 10795
rect 19809 10761 19843 10795
rect 10057 10693 10091 10727
rect 8217 10625 8251 10659
rect 8401 10557 8435 10591
rect 9873 10557 9907 10591
rect 10793 10625 10827 10659
rect 11621 10625 11655 10659
rect 12541 10693 12575 10727
rect 17693 10693 17727 10727
rect 17877 10693 17911 10727
rect 20821 10693 20855 10727
rect 13093 10625 13127 10659
rect 13277 10625 13311 10659
rect 17509 10557 17543 10591
rect 20361 10625 20395 10659
rect 18337 10557 18371 10591
rect 21005 10557 21039 10591
rect 8309 10489 8343 10523
rect 10057 10489 10091 10523
rect 10149 10489 10183 10523
rect 11437 10489 11471 10523
rect 11897 10489 11931 10523
rect 17264 10489 17298 10523
rect 17693 10489 17727 10523
rect 20177 10489 20211 10523
rect 9413 10421 9447 10455
rect 11529 10421 11563 10455
rect 12081 10421 12115 10455
rect 13369 10421 13403 10455
rect 14473 10421 14507 10455
rect 18981 10421 19015 10455
rect 20269 10421 20303 10455
rect 9965 10217 9999 10251
rect 13093 10217 13127 10251
rect 13553 10217 13587 10251
rect 20453 10217 20487 10251
rect 20913 10217 20947 10251
rect 8300 10149 8334 10183
rect 11100 10149 11134 10183
rect 13461 10149 13495 10183
rect 8033 10081 8067 10115
rect 11345 10081 11379 10115
rect 14361 10081 14395 10115
rect 18797 10081 18831 10115
rect 19064 10081 19098 10115
rect 21097 10081 21131 10115
rect 13645 10013 13679 10047
rect 14105 10013 14139 10047
rect 9413 9945 9447 9979
rect 15485 9877 15519 9911
rect 20177 9877 20211 9911
rect 9137 9673 9171 9707
rect 11805 9673 11839 9707
rect 13921 9673 13955 9707
rect 17233 9673 17267 9707
rect 19809 9673 19843 9707
rect 14841 9605 14875 9639
rect 20821 9605 20855 9639
rect 22017 9605 22051 9639
rect 15393 9537 15427 9571
rect 20361 9537 20395 9571
rect 12918 9469 12952 9503
rect 13185 9469 13219 9503
rect 13461 9469 13495 9503
rect 18613 9469 18647 9503
rect 21005 9469 21039 9503
rect 15209 9401 15243 9435
rect 15853 9401 15887 9435
rect 18368 9401 18402 9435
rect 20177 9401 20211 9435
rect 14473 9333 14507 9367
rect 15301 9333 15335 9367
rect 16405 9333 16439 9367
rect 19257 9333 19291 9367
rect 20269 9333 20303 9367
rect 12081 9129 12115 9163
rect 15761 9129 15795 9163
rect 20085 9129 20119 9163
rect 20545 9129 20579 9163
rect 11897 8993 11931 9027
rect 15945 8993 15979 9027
rect 19625 8993 19659 9027
rect 19901 8993 19935 9027
rect 20361 8993 20395 9027
rect 21005 8993 21039 9027
rect 21373 8925 21407 8959
rect 20821 8857 20855 8891
rect 11437 8585 11471 8619
rect 13277 8585 13311 8619
rect 16221 8585 16255 8619
rect 20085 8585 20119 8619
rect 21373 8585 21407 8619
rect 22017 8585 22051 8619
rect 13737 8517 13771 8551
rect 14565 8517 14599 8551
rect 20545 8517 20579 8551
rect 15117 8449 15151 8483
rect 11253 8381 11287 8415
rect 13461 8381 13495 8415
rect 13921 8381 13955 8415
rect 16405 8381 16439 8415
rect 19257 8381 19291 8415
rect 19901 8381 19935 8415
rect 20361 8381 20395 8415
rect 21005 8381 21039 8415
rect 15025 8313 15059 8347
rect 14933 8245 14967 8279
rect 17509 8245 17543 8279
rect 20821 8245 20855 8279
rect 11897 8041 11931 8075
rect 17141 8041 17175 8075
rect 17509 8041 17543 8075
rect 19625 8041 19659 8075
rect 20085 8041 20119 8075
rect 20545 8041 20579 8075
rect 12265 7905 12299 7939
rect 13645 7905 13679 7939
rect 13912 7905 13946 7939
rect 18501 7905 18535 7939
rect 19901 7905 19935 7939
rect 20361 7905 20395 7939
rect 21005 7905 21039 7939
rect 12357 7837 12391 7871
rect 12449 7837 12483 7871
rect 17601 7837 17635 7871
rect 17785 7837 17819 7871
rect 18245 7837 18279 7871
rect 15025 7701 15059 7735
rect 20821 7701 20855 7735
rect 21373 7701 21407 7735
rect 18429 7497 18463 7531
rect 19993 7497 20027 7531
rect 20821 7497 20855 7531
rect 20545 7429 20579 7463
rect 11621 7361 11655 7395
rect 14749 7361 14783 7395
rect 9689 7293 9723 7327
rect 11897 7293 11931 7327
rect 15393 7293 15427 7327
rect 17049 7293 17083 7327
rect 20361 7293 20395 7327
rect 21005 7293 21039 7327
rect 9956 7225 9990 7259
rect 12142 7225 12176 7259
rect 15638 7225 15672 7259
rect 17316 7225 17350 7259
rect 11069 7157 11103 7191
rect 13277 7157 13311 7191
rect 16773 7157 16807 7191
rect 21373 7157 21407 7191
rect 11897 6953 11931 6987
rect 12265 6953 12299 6987
rect 17693 6953 17727 6987
rect 18061 6953 18095 6987
rect 20361 6953 20395 6987
rect 14841 6885 14875 6919
rect 8473 6817 8507 6851
rect 11345 6817 11379 6851
rect 12357 6817 12391 6851
rect 14197 6817 14231 6851
rect 14749 6817 14783 6851
rect 17417 6817 17451 6851
rect 18153 6817 18187 6851
rect 20085 6817 20119 6851
rect 20545 6817 20579 6851
rect 21005 6817 21039 6851
rect 8217 6749 8251 6783
rect 12449 6749 12483 6783
rect 14565 6749 14599 6783
rect 18245 6749 18279 6783
rect 9597 6681 9631 6715
rect 15209 6681 15243 6715
rect 20821 6613 20855 6647
rect 21373 6613 21407 6647
rect 20913 6409 20947 6443
rect 21189 6341 21223 6375
rect 20453 6205 20487 6239
rect 20729 6205 20763 6239
rect 21373 6205 21407 6239
rect 1777 5865 1811 5899
rect 20821 5797 20855 5831
rect 1593 5729 1627 5763
rect 2053 5729 2087 5763
rect 21005 5729 21039 5763
rect 20913 5321 20947 5355
rect 21189 5321 21223 5355
rect 20453 5117 20487 5151
rect 20729 5117 20763 5151
rect 21373 5117 21407 5151
rect 20821 4777 20855 4811
rect 21373 4709 21407 4743
rect 21005 4641 21039 4675
rect 20821 4233 20855 4267
rect 21097 4097 21131 4131
rect 20361 4029 20395 4063
rect 20637 4029 20671 4063
rect 19993 3961 20027 3995
rect 21281 3961 21315 3995
rect 20637 3689 20671 3723
rect 21097 3621 21131 3655
rect 19349 3553 19383 3587
rect 20729 3553 20763 3587
rect 21281 3553 21315 3587
rect 20269 3485 20303 3519
rect 19625 3349 19659 3383
rect 20637 3145 20671 3179
rect 19993 3077 20027 3111
rect 19257 3009 19291 3043
rect 20913 3009 20947 3043
rect 19717 2941 19751 2975
rect 18889 2873 18923 2907
rect 20177 2873 20211 2907
rect 20729 2873 20763 2907
rect 20913 2873 20947 2907
rect 21281 2873 21315 2907
rect 21189 2805 21223 2839
rect 20637 2601 20671 2635
rect 18981 2533 19015 2567
rect 20729 2533 20763 2567
rect 22017 2533 22051 2567
rect 19257 2465 19291 2499
rect 19441 2465 19475 2499
rect 21281 2465 21315 2499
rect 20269 2397 20303 2431
rect 21097 2329 21131 2363
rect 22017 1377 22051 1411
<< metal1 >>
rect 3050 20816 3056 20868
rect 3108 20856 3114 20868
rect 4246 20856 4252 20868
rect 3108 20828 4252 20856
rect 3108 20816 3114 20828
rect 4246 20816 4252 20828
rect 4304 20816 4310 20868
rect 4706 20816 4712 20868
rect 4764 20856 4770 20868
rect 5442 20856 5448 20868
rect 4764 20828 5448 20856
rect 4764 20816 4770 20828
rect 5442 20816 5448 20828
rect 5500 20816 5506 20868
rect 4154 20748 4160 20800
rect 4212 20788 4218 20800
rect 5534 20788 5540 20800
rect 4212 20760 5540 20788
rect 4212 20748 4218 20760
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 2777 20587 2835 20593
rect 2777 20553 2789 20587
rect 2823 20584 2835 20587
rect 6730 20584 6736 20596
rect 2823 20556 6736 20584
rect 2823 20553 2835 20556
rect 2777 20547 2835 20553
rect 6730 20544 6736 20556
rect 6788 20544 6794 20596
rect 6914 20544 6920 20596
rect 6972 20584 6978 20596
rect 8846 20584 8852 20596
rect 6972 20556 8852 20584
rect 6972 20544 6978 20556
rect 8846 20544 8852 20556
rect 8904 20544 8910 20596
rect 11425 20587 11483 20593
rect 11425 20553 11437 20587
rect 11471 20584 11483 20587
rect 14274 20584 14280 20596
rect 11471 20556 14280 20584
rect 11471 20553 11483 20556
rect 11425 20547 11483 20553
rect 14274 20544 14280 20556
rect 14332 20544 14338 20596
rect 16209 20587 16267 20593
rect 16209 20553 16221 20587
rect 16255 20584 16267 20587
rect 18138 20584 18144 20596
rect 16255 20556 18144 20584
rect 16255 20553 16267 20556
rect 16209 20547 16267 20553
rect 18138 20544 18144 20556
rect 18196 20544 18202 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 20990 20584 20996 20596
rect 19484 20556 20996 20584
rect 19484 20544 19490 20556
rect 20990 20544 20996 20556
rect 21048 20544 21054 20596
rect 1394 20476 1400 20528
rect 1452 20516 1458 20528
rect 1452 20488 2636 20516
rect 1452 20476 1458 20488
rect 842 20408 848 20460
rect 900 20448 906 20460
rect 900 20420 2176 20448
rect 900 20408 906 20420
rect 290 20340 296 20392
rect 348 20380 354 20392
rect 1302 20380 1308 20392
rect 348 20352 1308 20380
rect 348 20340 354 20352
rect 1302 20340 1308 20352
rect 1360 20380 1366 20392
rect 1673 20383 1731 20389
rect 1673 20380 1685 20383
rect 1360 20352 1685 20380
rect 1360 20340 1366 20352
rect 1673 20349 1685 20352
rect 1719 20349 1731 20383
rect 1673 20343 1731 20349
rect 2038 20340 2044 20392
rect 2096 20380 2102 20392
rect 2148 20389 2176 20420
rect 2133 20383 2191 20389
rect 2133 20380 2145 20383
rect 2096 20352 2145 20380
rect 2096 20340 2102 20352
rect 2133 20349 2145 20352
rect 2179 20349 2191 20383
rect 2133 20343 2191 20349
rect 2498 20340 2504 20392
rect 2556 20380 2562 20392
rect 2608 20389 2636 20488
rect 3602 20476 3608 20528
rect 3660 20516 3666 20528
rect 4985 20519 5043 20525
rect 4985 20516 4997 20519
rect 3660 20488 4997 20516
rect 3660 20476 3666 20488
rect 4985 20485 4997 20488
rect 5031 20485 5043 20519
rect 4985 20479 5043 20485
rect 5166 20476 5172 20528
rect 5224 20516 5230 20528
rect 7742 20516 7748 20528
rect 5224 20488 7748 20516
rect 5224 20476 5230 20488
rect 7742 20476 7748 20488
rect 7800 20476 7806 20528
rect 7837 20519 7895 20525
rect 7837 20485 7849 20519
rect 7883 20516 7895 20519
rect 8202 20516 8208 20528
rect 7883 20488 8208 20516
rect 7883 20485 7895 20488
rect 7837 20479 7895 20485
rect 8202 20476 8208 20488
rect 8260 20476 8266 20528
rect 10045 20519 10103 20525
rect 10045 20485 10057 20519
rect 10091 20516 10103 20519
rect 11790 20516 11796 20528
rect 10091 20488 11796 20516
rect 10091 20485 10103 20488
rect 10045 20479 10103 20485
rect 11790 20476 11796 20488
rect 11848 20476 11854 20528
rect 12066 20516 12072 20528
rect 12027 20488 12072 20516
rect 12066 20476 12072 20488
rect 12124 20476 12130 20528
rect 12618 20516 12624 20528
rect 12579 20488 12624 20516
rect 12618 20476 12624 20488
rect 12676 20476 12682 20528
rect 13170 20516 13176 20528
rect 13131 20488 13176 20516
rect 13170 20476 13176 20488
rect 13228 20476 13234 20528
rect 13722 20516 13728 20528
rect 13683 20488 13728 20516
rect 13722 20476 13728 20488
rect 13780 20476 13786 20528
rect 16853 20519 16911 20525
rect 16853 20485 16865 20519
rect 16899 20516 16911 20519
rect 17678 20516 17684 20528
rect 16899 20488 17684 20516
rect 16899 20485 16911 20488
rect 16853 20479 16911 20485
rect 17678 20476 17684 20488
rect 17736 20476 17742 20528
rect 17865 20519 17923 20525
rect 17865 20485 17877 20519
rect 17911 20516 17923 20519
rect 17954 20516 17960 20528
rect 17911 20488 17960 20516
rect 17911 20485 17923 20488
rect 17865 20479 17923 20485
rect 17954 20476 17960 20488
rect 18012 20476 18018 20528
rect 18417 20519 18475 20525
rect 18417 20485 18429 20519
rect 18463 20516 18475 20519
rect 18598 20516 18604 20528
rect 18463 20488 18604 20516
rect 18463 20485 18475 20488
rect 18417 20479 18475 20485
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 18782 20476 18788 20528
rect 18840 20476 18846 20528
rect 18966 20516 18972 20528
rect 18927 20488 18972 20516
rect 18966 20476 18972 20488
rect 19024 20476 19030 20528
rect 19518 20516 19524 20528
rect 19479 20488 19524 20516
rect 19518 20476 19524 20488
rect 19576 20476 19582 20528
rect 2774 20408 2780 20460
rect 2832 20448 2838 20460
rect 3786 20448 3792 20460
rect 2832 20420 3792 20448
rect 2832 20408 2838 20420
rect 3786 20408 3792 20420
rect 3844 20448 3850 20460
rect 3844 20420 4108 20448
rect 3844 20408 3850 20420
rect 4080 20389 4108 20420
rect 4154 20408 4160 20460
rect 4212 20448 4218 20460
rect 4212 20420 5212 20448
rect 4212 20408 4218 20420
rect 2593 20383 2651 20389
rect 2593 20380 2605 20383
rect 2556 20352 2605 20380
rect 2556 20340 2562 20352
rect 2593 20349 2605 20352
rect 2639 20349 2651 20383
rect 2593 20343 2651 20349
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20349 3111 20383
rect 3053 20343 3111 20349
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20349 4123 20383
rect 4065 20343 4123 20349
rect 1946 20272 1952 20324
rect 2004 20312 2010 20324
rect 2866 20312 2872 20324
rect 2004 20284 2872 20312
rect 2004 20272 2010 20284
rect 2866 20272 2872 20284
rect 2924 20312 2930 20324
rect 3068 20312 3096 20343
rect 4246 20340 4252 20392
rect 4304 20380 4310 20392
rect 4525 20383 4583 20389
rect 4525 20380 4537 20383
rect 4304 20352 4537 20380
rect 4304 20340 4310 20352
rect 4525 20349 4537 20352
rect 4571 20380 4583 20383
rect 5074 20380 5080 20392
rect 4571 20352 5080 20380
rect 4571 20349 4583 20352
rect 4525 20343 4583 20349
rect 5074 20340 5080 20352
rect 5132 20340 5138 20392
rect 5184 20389 5212 20420
rect 5442 20408 5448 20460
rect 5500 20448 5506 20460
rect 5500 20420 5948 20448
rect 5500 20408 5506 20420
rect 5169 20383 5227 20389
rect 5169 20349 5181 20383
rect 5215 20380 5227 20383
rect 5350 20380 5356 20392
rect 5215 20352 5356 20380
rect 5215 20349 5227 20352
rect 5169 20343 5227 20349
rect 5350 20340 5356 20352
rect 5408 20340 5414 20392
rect 5534 20340 5540 20392
rect 5592 20380 5598 20392
rect 5920 20389 5948 20420
rect 6822 20408 6828 20460
rect 6880 20448 6886 20460
rect 7009 20451 7067 20457
rect 6880 20408 6914 20448
rect 7009 20417 7021 20451
rect 7055 20448 7067 20451
rect 12250 20448 12256 20460
rect 7055 20420 12256 20448
rect 7055 20417 7067 20420
rect 7009 20411 7067 20417
rect 12250 20408 12256 20420
rect 12308 20408 12314 20460
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20448 15807 20451
rect 18800 20448 18828 20476
rect 15795 20420 18828 20448
rect 15795 20417 15807 20420
rect 15749 20411 15807 20417
rect 6886 20392 6914 20408
rect 5629 20383 5687 20389
rect 5629 20380 5641 20383
rect 5592 20352 5641 20380
rect 5592 20340 5598 20352
rect 5629 20349 5641 20352
rect 5675 20349 5687 20383
rect 5629 20343 5687 20349
rect 5905 20383 5963 20389
rect 5905 20349 5917 20383
rect 5951 20349 5963 20383
rect 5905 20343 5963 20349
rect 6454 20340 6460 20392
rect 6512 20380 6518 20392
rect 6733 20383 6791 20389
rect 6733 20380 6745 20383
rect 6512 20352 6745 20380
rect 6512 20340 6518 20352
rect 6733 20349 6745 20352
rect 6779 20349 6791 20383
rect 6886 20352 6920 20392
rect 6733 20343 6791 20349
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 7193 20383 7251 20389
rect 7193 20380 7205 20383
rect 7156 20352 7205 20380
rect 7156 20340 7162 20352
rect 7193 20349 7205 20352
rect 7239 20349 7251 20383
rect 7193 20343 7251 20349
rect 7558 20340 7564 20392
rect 7616 20380 7622 20392
rect 7653 20383 7711 20389
rect 7653 20380 7665 20383
rect 7616 20352 7665 20380
rect 7616 20340 7622 20352
rect 7653 20349 7665 20352
rect 7699 20349 7711 20383
rect 8294 20380 8300 20392
rect 8255 20352 8300 20380
rect 7653 20343 7711 20349
rect 8294 20340 8300 20352
rect 8352 20340 8358 20392
rect 8662 20340 8668 20392
rect 8720 20380 8726 20392
rect 8849 20383 8907 20389
rect 8849 20380 8861 20383
rect 8720 20352 8861 20380
rect 8720 20340 8726 20352
rect 8849 20349 8861 20352
rect 8895 20380 8907 20383
rect 9122 20380 9128 20392
rect 8895 20352 9128 20380
rect 8895 20349 8907 20352
rect 8849 20343 8907 20349
rect 9122 20340 9128 20352
rect 9180 20340 9186 20392
rect 9214 20340 9220 20392
rect 9272 20380 9278 20392
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 9272 20352 9413 20380
rect 9272 20340 9278 20352
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 9766 20340 9772 20392
rect 9824 20380 9830 20392
rect 9861 20383 9919 20389
rect 9861 20380 9873 20383
rect 9824 20352 9873 20380
rect 9824 20340 9830 20352
rect 9861 20349 9873 20352
rect 9907 20349 9919 20383
rect 10318 20380 10324 20392
rect 10279 20352 10324 20380
rect 9861 20343 9919 20349
rect 10318 20340 10324 20352
rect 10376 20340 10382 20392
rect 10781 20383 10839 20389
rect 10781 20349 10793 20383
rect 10827 20380 10839 20383
rect 10870 20380 10876 20392
rect 10827 20352 10876 20380
rect 10827 20349 10839 20352
rect 10781 20343 10839 20349
rect 10870 20340 10876 20352
rect 10928 20340 10934 20392
rect 15013 20383 15071 20389
rect 15013 20349 15025 20383
rect 15059 20380 15071 20383
rect 15838 20380 15844 20392
rect 15059 20352 15844 20380
rect 15059 20349 15071 20352
rect 15013 20343 15071 20349
rect 15838 20340 15844 20352
rect 15896 20340 15902 20392
rect 16117 20383 16175 20389
rect 16117 20349 16129 20383
rect 16163 20380 16175 20383
rect 16206 20380 16212 20392
rect 16163 20352 16212 20380
rect 16163 20349 16175 20352
rect 16117 20343 16175 20349
rect 16206 20340 16212 20352
rect 16264 20340 16270 20392
rect 18785 20383 18843 20389
rect 16592 20352 18736 20380
rect 7009 20315 7067 20321
rect 7009 20312 7021 20315
rect 2924 20284 3096 20312
rect 3252 20284 7021 20312
rect 2924 20272 2930 20284
rect 1762 20244 1768 20256
rect 1723 20216 1768 20244
rect 1762 20204 1768 20216
rect 1820 20204 1826 20256
rect 2314 20244 2320 20256
rect 2275 20216 2320 20244
rect 2314 20204 2320 20216
rect 2372 20204 2378 20256
rect 3252 20253 3280 20284
rect 7009 20281 7021 20284
rect 7055 20281 7067 20315
rect 11238 20312 11244 20324
rect 7009 20275 7067 20281
rect 7300 20284 11244 20312
rect 3237 20247 3295 20253
rect 3237 20213 3249 20247
rect 3283 20213 3295 20247
rect 3237 20207 3295 20213
rect 4249 20247 4307 20253
rect 4249 20213 4261 20247
rect 4295 20244 4307 20247
rect 4614 20244 4620 20256
rect 4295 20216 4620 20244
rect 4295 20213 4307 20216
rect 4249 20207 4307 20213
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 4709 20247 4767 20253
rect 4709 20213 4721 20247
rect 4755 20244 4767 20247
rect 4890 20244 4896 20256
rect 4755 20216 4896 20244
rect 4755 20213 4767 20216
rect 4709 20207 4767 20213
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 5442 20244 5448 20256
rect 5403 20216 5448 20244
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 6086 20244 6092 20256
rect 6047 20216 6092 20244
rect 6086 20204 6092 20216
rect 6144 20204 6150 20256
rect 6917 20247 6975 20253
rect 6917 20213 6929 20247
rect 6963 20244 6975 20247
rect 7300 20244 7328 20284
rect 11238 20272 11244 20284
rect 11296 20272 11302 20324
rect 11333 20315 11391 20321
rect 11333 20281 11345 20315
rect 11379 20312 11391 20315
rect 11882 20312 11888 20324
rect 11379 20284 11888 20312
rect 11379 20281 11391 20284
rect 11333 20275 11391 20281
rect 11882 20272 11888 20284
rect 11940 20272 11946 20324
rect 12158 20272 12164 20324
rect 12216 20312 12222 20324
rect 12253 20315 12311 20321
rect 12253 20312 12265 20315
rect 12216 20284 12265 20312
rect 12216 20272 12222 20284
rect 12253 20281 12265 20284
rect 12299 20281 12311 20315
rect 12253 20275 12311 20281
rect 12805 20315 12863 20321
rect 12805 20281 12817 20315
rect 12851 20312 12863 20315
rect 12894 20312 12900 20324
rect 12851 20284 12900 20312
rect 12851 20281 12863 20284
rect 12805 20275 12863 20281
rect 12894 20272 12900 20284
rect 12952 20272 12958 20324
rect 13262 20272 13268 20324
rect 13320 20312 13326 20324
rect 13357 20315 13415 20321
rect 13357 20312 13369 20315
rect 13320 20284 13369 20312
rect 13320 20272 13326 20284
rect 13357 20281 13369 20284
rect 13403 20281 13415 20315
rect 13357 20275 13415 20281
rect 13909 20315 13967 20321
rect 13909 20281 13921 20315
rect 13955 20312 13967 20315
rect 15197 20315 15255 20321
rect 13955 20284 14412 20312
rect 13955 20281 13967 20284
rect 13909 20275 13967 20281
rect 14384 20256 14412 20284
rect 15197 20281 15209 20315
rect 15243 20281 15255 20315
rect 15197 20275 15255 20281
rect 15565 20315 15623 20321
rect 15565 20281 15577 20315
rect 15611 20312 15623 20315
rect 16592 20312 16620 20352
rect 15611 20284 16620 20312
rect 16669 20315 16727 20321
rect 15611 20281 15623 20284
rect 15565 20275 15623 20281
rect 16669 20281 16681 20315
rect 16715 20312 16727 20315
rect 17586 20312 17592 20324
rect 16715 20284 17592 20312
rect 16715 20281 16727 20284
rect 16669 20275 16727 20281
rect 6963 20216 7328 20244
rect 7377 20247 7435 20253
rect 6963 20213 6975 20216
rect 6917 20207 6975 20213
rect 7377 20213 7389 20247
rect 7423 20244 7435 20247
rect 7466 20244 7472 20256
rect 7423 20216 7472 20244
rect 7423 20213 7435 20216
rect 7377 20207 7435 20213
rect 7466 20204 7472 20216
rect 7524 20204 7530 20256
rect 7650 20204 7656 20256
rect 7708 20244 7714 20256
rect 8113 20247 8171 20253
rect 8113 20244 8125 20247
rect 7708 20216 8125 20244
rect 7708 20204 7714 20216
rect 8113 20213 8125 20216
rect 8159 20213 8171 20247
rect 8662 20244 8668 20256
rect 8623 20216 8668 20244
rect 8113 20207 8171 20213
rect 8662 20204 8668 20216
rect 8720 20204 8726 20256
rect 9582 20244 9588 20256
rect 9543 20216 9588 20244
rect 9582 20204 9588 20216
rect 9640 20204 9646 20256
rect 10505 20247 10563 20253
rect 10505 20213 10517 20247
rect 10551 20244 10563 20247
rect 10870 20244 10876 20256
rect 10551 20216 10876 20244
rect 10551 20213 10563 20216
rect 10505 20207 10563 20213
rect 10870 20204 10876 20216
rect 10928 20204 10934 20256
rect 10965 20247 11023 20253
rect 10965 20213 10977 20247
rect 11011 20244 11023 20247
rect 14182 20244 14188 20256
rect 11011 20216 14188 20244
rect 11011 20213 11023 20216
rect 10965 20207 11023 20213
rect 14182 20204 14188 20216
rect 14240 20204 14246 20256
rect 14366 20204 14372 20256
rect 14424 20244 14430 20256
rect 14553 20247 14611 20253
rect 14553 20244 14565 20247
rect 14424 20216 14565 20244
rect 14424 20204 14430 20216
rect 14553 20213 14565 20216
rect 14599 20213 14611 20247
rect 15212 20244 15240 20275
rect 17586 20272 17592 20284
rect 17644 20272 17650 20324
rect 17681 20315 17739 20321
rect 17681 20281 17693 20315
rect 17727 20312 17739 20315
rect 18138 20312 18144 20324
rect 17727 20284 18144 20312
rect 17727 20281 17739 20284
rect 17681 20275 17739 20281
rect 18138 20272 18144 20284
rect 18196 20272 18202 20324
rect 18233 20315 18291 20321
rect 18233 20281 18245 20315
rect 18279 20312 18291 20315
rect 18598 20312 18604 20324
rect 18279 20284 18604 20312
rect 18279 20281 18291 20284
rect 18233 20275 18291 20281
rect 18598 20272 18604 20284
rect 18656 20272 18662 20324
rect 18708 20312 18736 20352
rect 18785 20349 18797 20383
rect 18831 20380 18843 20383
rect 19518 20380 19524 20392
rect 18831 20352 19524 20380
rect 18831 20349 18843 20352
rect 18785 20343 18843 20349
rect 19518 20340 19524 20352
rect 19576 20340 19582 20392
rect 20254 20380 20260 20392
rect 20215 20352 20260 20380
rect 20254 20340 20260 20352
rect 20312 20340 20318 20392
rect 20530 20340 20536 20392
rect 20588 20380 20594 20392
rect 21177 20383 21235 20389
rect 21177 20380 21189 20383
rect 20588 20352 21189 20380
rect 20588 20340 20594 20352
rect 21177 20349 21189 20352
rect 21223 20349 21235 20383
rect 21177 20343 21235 20349
rect 18874 20312 18880 20324
rect 18708 20284 18880 20312
rect 18874 20272 18880 20284
rect 18932 20272 18938 20324
rect 19337 20315 19395 20321
rect 19337 20281 19349 20315
rect 19383 20312 19395 20315
rect 19383 20284 20116 20312
rect 19383 20281 19395 20284
rect 19337 20275 19395 20281
rect 19426 20244 19432 20256
rect 15212 20216 19432 20244
rect 14553 20207 14611 20213
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 20088 20253 20116 20284
rect 20162 20272 20168 20324
rect 20220 20312 20226 20324
rect 20625 20315 20683 20321
rect 20625 20312 20637 20315
rect 20220 20284 20637 20312
rect 20220 20272 20226 20284
rect 20625 20281 20637 20284
rect 20671 20281 20683 20315
rect 20806 20312 20812 20324
rect 20767 20284 20812 20312
rect 20625 20275 20683 20281
rect 20806 20272 20812 20284
rect 20864 20272 20870 20324
rect 21358 20312 21364 20324
rect 21319 20284 21364 20312
rect 21358 20272 21364 20284
rect 21416 20272 21422 20324
rect 20073 20247 20131 20253
rect 20073 20213 20085 20247
rect 20119 20213 20131 20247
rect 20073 20207 20131 20213
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 1302 20000 1308 20052
rect 1360 20040 1366 20052
rect 1397 20043 1455 20049
rect 1397 20040 1409 20043
rect 1360 20012 1409 20040
rect 1360 20000 1366 20012
rect 1397 20009 1409 20012
rect 1443 20009 1455 20043
rect 2038 20040 2044 20052
rect 1999 20012 2044 20040
rect 1397 20003 1455 20009
rect 2038 20000 2044 20012
rect 2096 20000 2102 20052
rect 2498 20040 2504 20052
rect 2459 20012 2504 20040
rect 2498 20000 2504 20012
rect 2556 20000 2562 20052
rect 2866 20040 2872 20052
rect 2827 20012 2872 20040
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 3786 20040 3792 20052
rect 3747 20012 3792 20040
rect 3786 20000 3792 20012
rect 3844 20000 3850 20052
rect 4433 20043 4491 20049
rect 4433 20009 4445 20043
rect 4479 20040 4491 20043
rect 5442 20040 5448 20052
rect 4479 20012 5448 20040
rect 4479 20009 4491 20012
rect 4433 20003 4491 20009
rect 5442 20000 5448 20012
rect 5500 20000 5506 20052
rect 6822 20040 6828 20052
rect 6783 20012 6828 20040
rect 6822 20000 6828 20012
rect 6880 20000 6886 20052
rect 8294 20000 8300 20052
rect 8352 20040 8358 20052
rect 9677 20043 9735 20049
rect 9677 20040 9689 20043
rect 8352 20012 9689 20040
rect 8352 20000 8358 20012
rect 9677 20009 9689 20012
rect 9723 20009 9735 20043
rect 9677 20003 9735 20009
rect 10318 20000 10324 20052
rect 10376 20040 10382 20052
rect 11149 20043 11207 20049
rect 11149 20040 11161 20043
rect 10376 20012 11161 20040
rect 10376 20000 10382 20012
rect 11149 20009 11161 20012
rect 11195 20009 11207 20043
rect 11149 20003 11207 20009
rect 12069 20043 12127 20049
rect 12069 20009 12081 20043
rect 12115 20040 12127 20043
rect 16298 20040 16304 20052
rect 12115 20012 16304 20040
rect 12115 20009 12127 20012
rect 12069 20003 12127 20009
rect 16298 20000 16304 20012
rect 16356 20000 16362 20052
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 17773 20043 17831 20049
rect 17773 20040 17785 20043
rect 16632 20012 17785 20040
rect 16632 20000 16638 20012
rect 17773 20009 17785 20012
rect 17819 20009 17831 20043
rect 17773 20003 17831 20009
rect 19334 20000 19340 20052
rect 19392 20040 19398 20052
rect 19889 20043 19947 20049
rect 19889 20040 19901 20043
rect 19392 20012 19901 20040
rect 19392 20000 19398 20012
rect 19889 20009 19901 20012
rect 19935 20009 19947 20043
rect 19889 20003 19947 20009
rect 3513 19975 3571 19981
rect 3513 19941 3525 19975
rect 3559 19972 3571 19975
rect 4706 19972 4712 19984
rect 3559 19944 4712 19972
rect 3559 19941 3571 19944
rect 3513 19935 3571 19941
rect 4706 19932 4712 19944
rect 4764 19932 4770 19984
rect 5074 19932 5080 19984
rect 5132 19972 5138 19984
rect 5169 19975 5227 19981
rect 5169 19972 5181 19975
rect 5132 19944 5181 19972
rect 5132 19932 5138 19944
rect 5169 19941 5181 19944
rect 5215 19941 5227 19975
rect 5169 19935 5227 19941
rect 5350 19932 5356 19984
rect 5408 19972 5414 19984
rect 5537 19975 5595 19981
rect 5537 19972 5549 19975
rect 5408 19944 5549 19972
rect 5408 19932 5414 19944
rect 5537 19941 5549 19944
rect 5583 19941 5595 19975
rect 5537 19935 5595 19941
rect 5810 19932 5816 19984
rect 5868 19972 5874 19984
rect 5868 19944 6408 19972
rect 5868 19932 5874 19944
rect 1762 19864 1768 19916
rect 1820 19904 1826 19916
rect 4525 19907 4583 19913
rect 1820 19876 4384 19904
rect 1820 19864 1826 19876
rect 4246 19836 4252 19848
rect 4207 19808 4252 19836
rect 4246 19796 4252 19808
rect 4304 19796 4310 19848
rect 4356 19836 4384 19876
rect 4525 19873 4537 19907
rect 4571 19904 4583 19907
rect 4798 19904 4804 19916
rect 4571 19876 4804 19904
rect 4571 19873 4583 19876
rect 4525 19867 4583 19873
rect 4798 19864 4804 19876
rect 4856 19864 4862 19916
rect 5258 19864 5264 19916
rect 5316 19904 5322 19916
rect 5718 19904 5724 19916
rect 5316 19876 5724 19904
rect 5316 19864 5322 19876
rect 5718 19864 5724 19876
rect 5776 19904 5782 19916
rect 5905 19907 5963 19913
rect 5905 19904 5917 19907
rect 5776 19876 5917 19904
rect 5776 19864 5782 19876
rect 5905 19873 5917 19876
rect 5951 19873 5963 19907
rect 6380 19904 6408 19944
rect 6454 19932 6460 19984
rect 6512 19972 6518 19984
rect 7101 19975 7159 19981
rect 7101 19972 7113 19975
rect 6512 19944 7113 19972
rect 6512 19932 6518 19944
rect 7101 19941 7113 19944
rect 7147 19941 7159 19975
rect 7101 19935 7159 19941
rect 7668 19944 9076 19972
rect 6641 19907 6699 19913
rect 6641 19904 6653 19907
rect 6380 19876 6653 19904
rect 5905 19867 5963 19873
rect 6641 19873 6653 19876
rect 6687 19904 6699 19907
rect 6730 19904 6736 19916
rect 6687 19876 6736 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 7668 19904 7696 19944
rect 7834 19913 7840 19916
rect 7828 19904 7840 19913
rect 6886 19876 7696 19904
rect 7795 19876 7840 19904
rect 5166 19836 5172 19848
rect 4356 19808 5172 19836
rect 5166 19796 5172 19808
rect 5224 19796 5230 19848
rect 4614 19728 4620 19780
rect 4672 19768 4678 19780
rect 6089 19771 6147 19777
rect 4672 19740 5672 19768
rect 4672 19728 4678 19740
rect 4890 19700 4896 19712
rect 4851 19672 4896 19700
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 5644 19700 5672 19740
rect 6089 19737 6101 19771
rect 6135 19768 6147 19771
rect 6886 19768 6914 19876
rect 7828 19867 7840 19876
rect 7834 19864 7840 19867
rect 7892 19864 7898 19916
rect 7190 19796 7196 19848
rect 7248 19836 7254 19848
rect 7561 19839 7619 19845
rect 7561 19836 7573 19839
rect 7248 19808 7573 19836
rect 7248 19796 7254 19808
rect 7561 19805 7573 19808
rect 7607 19805 7619 19839
rect 7561 19799 7619 19805
rect 6135 19740 6914 19768
rect 6135 19737 6147 19740
rect 6089 19731 6147 19737
rect 8570 19700 8576 19712
rect 5644 19672 8576 19700
rect 8570 19660 8576 19672
rect 8628 19660 8634 19712
rect 8938 19700 8944 19712
rect 8899 19672 8944 19700
rect 8938 19660 8944 19672
rect 8996 19660 9002 19712
rect 9048 19700 9076 19944
rect 9766 19932 9772 19984
rect 9824 19972 9830 19984
rect 10781 19975 10839 19981
rect 10781 19972 10793 19975
rect 9824 19944 10793 19972
rect 9824 19932 9830 19944
rect 10781 19941 10793 19944
rect 10827 19941 10839 19975
rect 10781 19935 10839 19941
rect 10870 19932 10876 19984
rect 10928 19972 10934 19984
rect 14553 19975 14611 19981
rect 14553 19972 14565 19975
rect 10928 19944 14565 19972
rect 10928 19932 10934 19944
rect 14553 19941 14565 19944
rect 14599 19941 14611 19975
rect 14553 19935 14611 19941
rect 15194 19932 15200 19984
rect 15252 19972 15258 19984
rect 15289 19975 15347 19981
rect 15289 19972 15301 19975
rect 15252 19944 15301 19972
rect 15252 19932 15258 19944
rect 15289 19941 15301 19944
rect 15335 19941 15347 19975
rect 15289 19935 15347 19941
rect 15378 19932 15384 19984
rect 15436 19972 15442 19984
rect 15841 19975 15899 19981
rect 15841 19972 15853 19975
rect 15436 19944 15853 19972
rect 15436 19932 15442 19944
rect 15841 19941 15853 19944
rect 15887 19941 15899 19975
rect 15841 19935 15899 19941
rect 15930 19932 15936 19984
rect 15988 19972 15994 19984
rect 17129 19975 17187 19981
rect 17129 19972 17141 19975
rect 15988 19944 17141 19972
rect 15988 19932 15994 19944
rect 17129 19941 17141 19944
rect 17175 19941 17187 19975
rect 19702 19972 19708 19984
rect 17129 19935 17187 19941
rect 19536 19944 19708 19972
rect 9214 19864 9220 19916
rect 9272 19904 9278 19916
rect 10413 19907 10471 19913
rect 10413 19904 10425 19907
rect 9272 19876 10425 19904
rect 9272 19864 9278 19876
rect 10413 19873 10425 19876
rect 10459 19873 10471 19907
rect 10413 19867 10471 19873
rect 11698 19864 11704 19916
rect 11756 19904 11762 19916
rect 11885 19907 11943 19913
rect 11885 19904 11897 19907
rect 11756 19876 11897 19904
rect 11756 19864 11762 19876
rect 11885 19873 11897 19876
rect 11931 19904 11943 19907
rect 12713 19907 12771 19913
rect 12713 19904 12725 19907
rect 11931 19876 12725 19904
rect 11931 19873 11943 19876
rect 11885 19867 11943 19873
rect 12713 19873 12725 19876
rect 12759 19873 12771 19907
rect 14642 19904 14648 19916
rect 14603 19876 14648 19904
rect 12713 19867 12771 19873
rect 14642 19864 14648 19876
rect 14700 19864 14706 19916
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19904 15531 19907
rect 15562 19904 15568 19916
rect 15519 19876 15568 19904
rect 15519 19873 15531 19876
rect 15473 19867 15531 19873
rect 15562 19864 15568 19876
rect 15620 19864 15626 19916
rect 16022 19904 16028 19916
rect 15983 19876 16028 19904
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 17313 19907 17371 19913
rect 17313 19873 17325 19907
rect 17359 19904 17371 19907
rect 17402 19904 17408 19916
rect 17359 19876 17408 19904
rect 17359 19873 17371 19876
rect 17313 19867 17371 19873
rect 17402 19864 17408 19876
rect 17460 19864 17466 19916
rect 17770 19864 17776 19916
rect 17828 19904 17834 19916
rect 19536 19913 19564 19944
rect 19702 19932 19708 19944
rect 19760 19932 19766 19984
rect 20346 19932 20352 19984
rect 20404 19972 20410 19984
rect 20533 19975 20591 19981
rect 20533 19972 20545 19975
rect 20404 19944 20545 19972
rect 20404 19932 20410 19944
rect 20533 19941 20545 19944
rect 20579 19941 20591 19975
rect 20533 19935 20591 19941
rect 17865 19907 17923 19913
rect 17865 19904 17877 19907
rect 17828 19876 17877 19904
rect 17828 19864 17834 19876
rect 17865 19873 17877 19876
rect 17911 19873 17923 19907
rect 17865 19867 17923 19873
rect 19521 19907 19579 19913
rect 19521 19873 19533 19907
rect 19567 19873 19579 19907
rect 19521 19867 19579 19873
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19668 19876 19993 19904
rect 19668 19864 19674 19876
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 19981 19867 20039 19873
rect 20622 19864 20628 19916
rect 20680 19904 20686 19916
rect 21177 19907 21235 19913
rect 21177 19904 21189 19907
rect 20680 19876 21189 19904
rect 20680 19864 20686 19876
rect 21177 19873 21189 19876
rect 21223 19873 21235 19907
rect 21177 19867 21235 19873
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19836 9459 19839
rect 9674 19836 9680 19848
rect 9447 19808 9680 19836
rect 9447 19805 9459 19808
rect 9401 19799 9459 19805
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 10962 19796 10968 19848
rect 11020 19836 11026 19848
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 11020 19808 12449 19836
rect 11020 19796 11026 19808
rect 12437 19805 12449 19808
rect 12483 19805 12495 19839
rect 12437 19799 12495 19805
rect 14461 19839 14519 19845
rect 14461 19805 14473 19839
rect 14507 19836 14519 19839
rect 14826 19836 14832 19848
rect 14507 19808 14832 19836
rect 14507 19805 14519 19808
rect 14461 19799 14519 19805
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 16574 19836 16580 19848
rect 16535 19808 16580 19836
rect 16574 19796 16580 19808
rect 16632 19796 16638 19848
rect 18690 19836 18696 19848
rect 18651 19808 18696 19836
rect 18690 19796 18696 19808
rect 18748 19796 18754 19848
rect 19886 19796 19892 19848
rect 19944 19836 19950 19848
rect 20349 19839 20407 19845
rect 20349 19836 20361 19839
rect 19944 19808 20361 19836
rect 19944 19796 19950 19808
rect 20349 19805 20361 19808
rect 20395 19805 20407 19839
rect 20349 19799 20407 19805
rect 9122 19728 9128 19780
rect 9180 19768 9186 19780
rect 10045 19771 10103 19777
rect 10045 19768 10057 19771
rect 9180 19740 10057 19768
rect 9180 19728 9186 19740
rect 10045 19737 10057 19740
rect 10091 19737 10103 19771
rect 10045 19731 10103 19737
rect 11238 19728 11244 19780
rect 11296 19768 11302 19780
rect 15013 19771 15071 19777
rect 11296 19740 14964 19768
rect 11296 19728 11302 19740
rect 11146 19700 11152 19712
rect 9048 19672 11152 19700
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 12894 19660 12900 19712
rect 12952 19700 12958 19712
rect 13081 19703 13139 19709
rect 13081 19700 13093 19703
rect 12952 19672 13093 19700
rect 12952 19660 12958 19672
rect 13081 19669 13093 19672
rect 13127 19669 13139 19703
rect 14936 19700 14964 19740
rect 15013 19737 15025 19771
rect 15059 19768 15071 19771
rect 16666 19768 16672 19780
rect 15059 19740 16672 19768
rect 15059 19737 15071 19740
rect 15013 19731 15071 19737
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 21358 19768 21364 19780
rect 21319 19740 21364 19768
rect 21358 19728 21364 19740
rect 21416 19728 21422 19780
rect 16758 19700 16764 19712
rect 14936 19672 16764 19700
rect 13081 19663 13139 19669
rect 16758 19660 16764 19672
rect 16816 19660 16822 19712
rect 17586 19660 17592 19712
rect 17644 19700 17650 19712
rect 20990 19700 20996 19712
rect 17644 19672 20996 19700
rect 17644 19660 17650 19672
rect 20990 19660 20996 19672
rect 21048 19660 21054 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 7098 19456 7104 19508
rect 7156 19496 7162 19508
rect 7561 19499 7619 19505
rect 7561 19496 7573 19499
rect 7156 19468 7573 19496
rect 7156 19456 7162 19468
rect 7561 19465 7573 19468
rect 7607 19465 7619 19499
rect 7561 19459 7619 19465
rect 7742 19456 7748 19508
rect 7800 19496 7806 19508
rect 12342 19496 12348 19508
rect 7800 19468 12348 19496
rect 7800 19456 7806 19468
rect 12342 19456 12348 19468
rect 12400 19456 12406 19508
rect 14274 19496 14280 19508
rect 12452 19468 14280 19496
rect 7285 19431 7343 19437
rect 7285 19397 7297 19431
rect 7331 19428 7343 19431
rect 7834 19428 7840 19440
rect 7331 19400 7840 19428
rect 7331 19397 7343 19400
rect 7285 19391 7343 19397
rect 7834 19388 7840 19400
rect 7892 19428 7898 19440
rect 12452 19428 12480 19468
rect 14274 19456 14280 19468
rect 14332 19456 14338 19508
rect 18598 19496 18604 19508
rect 18559 19468 18604 19496
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 19245 19499 19303 19505
rect 19245 19465 19257 19499
rect 19291 19496 19303 19499
rect 20530 19496 20536 19508
rect 19291 19468 20536 19496
rect 19291 19465 19303 19468
rect 19245 19459 19303 19465
rect 20530 19456 20536 19468
rect 20588 19456 20594 19508
rect 7892 19400 8156 19428
rect 7892 19388 7898 19400
rect 6914 19320 6920 19372
rect 6972 19360 6978 19372
rect 8128 19369 8156 19400
rect 8220 19400 10732 19428
rect 8113 19363 8171 19369
rect 6972 19332 8064 19360
rect 6972 19320 6978 19332
rect 3878 19252 3884 19304
rect 3936 19292 3942 19304
rect 4065 19295 4123 19301
rect 4065 19292 4077 19295
rect 3936 19264 4077 19292
rect 3936 19252 3942 19264
rect 4065 19261 4077 19264
rect 4111 19261 4123 19295
rect 4798 19292 4804 19304
rect 4065 19255 4123 19261
rect 4172 19264 4804 19292
rect 3513 19227 3571 19233
rect 3513 19193 3525 19227
rect 3559 19224 3571 19227
rect 4172 19224 4200 19264
rect 4798 19252 4804 19264
rect 4856 19292 4862 19304
rect 5902 19292 5908 19304
rect 4856 19264 5580 19292
rect 5863 19264 5908 19292
rect 4856 19252 4862 19264
rect 3559 19196 4200 19224
rect 3559 19193 3571 19196
rect 3513 19187 3571 19193
rect 4246 19184 4252 19236
rect 4304 19233 4310 19236
rect 4304 19227 4368 19233
rect 4304 19193 4322 19227
rect 4356 19193 4368 19227
rect 4304 19187 4368 19193
rect 4304 19184 4310 19187
rect 4798 19116 4804 19168
rect 4856 19156 4862 19168
rect 5445 19159 5503 19165
rect 5445 19156 5457 19159
rect 4856 19128 5457 19156
rect 4856 19116 4862 19128
rect 5445 19125 5457 19128
rect 5491 19125 5503 19159
rect 5552 19156 5580 19264
rect 5902 19252 5908 19264
rect 5960 19292 5966 19304
rect 7190 19292 7196 19304
rect 5960 19264 7196 19292
rect 5960 19252 5966 19264
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 8036 19292 8064 19332
rect 8113 19329 8125 19363
rect 8159 19329 8171 19363
rect 8113 19323 8171 19329
rect 8220 19292 8248 19400
rect 8297 19363 8355 19369
rect 8297 19329 8309 19363
rect 8343 19360 8355 19363
rect 8662 19360 8668 19372
rect 8343 19332 8668 19360
rect 8343 19329 8355 19332
rect 8297 19323 8355 19329
rect 8662 19320 8668 19332
rect 8720 19320 8726 19372
rect 8938 19320 8944 19372
rect 8996 19360 9002 19372
rect 9398 19360 9404 19372
rect 8996 19332 9404 19360
rect 8996 19320 9002 19332
rect 9398 19320 9404 19332
rect 9456 19320 9462 19372
rect 9674 19292 9680 19304
rect 8036 19264 8248 19292
rect 9635 19264 9680 19292
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 6172 19227 6230 19233
rect 6172 19193 6184 19227
rect 6218 19224 6230 19227
rect 6638 19224 6644 19236
rect 6218 19196 6644 19224
rect 6218 19193 6230 19196
rect 6172 19187 6230 19193
rect 6638 19184 6644 19196
rect 6696 19184 6702 19236
rect 8389 19227 8447 19233
rect 8389 19224 8401 19227
rect 6886 19196 8401 19224
rect 6886 19156 6914 19196
rect 8389 19193 8401 19196
rect 8435 19224 8447 19227
rect 8938 19224 8944 19236
rect 8435 19196 8944 19224
rect 8435 19193 8447 19196
rect 8389 19187 8447 19193
rect 8938 19184 8944 19196
rect 8996 19184 9002 19236
rect 10704 19224 10732 19400
rect 11808 19400 12480 19428
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19292 10839 19295
rect 10870 19292 10876 19304
rect 10827 19264 10876 19292
rect 10827 19261 10839 19264
rect 10781 19255 10839 19261
rect 10870 19252 10876 19264
rect 10928 19252 10934 19304
rect 11808 19292 11836 19400
rect 15838 19388 15844 19440
rect 15896 19428 15902 19440
rect 18325 19431 18383 19437
rect 15896 19400 18276 19428
rect 15896 19388 15902 19400
rect 16301 19363 16359 19369
rect 16301 19329 16313 19363
rect 16347 19329 16359 19363
rect 16301 19323 16359 19329
rect 16485 19363 16543 19369
rect 16485 19329 16497 19363
rect 16531 19360 16543 19363
rect 16666 19360 16672 19372
rect 16531 19332 16672 19360
rect 16531 19329 16543 19332
rect 16485 19323 16543 19329
rect 10980 19264 11836 19292
rect 12437 19295 12495 19301
rect 10980 19224 11008 19264
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 13170 19292 13176 19304
rect 12483 19264 13176 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 13170 19252 13176 19264
rect 13228 19292 13234 19304
rect 14550 19292 14556 19304
rect 13228 19264 14556 19292
rect 13228 19252 13234 19264
rect 14550 19252 14556 19264
rect 14608 19252 14614 19304
rect 14826 19301 14832 19304
rect 14820 19292 14832 19301
rect 14787 19264 14832 19292
rect 14820 19255 14832 19264
rect 14826 19252 14832 19255
rect 14884 19252 14890 19304
rect 16316 19292 16344 19323
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 18248 19360 18276 19400
rect 18325 19397 18337 19431
rect 18371 19428 18383 19431
rect 20162 19428 20168 19440
rect 18371 19400 20168 19428
rect 18371 19397 18383 19400
rect 18325 19391 18383 19397
rect 20162 19388 20168 19400
rect 20220 19388 20226 19440
rect 19886 19360 19892 19372
rect 18248 19332 19892 19360
rect 19886 19320 19892 19332
rect 19944 19320 19950 19372
rect 16574 19292 16580 19304
rect 15948 19264 16344 19292
rect 16535 19264 16580 19292
rect 10704 19196 11008 19224
rect 11048 19227 11106 19233
rect 11048 19193 11060 19227
rect 11094 19224 11106 19227
rect 11330 19224 11336 19236
rect 11094 19196 11336 19224
rect 11094 19193 11106 19196
rect 11048 19187 11106 19193
rect 11330 19184 11336 19196
rect 11388 19184 11394 19236
rect 12682 19227 12740 19233
rect 12682 19224 12694 19227
rect 12176 19196 12694 19224
rect 5552 19128 6914 19156
rect 8757 19159 8815 19165
rect 5445 19119 5503 19125
rect 8757 19125 8769 19159
rect 8803 19156 8815 19159
rect 9585 19159 9643 19165
rect 9585 19156 9597 19159
rect 8803 19128 9597 19156
rect 8803 19125 8815 19128
rect 8757 19119 8815 19125
rect 9585 19125 9597 19128
rect 9631 19125 9643 19159
rect 9585 19119 9643 19125
rect 10045 19159 10103 19165
rect 10045 19125 10057 19159
rect 10091 19156 10103 19159
rect 11974 19156 11980 19168
rect 10091 19128 11980 19156
rect 10091 19125 10103 19128
rect 10045 19119 10103 19125
rect 11974 19116 11980 19128
rect 12032 19116 12038 19168
rect 12066 19116 12072 19168
rect 12124 19156 12130 19168
rect 12176 19165 12204 19196
rect 12682 19193 12694 19196
rect 12728 19193 12740 19227
rect 12682 19187 12740 19193
rect 12161 19159 12219 19165
rect 12161 19156 12173 19159
rect 12124 19128 12173 19156
rect 12124 19116 12130 19128
rect 12161 19125 12173 19128
rect 12207 19125 12219 19159
rect 13814 19156 13820 19168
rect 13775 19128 13820 19156
rect 12161 19119 12219 19125
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 15948 19165 15976 19264
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 17034 19252 17040 19304
rect 17092 19292 17098 19304
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 17092 19264 17233 19292
rect 17092 19252 17098 19264
rect 17221 19261 17233 19264
rect 17267 19261 17279 19295
rect 17221 19255 17279 19261
rect 17494 19252 17500 19304
rect 17552 19292 17558 19304
rect 18141 19295 18199 19301
rect 18141 19292 18153 19295
rect 17552 19264 18153 19292
rect 17552 19252 17558 19264
rect 18141 19261 18153 19264
rect 18187 19261 18199 19295
rect 18141 19255 18199 19261
rect 18785 19295 18843 19301
rect 18785 19261 18797 19295
rect 18831 19261 18843 19295
rect 19058 19292 19064 19304
rect 19019 19264 19064 19292
rect 18785 19255 18843 19261
rect 17310 19184 17316 19236
rect 17368 19224 17374 19236
rect 17405 19227 17463 19233
rect 17405 19224 17417 19227
rect 17368 19196 17417 19224
rect 17368 19184 17374 19196
rect 17405 19193 17417 19196
rect 17451 19193 17463 19227
rect 18800 19224 18828 19255
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 19981 19295 20039 19301
rect 19981 19261 19993 19295
rect 20027 19292 20039 19295
rect 20070 19292 20076 19304
rect 20027 19264 20076 19292
rect 20027 19261 20039 19264
rect 19981 19255 20039 19261
rect 20070 19252 20076 19264
rect 20128 19252 20134 19304
rect 20438 19292 20444 19304
rect 20399 19264 20444 19292
rect 20438 19252 20444 19264
rect 20496 19252 20502 19304
rect 17405 19187 17463 19193
rect 17512 19196 18828 19224
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 15896 19128 15945 19156
rect 15896 19116 15902 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 16942 19156 16948 19168
rect 16903 19128 16948 19156
rect 15933 19119 15991 19125
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 17034 19116 17040 19168
rect 17092 19156 17098 19168
rect 17512 19156 17540 19196
rect 20530 19184 20536 19236
rect 20588 19224 20594 19236
rect 20625 19227 20683 19233
rect 20625 19224 20637 19227
rect 20588 19196 20637 19224
rect 20588 19184 20594 19196
rect 20625 19193 20637 19196
rect 20671 19193 20683 19227
rect 20625 19187 20683 19193
rect 20898 19184 20904 19236
rect 20956 19224 20962 19236
rect 21177 19227 21235 19233
rect 21177 19224 21189 19227
rect 20956 19196 21189 19224
rect 20956 19184 20962 19196
rect 21177 19193 21189 19196
rect 21223 19193 21235 19227
rect 21358 19224 21364 19236
rect 21319 19196 21364 19224
rect 21177 19187 21235 19193
rect 21358 19184 21364 19196
rect 21416 19184 21422 19236
rect 17092 19128 17540 19156
rect 20073 19159 20131 19165
rect 17092 19116 17098 19128
rect 20073 19125 20085 19159
rect 20119 19156 20131 19159
rect 21542 19156 21548 19168
rect 20119 19128 21548 19156
rect 20119 19125 20131 19128
rect 20073 19119 20131 19125
rect 21542 19116 21548 19128
rect 21600 19116 21606 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 3697 18955 3755 18961
rect 3697 18921 3709 18955
rect 3743 18952 3755 18955
rect 4246 18952 4252 18964
rect 3743 18924 4252 18952
rect 3743 18921 3755 18924
rect 3697 18915 3755 18921
rect 4246 18912 4252 18924
rect 4304 18912 4310 18964
rect 4709 18955 4767 18961
rect 4709 18921 4721 18955
rect 4755 18952 4767 18955
rect 4890 18952 4896 18964
rect 4755 18924 4896 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 4890 18912 4896 18924
rect 4948 18912 4954 18964
rect 5534 18912 5540 18964
rect 5592 18952 5598 18964
rect 5721 18955 5779 18961
rect 5721 18952 5733 18955
rect 5592 18924 5733 18952
rect 5592 18912 5598 18924
rect 5721 18921 5733 18924
rect 5767 18921 5779 18955
rect 5721 18915 5779 18921
rect 7558 18912 7564 18964
rect 7616 18952 7622 18964
rect 7653 18955 7711 18961
rect 7653 18952 7665 18955
rect 7616 18924 7665 18952
rect 7616 18912 7622 18924
rect 7653 18921 7665 18924
rect 7699 18921 7711 18955
rect 11330 18952 11336 18964
rect 11291 18924 11336 18952
rect 7653 18915 7711 18921
rect 11330 18912 11336 18924
rect 11388 18912 11394 18964
rect 11974 18912 11980 18964
rect 12032 18952 12038 18964
rect 14734 18952 14740 18964
rect 12032 18924 14596 18952
rect 14695 18924 14740 18952
rect 12032 18912 12038 18924
rect 6730 18844 6736 18896
rect 6788 18884 6794 18896
rect 8021 18887 8079 18893
rect 8021 18884 8033 18887
rect 6788 18856 8033 18884
rect 6788 18844 6794 18856
rect 8021 18853 8033 18856
rect 8067 18853 8079 18887
rect 13624 18887 13682 18893
rect 8021 18847 8079 18853
rect 10060 18856 10916 18884
rect 1762 18776 1768 18828
rect 1820 18816 1826 18828
rect 2573 18819 2631 18825
rect 2573 18816 2585 18819
rect 1820 18788 2585 18816
rect 1820 18776 1826 18788
rect 2573 18785 2585 18788
rect 2619 18785 2631 18819
rect 2573 18779 2631 18785
rect 4617 18819 4675 18825
rect 4617 18785 4629 18819
rect 4663 18816 4675 18819
rect 5261 18819 5319 18825
rect 5261 18816 5273 18819
rect 4663 18788 5273 18816
rect 4663 18785 4675 18788
rect 4617 18779 4675 18785
rect 5261 18785 5273 18788
rect 5307 18785 5319 18819
rect 7190 18816 7196 18828
rect 7151 18788 7196 18816
rect 5261 18779 5319 18785
rect 7190 18776 7196 18788
rect 7248 18776 7254 18828
rect 10060 18816 10088 18856
rect 10226 18825 10232 18828
rect 10220 18816 10232 18825
rect 7392 18788 10088 18816
rect 10187 18788 10232 18816
rect 2317 18751 2375 18757
rect 2317 18717 2329 18751
rect 2363 18717 2375 18751
rect 4798 18748 4804 18760
rect 4759 18720 4804 18748
rect 2317 18711 2375 18717
rect 2332 18612 2360 18711
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 6917 18751 6975 18757
rect 6917 18717 6929 18751
rect 6963 18748 6975 18751
rect 7282 18748 7288 18760
rect 6963 18720 7288 18748
rect 6963 18717 6975 18720
rect 6917 18711 6975 18717
rect 7282 18708 7288 18720
rect 7340 18708 7346 18760
rect 7392 18689 7420 18788
rect 10220 18779 10232 18788
rect 10226 18776 10232 18779
rect 10284 18776 10290 18828
rect 10888 18816 10916 18856
rect 11716 18856 13584 18884
rect 11716 18816 11744 18856
rect 10888 18788 11744 18816
rect 11790 18776 11796 18828
rect 11848 18816 11854 18828
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11848 18788 12173 18816
rect 11848 18776 11854 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 12253 18819 12311 18825
rect 12253 18785 12265 18819
rect 12299 18816 12311 18819
rect 12434 18816 12440 18828
rect 12299 18788 12440 18816
rect 12299 18785 12311 18788
rect 12253 18779 12311 18785
rect 12434 18776 12440 18788
rect 12492 18776 12498 18828
rect 13170 18776 13176 18828
rect 13228 18816 13234 18828
rect 13357 18819 13415 18825
rect 13357 18816 13369 18819
rect 13228 18788 13369 18816
rect 13228 18776 13234 18788
rect 13357 18785 13369 18788
rect 13403 18785 13415 18819
rect 13556 18816 13584 18856
rect 13624 18853 13636 18887
rect 13670 18884 13682 18887
rect 13814 18884 13820 18896
rect 13670 18856 13820 18884
rect 13670 18853 13682 18856
rect 13624 18847 13682 18853
rect 13814 18844 13820 18856
rect 13872 18844 13878 18896
rect 14568 18884 14596 18924
rect 14734 18912 14740 18924
rect 14792 18912 14798 18964
rect 16577 18955 16635 18961
rect 16577 18921 16589 18955
rect 16623 18952 16635 18955
rect 17034 18952 17040 18964
rect 16623 18924 17040 18952
rect 16623 18921 16635 18924
rect 16577 18915 16635 18921
rect 17034 18912 17040 18924
rect 17092 18912 17098 18964
rect 17494 18952 17500 18964
rect 17455 18924 17500 18952
rect 17494 18912 17500 18924
rect 17552 18912 17558 18964
rect 18138 18912 18144 18964
rect 18196 18952 18202 18964
rect 19061 18955 19119 18961
rect 19061 18952 19073 18955
rect 18196 18924 19073 18952
rect 18196 18912 18202 18924
rect 19061 18921 19073 18924
rect 19107 18921 19119 18955
rect 19518 18952 19524 18964
rect 19479 18924 19524 18952
rect 19061 18915 19119 18921
rect 19518 18912 19524 18924
rect 19576 18912 19582 18964
rect 20165 18955 20223 18961
rect 20165 18921 20177 18955
rect 20211 18952 20223 18955
rect 22646 18952 22652 18964
rect 20211 18924 22652 18952
rect 20211 18921 20223 18924
rect 20165 18915 20223 18921
rect 22646 18912 22652 18924
rect 22704 18912 22710 18964
rect 20809 18887 20867 18893
rect 14568 18856 17356 18884
rect 16393 18819 16451 18825
rect 13556 18788 14412 18816
rect 13357 18779 13415 18785
rect 9953 18751 10011 18757
rect 9953 18717 9965 18751
rect 9999 18717 10011 18751
rect 12066 18748 12072 18760
rect 12027 18720 12072 18748
rect 9953 18711 10011 18717
rect 7377 18683 7435 18689
rect 7377 18649 7389 18683
rect 7423 18649 7435 18683
rect 7377 18643 7435 18649
rect 3878 18612 3884 18624
rect 2332 18584 3884 18612
rect 3878 18572 3884 18584
rect 3936 18572 3942 18624
rect 4246 18612 4252 18624
rect 4207 18584 4252 18612
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 8938 18612 8944 18624
rect 8899 18584 8944 18612
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 9968 18612 9996 18711
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 13078 18748 13084 18760
rect 13039 18720 13084 18748
rect 13078 18708 13084 18720
rect 13136 18708 13142 18760
rect 14384 18748 14412 18788
rect 16393 18785 16405 18819
rect 16439 18816 16451 18819
rect 16942 18816 16948 18828
rect 16439 18788 16948 18816
rect 16439 18785 16451 18788
rect 16393 18779 16451 18785
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 17328 18825 17356 18856
rect 20809 18853 20821 18887
rect 20855 18884 20867 18887
rect 22094 18884 22100 18896
rect 20855 18856 22100 18884
rect 20855 18853 20867 18856
rect 20809 18847 20867 18853
rect 22094 18844 22100 18856
rect 22152 18844 22158 18896
rect 17313 18819 17371 18825
rect 17313 18785 17325 18819
rect 17359 18785 17371 18819
rect 18046 18816 18052 18828
rect 18007 18788 18052 18816
rect 17313 18779 17371 18785
rect 18046 18776 18052 18788
rect 18104 18776 18110 18828
rect 19058 18816 19064 18828
rect 18156 18788 19064 18816
rect 18156 18748 18184 18788
rect 19058 18776 19064 18788
rect 19116 18776 19122 18828
rect 19242 18816 19248 18828
rect 19203 18788 19248 18816
rect 19242 18776 19248 18788
rect 19300 18776 19306 18828
rect 19702 18816 19708 18828
rect 19663 18788 19708 18816
rect 19702 18776 19708 18788
rect 19760 18776 19766 18828
rect 19978 18776 19984 18828
rect 20036 18816 20042 18828
rect 20073 18819 20131 18825
rect 20073 18816 20085 18819
rect 20036 18788 20085 18816
rect 20036 18776 20042 18788
rect 20073 18785 20085 18788
rect 20119 18785 20131 18819
rect 20073 18779 20131 18785
rect 20438 18776 20444 18828
rect 20496 18816 20502 18828
rect 20625 18819 20683 18825
rect 20625 18816 20637 18819
rect 20496 18788 20637 18816
rect 20496 18776 20502 18788
rect 20625 18785 20637 18788
rect 20671 18785 20683 18819
rect 21174 18816 21180 18828
rect 21135 18788 21180 18816
rect 20625 18779 20683 18785
rect 21174 18776 21180 18788
rect 21232 18776 21238 18828
rect 14384 18720 18184 18748
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18748 18567 18751
rect 18598 18748 18604 18760
rect 18555 18720 18604 18748
rect 18555 18717 18567 18720
rect 18509 18711 18567 18717
rect 18598 18708 18604 18720
rect 18656 18708 18662 18760
rect 18233 18683 18291 18689
rect 18233 18649 18245 18683
rect 18279 18680 18291 18683
rect 20254 18680 20260 18692
rect 18279 18652 20260 18680
rect 18279 18649 18291 18652
rect 18233 18643 18291 18649
rect 20254 18640 20260 18652
rect 20312 18640 20318 18692
rect 21358 18680 21364 18692
rect 21319 18652 21364 18680
rect 21358 18640 21364 18652
rect 21416 18640 21422 18692
rect 10962 18612 10968 18624
rect 9968 18584 10968 18612
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 12621 18615 12679 18621
rect 12621 18581 12633 18615
rect 12667 18612 12679 18615
rect 13354 18612 13360 18624
rect 12667 18584 13360 18612
rect 12667 18581 12679 18584
rect 12621 18575 12679 18581
rect 13354 18572 13360 18584
rect 13412 18572 13418 18624
rect 14642 18572 14648 18624
rect 14700 18612 14706 18624
rect 15197 18615 15255 18621
rect 15197 18612 15209 18615
rect 14700 18584 15209 18612
rect 14700 18572 14706 18584
rect 15197 18581 15209 18584
rect 15243 18581 15255 18615
rect 15197 18575 15255 18581
rect 17310 18572 17316 18624
rect 17368 18612 17374 18624
rect 21082 18612 21088 18624
rect 17368 18584 21088 18612
rect 17368 18572 17374 18584
rect 21082 18572 21088 18584
rect 21140 18572 21146 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 6638 18408 6644 18420
rect 6599 18380 6644 18408
rect 6638 18368 6644 18380
rect 6696 18368 6702 18420
rect 6917 18411 6975 18417
rect 6917 18377 6929 18411
rect 6963 18408 6975 18411
rect 7190 18408 7196 18420
rect 6963 18380 7196 18408
rect 6963 18377 6975 18380
rect 6917 18371 6975 18377
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 8938 18368 8944 18420
rect 8996 18408 9002 18420
rect 11701 18411 11759 18417
rect 8996 18380 10272 18408
rect 8996 18368 9002 18380
rect 6656 18272 6684 18368
rect 10244 18340 10272 18380
rect 11701 18377 11713 18411
rect 11747 18408 11759 18411
rect 18046 18408 18052 18420
rect 11747 18380 18052 18408
rect 11747 18377 11759 18380
rect 11701 18371 11759 18377
rect 18046 18368 18052 18380
rect 18104 18368 18110 18420
rect 19705 18411 19763 18417
rect 19705 18377 19717 18411
rect 19751 18408 19763 18411
rect 19794 18408 19800 18420
rect 19751 18380 19800 18408
rect 19751 18377 19763 18380
rect 19705 18371 19763 18377
rect 19794 18368 19800 18380
rect 19852 18368 19858 18420
rect 20349 18411 20407 18417
rect 20349 18377 20361 18411
rect 20395 18408 20407 18411
rect 20622 18408 20628 18420
rect 20395 18380 20628 18408
rect 20395 18377 20407 18380
rect 20349 18371 20407 18377
rect 20622 18368 20628 18380
rect 20680 18368 20686 18420
rect 20809 18411 20867 18417
rect 20809 18377 20821 18411
rect 20855 18408 20867 18411
rect 21174 18408 21180 18420
rect 20855 18380 21180 18408
rect 20855 18377 20867 18380
rect 20809 18371 20867 18377
rect 21174 18368 21180 18380
rect 21232 18368 21238 18420
rect 12710 18340 12716 18352
rect 10244 18312 12716 18340
rect 12710 18300 12716 18312
rect 12768 18300 12774 18352
rect 13814 18340 13820 18352
rect 13188 18312 13820 18340
rect 7469 18275 7527 18281
rect 7469 18272 7481 18275
rect 6656 18244 7481 18272
rect 7469 18241 7481 18244
rect 7515 18241 7527 18275
rect 7469 18235 7527 18241
rect 11149 18275 11207 18281
rect 11149 18241 11161 18275
rect 11195 18272 11207 18275
rect 11238 18272 11244 18284
rect 11195 18244 11244 18272
rect 11195 18241 11207 18244
rect 11149 18235 11207 18241
rect 11238 18232 11244 18244
rect 11296 18232 11302 18284
rect 13188 18281 13216 18312
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 16945 18343 17003 18349
rect 16945 18309 16957 18343
rect 16991 18340 17003 18343
rect 16991 18312 17356 18340
rect 16991 18309 17003 18312
rect 16945 18303 17003 18309
rect 17328 18284 17356 18312
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18241 13231 18275
rect 13354 18272 13360 18284
rect 13315 18244 13360 18272
rect 13173 18235 13231 18241
rect 13354 18232 13360 18244
rect 13412 18232 13418 18284
rect 14550 18232 14556 18284
rect 14608 18272 14614 18284
rect 15565 18275 15623 18281
rect 15565 18272 15577 18275
rect 14608 18244 15577 18272
rect 14608 18232 14614 18244
rect 15565 18241 15577 18244
rect 15611 18241 15623 18275
rect 17310 18272 17316 18284
rect 17223 18244 17316 18272
rect 15565 18235 15623 18241
rect 17310 18232 17316 18244
rect 17368 18232 17374 18284
rect 18322 18272 18328 18284
rect 18283 18244 18328 18272
rect 18322 18232 18328 18244
rect 18380 18232 18386 18284
rect 19334 18232 19340 18284
rect 19392 18272 19398 18284
rect 19392 18244 20668 18272
rect 19392 18232 19398 18244
rect 5258 18204 5264 18216
rect 5219 18176 5264 18204
rect 5258 18164 5264 18176
rect 5316 18204 5322 18216
rect 5902 18204 5908 18216
rect 5316 18176 5908 18204
rect 5316 18164 5322 18176
rect 5902 18164 5908 18176
rect 5960 18164 5966 18216
rect 7282 18204 7288 18216
rect 7243 18176 7288 18204
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 9309 18207 9367 18213
rect 9309 18173 9321 18207
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 5534 18145 5540 18148
rect 5528 18136 5540 18145
rect 5495 18108 5540 18136
rect 5528 18099 5540 18108
rect 5534 18096 5540 18099
rect 5592 18096 5598 18148
rect 9324 18136 9352 18167
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 9565 18207 9623 18213
rect 9565 18204 9577 18207
rect 9456 18176 9577 18204
rect 9456 18164 9462 18176
rect 9565 18173 9577 18176
rect 9611 18173 9623 18207
rect 9565 18167 9623 18173
rect 13078 18164 13084 18216
rect 13136 18204 13142 18216
rect 15838 18213 15844 18216
rect 13449 18207 13507 18213
rect 13449 18204 13461 18207
rect 13136 18176 13461 18204
rect 13136 18164 13142 18176
rect 13449 18173 13461 18176
rect 13495 18173 13507 18207
rect 13449 18167 13507 18173
rect 15832 18167 15844 18213
rect 15896 18204 15902 18216
rect 18598 18204 18604 18216
rect 15896 18176 15932 18204
rect 18559 18176 18604 18204
rect 15838 18164 15844 18167
rect 15896 18164 15902 18176
rect 18598 18164 18604 18176
rect 18656 18164 18662 18216
rect 20162 18204 20168 18216
rect 20123 18176 20168 18204
rect 20162 18164 20168 18176
rect 20220 18164 20226 18216
rect 20640 18213 20668 18244
rect 20625 18207 20683 18213
rect 20625 18173 20637 18207
rect 20671 18173 20683 18207
rect 20625 18167 20683 18173
rect 10962 18136 10968 18148
rect 9324 18108 10968 18136
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 11333 18139 11391 18145
rect 11333 18105 11345 18139
rect 11379 18136 11391 18139
rect 11977 18139 12035 18145
rect 11977 18136 11989 18139
rect 11379 18108 11989 18136
rect 11379 18105 11391 18108
rect 11333 18099 11391 18105
rect 11977 18105 11989 18108
rect 12023 18105 12035 18139
rect 11977 18099 12035 18105
rect 14182 18096 14188 18148
rect 14240 18136 14246 18148
rect 17497 18139 17555 18145
rect 17497 18136 17509 18139
rect 14240 18108 17509 18136
rect 14240 18096 14246 18108
rect 17497 18105 17509 18108
rect 17543 18105 17555 18139
rect 17497 18099 17555 18105
rect 20254 18096 20260 18148
rect 20312 18136 20318 18148
rect 21177 18139 21235 18145
rect 21177 18136 21189 18139
rect 20312 18108 21189 18136
rect 20312 18096 20318 18108
rect 21177 18105 21189 18108
rect 21223 18105 21235 18139
rect 21358 18136 21364 18148
rect 21319 18108 21364 18136
rect 21177 18099 21235 18105
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 7374 18068 7380 18080
rect 7335 18040 7380 18068
rect 7374 18028 7380 18040
rect 7432 18028 7438 18080
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 10226 18068 10232 18080
rect 9824 18040 10232 18068
rect 9824 18028 9830 18040
rect 10226 18028 10232 18040
rect 10284 18068 10290 18080
rect 10689 18071 10747 18077
rect 10689 18068 10701 18071
rect 10284 18040 10701 18068
rect 10284 18028 10290 18040
rect 10689 18037 10701 18040
rect 10735 18037 10747 18071
rect 11238 18068 11244 18080
rect 11199 18040 11244 18068
rect 10689 18031 10747 18037
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12713 18071 12771 18077
rect 12713 18068 12725 18071
rect 12492 18040 12725 18068
rect 12492 18028 12498 18040
rect 12713 18037 12725 18040
rect 12759 18037 12771 18071
rect 12713 18031 12771 18037
rect 13817 18071 13875 18077
rect 13817 18037 13829 18071
rect 13863 18068 13875 18071
rect 16482 18068 16488 18080
rect 13863 18040 16488 18068
rect 13863 18037 13875 18040
rect 13817 18031 13875 18037
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 17586 18068 17592 18080
rect 17547 18040 17592 18068
rect 17586 18028 17592 18040
rect 17644 18028 17650 18080
rect 17957 18071 18015 18077
rect 17957 18037 17969 18071
rect 18003 18068 18015 18071
rect 18509 18071 18567 18077
rect 18509 18068 18521 18071
rect 18003 18040 18521 18068
rect 18003 18037 18015 18040
rect 17957 18031 18015 18037
rect 18509 18037 18521 18040
rect 18555 18037 18567 18071
rect 18509 18031 18567 18037
rect 18969 18071 19027 18077
rect 18969 18037 18981 18071
rect 19015 18068 19027 18071
rect 19058 18068 19064 18080
rect 19015 18040 19064 18068
rect 19015 18037 19027 18040
rect 18969 18031 19027 18037
rect 19058 18028 19064 18040
rect 19116 18028 19122 18080
rect 19794 18028 19800 18080
rect 19852 18068 19858 18080
rect 19978 18068 19984 18080
rect 19852 18040 19984 18068
rect 19852 18028 19858 18040
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 3602 17864 3608 17876
rect 3563 17836 3608 17864
rect 3602 17824 3608 17836
rect 3660 17824 3666 17876
rect 5718 17864 5724 17876
rect 5679 17836 5724 17864
rect 5718 17824 5724 17836
rect 5776 17824 5782 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 7561 17867 7619 17873
rect 7561 17864 7573 17867
rect 7432 17836 7573 17864
rect 7432 17824 7438 17836
rect 7561 17833 7573 17836
rect 7607 17833 7619 17867
rect 7561 17827 7619 17833
rect 9582 17824 9588 17876
rect 9640 17864 9646 17876
rect 9861 17867 9919 17873
rect 9861 17864 9873 17867
rect 9640 17836 9873 17864
rect 9640 17824 9646 17836
rect 9861 17833 9873 17836
rect 9907 17833 9919 17867
rect 9861 17827 9919 17833
rect 10321 17867 10379 17873
rect 10321 17833 10333 17867
rect 10367 17864 10379 17867
rect 11238 17864 11244 17876
rect 10367 17836 11244 17864
rect 10367 17833 10379 17836
rect 10321 17827 10379 17833
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 18322 17864 18328 17876
rect 12406 17836 18328 17864
rect 1765 17799 1823 17805
rect 1765 17765 1777 17799
rect 1811 17796 1823 17799
rect 1811 17768 11744 17796
rect 1811 17765 1823 17768
rect 1765 17759 1823 17765
rect 3513 17731 3571 17737
rect 3513 17697 3525 17731
rect 3559 17728 3571 17731
rect 4249 17731 4307 17737
rect 4249 17728 4261 17731
rect 3559 17700 4261 17728
rect 3559 17697 3571 17700
rect 3513 17691 3571 17697
rect 4249 17697 4261 17700
rect 4295 17728 4307 17731
rect 7193 17731 7251 17737
rect 7193 17728 7205 17731
rect 4295 17700 7205 17728
rect 4295 17697 4307 17700
rect 4249 17691 4307 17697
rect 7193 17697 7205 17700
rect 7239 17728 7251 17731
rect 7742 17728 7748 17740
rect 7239 17700 7748 17728
rect 7239 17697 7251 17700
rect 7193 17691 7251 17697
rect 7742 17688 7748 17700
rect 7800 17688 7806 17740
rect 8478 17688 8484 17740
rect 8536 17728 8542 17740
rect 9122 17728 9128 17740
rect 8536 17700 9128 17728
rect 8536 17688 8542 17700
rect 9122 17688 9128 17700
rect 9180 17728 9186 17740
rect 9953 17731 10011 17737
rect 9953 17728 9965 17731
rect 9180 17700 9965 17728
rect 9180 17688 9186 17700
rect 9953 17697 9965 17700
rect 9999 17728 10011 17731
rect 10597 17731 10655 17737
rect 10597 17728 10609 17731
rect 9999 17700 10609 17728
rect 9999 17697 10011 17700
rect 9953 17691 10011 17697
rect 10597 17697 10609 17700
rect 10643 17697 10655 17731
rect 11716 17728 11744 17768
rect 12406 17728 12434 17836
rect 18322 17824 18328 17836
rect 18380 17864 18386 17876
rect 18509 17867 18567 17873
rect 18509 17864 18521 17867
rect 18380 17836 18521 17864
rect 18380 17824 18386 17836
rect 18509 17833 18521 17836
rect 18555 17833 18567 17867
rect 18509 17827 18567 17833
rect 19337 17867 19395 17873
rect 19337 17833 19349 17867
rect 19383 17864 19395 17867
rect 19702 17864 19708 17876
rect 19383 17836 19708 17864
rect 19383 17833 19395 17836
rect 19337 17827 19395 17833
rect 19702 17824 19708 17836
rect 19760 17824 19766 17876
rect 20254 17864 20260 17876
rect 20215 17836 20260 17864
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 17310 17756 17316 17808
rect 17368 17805 17374 17808
rect 17368 17799 17432 17805
rect 17368 17765 17386 17799
rect 17420 17765 17432 17799
rect 17368 17759 17432 17765
rect 17368 17756 17374 17759
rect 17586 17756 17592 17808
rect 17644 17796 17650 17808
rect 18785 17799 18843 17805
rect 18785 17796 18797 17799
rect 17644 17768 18797 17796
rect 17644 17756 17650 17768
rect 18785 17765 18797 17768
rect 18831 17765 18843 17799
rect 18785 17759 18843 17765
rect 11716 17700 12434 17728
rect 10597 17691 10655 17697
rect 16482 17688 16488 17740
rect 16540 17728 16546 17740
rect 19153 17731 19211 17737
rect 19153 17728 19165 17731
rect 16540 17700 19165 17728
rect 16540 17688 16546 17700
rect 19153 17697 19165 17700
rect 19199 17697 19211 17731
rect 19153 17691 19211 17697
rect 19613 17731 19671 17737
rect 19613 17697 19625 17731
rect 19659 17697 19671 17731
rect 20073 17731 20131 17737
rect 20073 17728 20085 17731
rect 19613 17691 19671 17697
rect 19812 17700 20085 17728
rect 3694 17660 3700 17672
rect 3655 17632 3700 17660
rect 3694 17620 3700 17632
rect 3752 17620 3758 17672
rect 5534 17620 5540 17672
rect 5592 17660 5598 17672
rect 6917 17663 6975 17669
rect 6917 17660 6929 17663
rect 5592 17632 6929 17660
rect 5592 17620 5598 17632
rect 6917 17629 6929 17632
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 7101 17663 7159 17669
rect 7101 17629 7113 17663
rect 7147 17660 7159 17663
rect 7650 17660 7656 17672
rect 7147 17632 7656 17660
rect 7147 17629 7159 17632
rect 7101 17623 7159 17629
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 9766 17660 9772 17672
rect 9727 17632 9772 17660
rect 9766 17620 9772 17632
rect 9824 17620 9830 17672
rect 17126 17660 17132 17672
rect 17087 17632 17132 17660
rect 17126 17620 17132 17632
rect 17184 17620 17190 17672
rect 18138 17620 18144 17672
rect 18196 17660 18202 17672
rect 19628 17660 19656 17691
rect 18196 17632 19656 17660
rect 18196 17620 18202 17632
rect 12161 17595 12219 17601
rect 12161 17561 12173 17595
rect 12207 17592 12219 17595
rect 12434 17592 12440 17604
rect 12207 17564 12440 17592
rect 12207 17561 12219 17564
rect 12161 17555 12219 17561
rect 12434 17552 12440 17564
rect 12492 17552 12498 17604
rect 19812 17601 19840 17700
rect 20073 17697 20085 17700
rect 20119 17697 20131 17731
rect 20622 17728 20628 17740
rect 20583 17700 20628 17728
rect 20073 17691 20131 17697
rect 20622 17688 20628 17700
rect 20680 17688 20686 17740
rect 20714 17688 20720 17740
rect 20772 17728 20778 17740
rect 21177 17731 21235 17737
rect 21177 17728 21189 17731
rect 20772 17700 21189 17728
rect 20772 17688 20778 17700
rect 21177 17697 21189 17700
rect 21223 17697 21235 17731
rect 21177 17691 21235 17697
rect 19797 17595 19855 17601
rect 19797 17561 19809 17595
rect 19843 17561 19855 17595
rect 20806 17592 20812 17604
rect 20767 17564 20812 17592
rect 19797 17555 19855 17561
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 21358 17592 21364 17604
rect 21319 17564 21364 17592
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 1670 17524 1676 17536
rect 1631 17496 1676 17524
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 3050 17484 3056 17536
rect 3108 17524 3114 17536
rect 3145 17527 3203 17533
rect 3145 17524 3157 17527
rect 3108 17496 3157 17524
rect 3108 17484 3114 17496
rect 3145 17493 3157 17496
rect 3191 17493 3203 17527
rect 3145 17487 3203 17493
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 7837 17527 7895 17533
rect 7837 17524 7849 17527
rect 7800 17496 7849 17524
rect 7800 17484 7806 17496
rect 7837 17493 7849 17496
rect 7883 17493 7895 17527
rect 7837 17487 7895 17493
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 1762 17320 1768 17332
rect 1723 17292 1768 17320
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 3510 17280 3516 17332
rect 3568 17320 3574 17332
rect 15473 17323 15531 17329
rect 3568 17292 15424 17320
rect 3568 17280 3574 17292
rect 4709 17255 4767 17261
rect 4709 17221 4721 17255
rect 4755 17252 4767 17255
rect 12989 17255 13047 17261
rect 4755 17224 12848 17252
rect 4755 17221 4767 17224
rect 4709 17215 4767 17221
rect 7466 17184 7472 17196
rect 7427 17156 7472 17184
rect 7466 17144 7472 17156
rect 7524 17144 7530 17196
rect 8478 17184 8484 17196
rect 8439 17156 8484 17184
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 11238 17144 11244 17196
rect 11296 17184 11302 17196
rect 11333 17187 11391 17193
rect 11333 17184 11345 17187
rect 11296 17156 11345 17184
rect 11296 17144 11302 17156
rect 11333 17153 11345 17156
rect 11379 17153 11391 17187
rect 11333 17147 11391 17153
rect 12437 17187 12495 17193
rect 12437 17153 12449 17187
rect 12483 17184 12495 17187
rect 12526 17184 12532 17196
rect 12483 17156 12532 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 3145 17119 3203 17125
rect 3145 17085 3157 17119
rect 3191 17116 3203 17119
rect 3878 17116 3884 17128
rect 3191 17088 3884 17116
rect 3191 17085 3203 17088
rect 3145 17079 3203 17085
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 4246 17076 4252 17128
rect 4304 17116 4310 17128
rect 4525 17119 4583 17125
rect 4525 17116 4537 17119
rect 4304 17088 4537 17116
rect 4304 17076 4310 17088
rect 4525 17085 4537 17088
rect 4571 17085 4583 17119
rect 4525 17079 4583 17085
rect 6086 17076 6092 17128
rect 6144 17116 6150 17128
rect 7653 17119 7711 17125
rect 7653 17116 7665 17119
rect 6144 17088 7665 17116
rect 6144 17076 6150 17088
rect 7653 17085 7665 17088
rect 7699 17085 7711 17119
rect 7653 17079 7711 17085
rect 7745 17119 7803 17125
rect 7745 17085 7757 17119
rect 7791 17116 7803 17119
rect 8496 17116 8524 17144
rect 7791 17088 8524 17116
rect 7791 17085 7803 17088
rect 7745 17079 7803 17085
rect 11146 17076 11152 17128
rect 11204 17116 11210 17128
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 11204 17088 11529 17116
rect 11204 17076 11210 17088
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 11609 17119 11667 17125
rect 11609 17085 11621 17119
rect 11655 17116 11667 17119
rect 11655 17088 12434 17116
rect 11655 17085 11667 17088
rect 11609 17079 11667 17085
rect 12406 17060 12434 17088
rect 2866 17048 2872 17060
rect 2924 17057 2930 17060
rect 2924 17051 2958 17057
rect 2810 17020 2872 17048
rect 2866 17008 2872 17020
rect 2946 17048 2958 17051
rect 3694 17048 3700 17060
rect 2946 17020 3700 17048
rect 2946 17017 2958 17020
rect 2924 17011 2958 17017
rect 2924 17008 2930 17011
rect 3694 17008 3700 17020
rect 3752 17008 3758 17060
rect 12406 17020 12440 17060
rect 12434 17008 12440 17020
rect 12492 17008 12498 17060
rect 12820 17048 12848 17224
rect 12989 17221 13001 17255
rect 13035 17252 13047 17255
rect 13035 17224 15332 17252
rect 13035 17221 13047 17224
rect 12989 17215 13047 17221
rect 14921 17187 14979 17193
rect 14921 17153 14933 17187
rect 14967 17184 14979 17187
rect 15194 17184 15200 17196
rect 14967 17156 15200 17184
rect 14967 17153 14979 17156
rect 14921 17147 14979 17153
rect 15194 17144 15200 17156
rect 15252 17144 15258 17196
rect 15105 17119 15163 17125
rect 15105 17085 15117 17119
rect 15151 17116 15163 17119
rect 15304 17116 15332 17224
rect 15396 17184 15424 17292
rect 15473 17289 15485 17323
rect 15519 17320 15531 17323
rect 18138 17320 18144 17332
rect 15519 17292 18144 17320
rect 15519 17289 15531 17292
rect 15473 17283 15531 17289
rect 18138 17280 18144 17292
rect 18196 17280 18202 17332
rect 19242 17320 19248 17332
rect 19203 17292 19248 17320
rect 19242 17280 19248 17292
rect 19300 17280 19306 17332
rect 20622 17320 20628 17332
rect 20583 17292 20628 17320
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 19702 17184 19708 17196
rect 15396 17156 19708 17184
rect 19702 17144 19708 17156
rect 19760 17144 19766 17196
rect 19058 17116 19064 17128
rect 15151 17088 15240 17116
rect 15304 17088 18920 17116
rect 19019 17088 19064 17116
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 15212 17048 15240 17088
rect 15749 17051 15807 17057
rect 15749 17048 15761 17051
rect 12820 17020 15148 17048
rect 15212 17020 15761 17048
rect 8113 16983 8171 16989
rect 8113 16949 8125 16983
rect 8159 16980 8171 16983
rect 8294 16980 8300 16992
rect 8159 16952 8300 16980
rect 8159 16949 8171 16952
rect 8113 16943 8171 16949
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 11977 16983 12035 16989
rect 11977 16949 11989 16983
rect 12023 16980 12035 16983
rect 12529 16983 12587 16989
rect 12529 16980 12541 16983
rect 12023 16952 12541 16980
rect 12023 16949 12035 16952
rect 11977 16943 12035 16949
rect 12529 16949 12541 16952
rect 12575 16949 12587 16983
rect 12529 16943 12587 16949
rect 12618 16940 12624 16992
rect 12676 16980 12682 16992
rect 12676 16952 12721 16980
rect 12676 16940 12682 16952
rect 14734 16940 14740 16992
rect 14792 16980 14798 16992
rect 15013 16983 15071 16989
rect 15013 16980 15025 16983
rect 14792 16952 15025 16980
rect 14792 16940 14798 16952
rect 15013 16949 15025 16952
rect 15059 16949 15071 16983
rect 15120 16980 15148 17020
rect 15749 17017 15761 17020
rect 15795 17017 15807 17051
rect 18892 17048 18920 17088
rect 19058 17076 19064 17088
rect 19116 17076 19122 17128
rect 19797 17119 19855 17125
rect 19797 17085 19809 17119
rect 19843 17085 19855 17119
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 19797 17079 19855 17085
rect 19996 17088 20821 17116
rect 19812 17048 19840 17079
rect 18892 17020 19840 17048
rect 15749 17011 15807 17017
rect 19426 16980 19432 16992
rect 15120 16952 19432 16980
rect 15013 16943 15071 16949
rect 19426 16940 19432 16952
rect 19484 16940 19490 16992
rect 19996 16989 20024 17088
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 20809 17079 20867 17085
rect 21174 17048 21180 17060
rect 21135 17020 21180 17048
rect 21174 17008 21180 17020
rect 21232 17008 21238 17060
rect 21361 17051 21419 17057
rect 21361 17017 21373 17051
rect 21407 17048 21419 17051
rect 21450 17048 21456 17060
rect 21407 17020 21456 17048
rect 21407 17017 21419 17020
rect 21361 17011 21419 17017
rect 21450 17008 21456 17020
rect 21508 17008 21514 17060
rect 19981 16983 20039 16989
rect 19981 16949 19993 16983
rect 20027 16949 20039 16983
rect 19981 16943 20039 16949
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 3050 16776 3056 16788
rect 3011 16748 3056 16776
rect 3050 16736 3056 16748
rect 3108 16736 3114 16788
rect 3510 16776 3516 16788
rect 3471 16748 3516 16776
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 5905 16779 5963 16785
rect 5905 16745 5917 16779
rect 5951 16745 5963 16779
rect 5905 16739 5963 16745
rect 4798 16717 4804 16720
rect 4792 16671 4804 16717
rect 4856 16708 4862 16720
rect 5920 16708 5948 16739
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 9217 16779 9275 16785
rect 9217 16776 9229 16779
rect 8352 16748 9229 16776
rect 8352 16736 8358 16748
rect 9217 16745 9229 16748
rect 9263 16745 9275 16779
rect 9217 16739 9275 16745
rect 9677 16779 9735 16785
rect 9677 16745 9689 16779
rect 9723 16776 9735 16779
rect 10597 16779 10655 16785
rect 9723 16748 10456 16776
rect 9723 16745 9735 16748
rect 9677 16739 9735 16745
rect 7466 16708 7472 16720
rect 4856 16680 4892 16708
rect 5920 16680 7472 16708
rect 4798 16668 4804 16671
rect 4856 16668 4862 16680
rect 7466 16668 7472 16680
rect 7524 16717 7530 16720
rect 7524 16711 7588 16717
rect 7524 16677 7542 16711
rect 7576 16677 7588 16711
rect 7524 16671 7588 16677
rect 7524 16668 7530 16671
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16640 3203 16643
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3191 16612 3801 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 3789 16609 3801 16612
rect 3835 16609 3847 16643
rect 3789 16603 3847 16609
rect 3878 16600 3884 16652
rect 3936 16640 3942 16652
rect 4525 16643 4583 16649
rect 4525 16640 4537 16643
rect 3936 16612 4537 16640
rect 3936 16600 3942 16612
rect 4525 16609 4537 16612
rect 4571 16640 4583 16643
rect 5258 16640 5264 16652
rect 4571 16612 5264 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 5258 16600 5264 16612
rect 5316 16640 5322 16652
rect 7282 16640 7288 16652
rect 5316 16612 7288 16640
rect 5316 16600 5322 16612
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 10428 16649 10456 16748
rect 10597 16745 10609 16779
rect 10643 16745 10655 16779
rect 10597 16739 10655 16745
rect 12161 16779 12219 16785
rect 12161 16745 12173 16779
rect 12207 16776 12219 16779
rect 12618 16776 12624 16788
rect 12207 16748 12624 16776
rect 12207 16745 12219 16748
rect 12161 16739 12219 16745
rect 10612 16708 10640 16739
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 14274 16736 14280 16788
rect 14332 16776 14338 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 14332 16748 14381 16776
rect 14332 16736 14338 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 14369 16739 14427 16745
rect 14734 16736 14740 16788
rect 14792 16776 14798 16788
rect 14829 16779 14887 16785
rect 14829 16776 14841 16779
rect 14792 16748 14841 16776
rect 14792 16736 14798 16748
rect 14829 16745 14841 16748
rect 14875 16745 14887 16779
rect 14829 16739 14887 16745
rect 18877 16779 18935 16785
rect 18877 16745 18889 16779
rect 18923 16776 18935 16779
rect 19334 16776 19340 16788
rect 18923 16748 19340 16776
rect 18923 16745 18935 16748
rect 18877 16739 18935 16745
rect 19334 16736 19340 16748
rect 19392 16736 19398 16788
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 20349 16779 20407 16785
rect 19484 16748 20300 16776
rect 19484 16736 19490 16748
rect 20272 16708 20300 16748
rect 20349 16745 20361 16779
rect 20395 16776 20407 16779
rect 20714 16776 20720 16788
rect 20395 16748 20720 16776
rect 20395 16745 20407 16748
rect 20349 16739 20407 16745
rect 20714 16736 20720 16748
rect 20772 16736 20778 16788
rect 20809 16779 20867 16785
rect 20809 16745 20821 16779
rect 20855 16776 20867 16779
rect 21174 16776 21180 16788
rect 20855 16748 21180 16776
rect 20855 16745 20867 16748
rect 20809 16739 20867 16745
rect 21174 16736 21180 16748
rect 21232 16736 21238 16788
rect 10612 16680 20208 16708
rect 20272 16680 20668 16708
rect 9309 16643 9367 16649
rect 9309 16609 9321 16643
rect 9355 16640 9367 16643
rect 9953 16643 10011 16649
rect 9953 16640 9965 16643
rect 9355 16612 9965 16640
rect 9355 16609 9367 16612
rect 9309 16603 9367 16609
rect 9953 16609 9965 16612
rect 9999 16609 10011 16643
rect 9953 16603 10011 16609
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16609 10471 16643
rect 10413 16603 10471 16609
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16609 12495 16643
rect 12437 16603 12495 16609
rect 1762 16532 1768 16584
rect 1820 16572 1826 16584
rect 2869 16575 2927 16581
rect 2869 16572 2881 16575
rect 1820 16544 2881 16572
rect 1820 16532 1826 16544
rect 2869 16541 2881 16544
rect 2915 16541 2927 16575
rect 9125 16575 9183 16581
rect 9125 16572 9137 16575
rect 2869 16535 2927 16541
rect 8680 16544 9137 16572
rect 8680 16513 8708 16544
rect 9125 16541 9137 16544
rect 9171 16572 9183 16575
rect 9398 16572 9404 16584
rect 9171 16544 9404 16572
rect 9171 16541 9183 16544
rect 9125 16535 9183 16541
rect 9398 16532 9404 16544
rect 9456 16532 9462 16584
rect 8665 16507 8723 16513
rect 8665 16473 8677 16507
rect 8711 16473 8723 16507
rect 8665 16467 8723 16473
rect 12452 16436 12480 16603
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 12693 16643 12751 16649
rect 12693 16640 12705 16643
rect 12584 16612 12705 16640
rect 12584 16600 12590 16612
rect 12693 16609 12705 16612
rect 12739 16609 12751 16643
rect 12693 16603 12751 16609
rect 14461 16643 14519 16649
rect 14461 16609 14473 16643
rect 14507 16640 14519 16643
rect 14642 16640 14648 16652
rect 14507 16612 14648 16640
rect 14507 16609 14519 16612
rect 14461 16603 14519 16609
rect 14642 16600 14648 16612
rect 14700 16600 14706 16652
rect 15197 16643 15255 16649
rect 15197 16640 15209 16643
rect 15120 16612 15209 16640
rect 14274 16572 14280 16584
rect 13832 16544 14280 16572
rect 13832 16513 13860 16544
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 14550 16532 14556 16584
rect 14608 16572 14614 16584
rect 15120 16572 15148 16612
rect 15197 16609 15209 16612
rect 15243 16609 15255 16643
rect 15197 16603 15255 16609
rect 15286 16600 15292 16652
rect 15344 16640 15350 16652
rect 15464 16643 15522 16649
rect 15464 16640 15476 16643
rect 15344 16612 15476 16640
rect 15344 16600 15350 16612
rect 15464 16609 15476 16612
rect 15510 16640 15522 16643
rect 15930 16640 15936 16652
rect 15510 16612 15936 16640
rect 15510 16609 15522 16612
rect 15464 16603 15522 16609
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 18690 16640 18696 16652
rect 18651 16612 18696 16640
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 19702 16640 19708 16652
rect 19663 16612 19708 16640
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 20180 16649 20208 16680
rect 20640 16649 20668 16680
rect 20165 16643 20223 16649
rect 20165 16609 20177 16643
rect 20211 16609 20223 16643
rect 20165 16603 20223 16609
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16609 20683 16643
rect 21174 16640 21180 16652
rect 21135 16612 21180 16640
rect 20625 16603 20683 16609
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 21358 16640 21364 16652
rect 21319 16612 21364 16640
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 14608 16544 15148 16572
rect 14608 16532 14614 16544
rect 13817 16507 13875 16513
rect 13817 16473 13829 16507
rect 13863 16473 13875 16507
rect 13817 16467 13875 16473
rect 14550 16436 14556 16448
rect 12452 16408 14556 16436
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 16574 16436 16580 16448
rect 16535 16408 16580 16436
rect 16574 16396 16580 16408
rect 16632 16396 16638 16448
rect 19889 16439 19947 16445
rect 19889 16405 19901 16439
rect 19935 16436 19947 16439
rect 20254 16436 20260 16448
rect 19935 16408 20260 16436
rect 19935 16405 19947 16408
rect 19889 16399 19947 16405
rect 20254 16396 20260 16408
rect 20312 16396 20318 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 4893 16235 4951 16241
rect 4893 16201 4905 16235
rect 4939 16232 4951 16235
rect 5534 16232 5540 16244
rect 4939 16204 5540 16232
rect 4939 16201 4951 16204
rect 4893 16195 4951 16201
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 10689 16235 10747 16241
rect 10689 16201 10701 16235
rect 10735 16232 10747 16235
rect 11238 16232 11244 16244
rect 10735 16204 11244 16232
rect 10735 16201 10747 16204
rect 10689 16195 10747 16201
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 12345 16235 12403 16241
rect 12345 16201 12357 16235
rect 12391 16232 12403 16235
rect 12526 16232 12532 16244
rect 12391 16204 12532 16232
rect 12391 16201 12403 16204
rect 12345 16195 12403 16201
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 15930 16232 15936 16244
rect 15891 16204 15936 16232
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 16666 16192 16672 16244
rect 16724 16232 16730 16244
rect 17405 16235 17463 16241
rect 17405 16232 17417 16235
rect 16724 16204 17417 16232
rect 16724 16192 16730 16204
rect 17405 16201 17417 16204
rect 17451 16232 17463 16235
rect 17586 16232 17592 16244
rect 17451 16204 17592 16232
rect 17451 16201 17463 16204
rect 17405 16195 17463 16201
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 18509 16235 18567 16241
rect 18509 16201 18521 16235
rect 18555 16232 18567 16235
rect 18690 16232 18696 16244
rect 18555 16204 18696 16232
rect 18555 16201 18567 16204
rect 18509 16195 18567 16201
rect 18690 16192 18696 16204
rect 18748 16192 18754 16244
rect 20073 16235 20131 16241
rect 20073 16201 20085 16235
rect 20119 16232 20131 16235
rect 20162 16232 20168 16244
rect 20119 16204 20168 16232
rect 20119 16201 20131 16204
rect 20073 16195 20131 16201
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 21174 16232 21180 16244
rect 20855 16204 21180 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 6273 16099 6331 16105
rect 6273 16065 6285 16099
rect 6319 16096 6331 16099
rect 7282 16096 7288 16108
rect 6319 16068 7288 16096
rect 6319 16065 6331 16068
rect 6273 16059 6331 16065
rect 7282 16056 7288 16068
rect 7340 16056 7346 16108
rect 10962 16096 10968 16108
rect 10923 16068 10968 16096
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 14550 16096 14556 16108
rect 14511 16068 14556 16096
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 16485 16099 16543 16105
rect 16485 16065 16497 16099
rect 16531 16096 16543 16099
rect 16574 16096 16580 16108
rect 16531 16068 16580 16096
rect 16531 16065 16543 16068
rect 16485 16059 16543 16065
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 17954 16096 17960 16108
rect 17915 16068 17960 16096
rect 17954 16056 17960 16068
rect 18012 16056 18018 16108
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 9309 16031 9367 16037
rect 9309 16028 9321 16031
rect 7524 16000 9321 16028
rect 7524 15988 7530 16000
rect 9309 15997 9321 16000
rect 9355 15997 9367 16031
rect 9309 15991 9367 15997
rect 9398 15988 9404 16040
rect 9456 16028 9462 16040
rect 11238 16037 11244 16040
rect 9565 16031 9623 16037
rect 9565 16028 9577 16031
rect 9456 16000 9577 16028
rect 9456 15988 9462 16000
rect 9565 15997 9577 16000
rect 9611 15997 9623 16031
rect 11232 16028 11244 16037
rect 11199 16000 11244 16028
rect 9565 15991 9623 15997
rect 11232 15991 11244 16000
rect 11238 15988 11244 15991
rect 11296 15988 11302 16040
rect 16114 15988 16120 16040
rect 16172 16028 16178 16040
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 16172 16000 19901 16028
rect 16172 15988 16178 16000
rect 19889 15997 19901 16000
rect 19935 15997 19947 16031
rect 19889 15991 19947 15997
rect 20254 15988 20260 16040
rect 20312 16028 20318 16040
rect 20625 16031 20683 16037
rect 20625 16028 20637 16031
rect 20312 16000 20637 16028
rect 20312 15988 20318 16000
rect 20625 15997 20637 16000
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 6086 15969 6092 15972
rect 6028 15963 6092 15969
rect 6028 15929 6040 15963
rect 6074 15929 6092 15963
rect 6028 15923 6092 15929
rect 6086 15920 6092 15923
rect 6144 15920 6150 15972
rect 14274 15920 14280 15972
rect 14332 15960 14338 15972
rect 14798 15963 14856 15969
rect 14798 15960 14810 15963
rect 14332 15932 14810 15960
rect 14332 15920 14338 15932
rect 14798 15929 14810 15932
rect 14844 15929 14856 15963
rect 14798 15923 14856 15929
rect 16577 15963 16635 15969
rect 16577 15929 16589 15963
rect 16623 15960 16635 15963
rect 16758 15960 16764 15972
rect 16623 15932 16764 15960
rect 16623 15929 16635 15932
rect 16577 15923 16635 15929
rect 16758 15920 16764 15932
rect 16816 15920 16822 15972
rect 18049 15963 18107 15969
rect 18049 15960 18061 15963
rect 17052 15932 18061 15960
rect 16666 15892 16672 15904
rect 16627 15864 16672 15892
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 17052 15901 17080 15932
rect 18049 15929 18061 15932
rect 18095 15929 18107 15963
rect 18049 15923 18107 15929
rect 20806 15920 20812 15972
rect 20864 15960 20870 15972
rect 21177 15963 21235 15969
rect 21177 15960 21189 15963
rect 20864 15932 21189 15960
rect 20864 15920 20870 15932
rect 21177 15929 21189 15932
rect 21223 15929 21235 15963
rect 21358 15960 21364 15972
rect 21319 15932 21364 15960
rect 21177 15923 21235 15929
rect 21358 15920 21364 15932
rect 21416 15920 21422 15972
rect 17037 15895 17095 15901
rect 17037 15861 17049 15895
rect 17083 15861 17095 15895
rect 17037 15855 17095 15861
rect 18141 15895 18199 15901
rect 18141 15861 18153 15895
rect 18187 15892 18199 15895
rect 18785 15895 18843 15901
rect 18785 15892 18797 15895
rect 18187 15864 18797 15892
rect 18187 15861 18199 15864
rect 18141 15855 18199 15861
rect 18785 15861 18797 15864
rect 18831 15861 18843 15895
rect 18785 15855 18843 15861
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 2866 15648 2872 15700
rect 2924 15688 2930 15700
rect 3237 15691 3295 15697
rect 3237 15688 3249 15691
rect 2924 15660 3249 15688
rect 2924 15648 2930 15660
rect 3237 15657 3249 15660
rect 3283 15657 3295 15691
rect 3237 15651 3295 15657
rect 7837 15691 7895 15697
rect 7837 15657 7849 15691
rect 7883 15688 7895 15691
rect 16114 15688 16120 15700
rect 7883 15660 16120 15688
rect 7883 15657 7895 15660
rect 7837 15651 7895 15657
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 17954 15648 17960 15700
rect 18012 15688 18018 15700
rect 18509 15691 18567 15697
rect 18509 15688 18521 15691
rect 18012 15660 18521 15688
rect 18012 15648 18018 15660
rect 18509 15657 18521 15660
rect 18555 15657 18567 15691
rect 20806 15688 20812 15700
rect 20767 15660 20812 15688
rect 18509 15651 18567 15657
rect 20806 15648 20812 15660
rect 20864 15648 20870 15700
rect 3878 15620 3884 15632
rect 1872 15592 3884 15620
rect 1872 15561 1900 15592
rect 3878 15580 3884 15592
rect 3936 15580 3942 15632
rect 8849 15623 8907 15629
rect 8849 15589 8861 15623
rect 8895 15620 8907 15623
rect 10962 15620 10968 15632
rect 8895 15592 10968 15620
rect 8895 15589 8907 15592
rect 8849 15583 8907 15589
rect 10962 15580 10968 15592
rect 11020 15580 11026 15632
rect 12406 15592 20024 15620
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15521 1915 15555
rect 1857 15515 1915 15521
rect 2124 15555 2182 15561
rect 2124 15521 2136 15555
rect 2170 15552 2182 15555
rect 2498 15552 2504 15564
rect 2170 15524 2504 15552
rect 2170 15521 2182 15524
rect 2124 15515 2182 15521
rect 2498 15512 2504 15524
rect 2556 15512 2562 15564
rect 7469 15555 7527 15561
rect 7469 15521 7481 15555
rect 7515 15552 7527 15555
rect 8113 15555 8171 15561
rect 8113 15552 8125 15555
rect 7515 15524 8125 15552
rect 7515 15521 7527 15524
rect 7469 15515 7527 15521
rect 8113 15521 8125 15524
rect 8159 15521 8171 15555
rect 8113 15515 8171 15521
rect 8757 15555 8815 15561
rect 8757 15521 8769 15555
rect 8803 15552 8815 15555
rect 9306 15552 9312 15564
rect 8803 15524 9312 15552
rect 8803 15521 8815 15524
rect 8757 15515 8815 15521
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 6086 15444 6092 15496
rect 6144 15484 6150 15496
rect 7193 15487 7251 15493
rect 7193 15484 7205 15487
rect 6144 15456 7205 15484
rect 6144 15444 6150 15456
rect 7193 15453 7205 15456
rect 7239 15453 7251 15487
rect 7193 15447 7251 15453
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15484 7435 15487
rect 7742 15484 7748 15496
rect 7423 15456 7748 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 4798 15376 4804 15428
rect 4856 15416 4862 15428
rect 12406 15416 12434 15592
rect 16574 15512 16580 15564
rect 16632 15552 16638 15564
rect 19996 15561 20024 15592
rect 20346 15580 20352 15632
rect 20404 15620 20410 15632
rect 21177 15623 21235 15629
rect 21177 15620 21189 15623
rect 20404 15592 21189 15620
rect 20404 15580 20410 15592
rect 21177 15589 21189 15592
rect 21223 15589 21235 15623
rect 21177 15583 21235 15589
rect 17385 15555 17443 15561
rect 17385 15552 17397 15555
rect 16632 15524 17397 15552
rect 16632 15512 16638 15524
rect 17385 15521 17397 15524
rect 17431 15521 17443 15555
rect 17385 15515 17443 15521
rect 19981 15555 20039 15561
rect 19981 15521 19993 15555
rect 20027 15521 20039 15555
rect 20625 15555 20683 15561
rect 20625 15552 20637 15555
rect 19981 15515 20039 15521
rect 20180 15524 20637 15552
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 17126 15484 17132 15496
rect 14608 15456 17132 15484
rect 14608 15444 14614 15456
rect 17126 15444 17132 15456
rect 17184 15444 17190 15496
rect 20180 15425 20208 15524
rect 20625 15521 20637 15524
rect 20671 15521 20683 15555
rect 20625 15515 20683 15521
rect 4856 15388 12434 15416
rect 20165 15419 20223 15425
rect 4856 15376 4862 15388
rect 20165 15385 20177 15419
rect 20211 15385 20223 15419
rect 21358 15416 21364 15428
rect 21319 15388 21364 15416
rect 20165 15379 20223 15385
rect 21358 15376 21364 15388
rect 21416 15376 21422 15428
rect 7282 15308 7288 15360
rect 7340 15348 7346 15360
rect 8573 15351 8631 15357
rect 8573 15348 8585 15351
rect 7340 15320 8585 15348
rect 7340 15308 7346 15320
rect 8573 15317 8585 15320
rect 8619 15348 8631 15351
rect 8849 15351 8907 15357
rect 8849 15348 8861 15351
rect 8619 15320 8861 15348
rect 8619 15317 8631 15320
rect 8573 15311 8631 15317
rect 8849 15317 8861 15320
rect 8895 15317 8907 15351
rect 9122 15348 9128 15360
rect 9035 15320 9128 15348
rect 8849 15311 8907 15317
rect 9122 15308 9128 15320
rect 9180 15348 9186 15360
rect 9582 15348 9588 15360
rect 9180 15320 9588 15348
rect 9180 15308 9186 15320
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 14642 15308 14648 15360
rect 14700 15348 14706 15360
rect 14921 15351 14979 15357
rect 14921 15348 14933 15351
rect 14700 15320 14933 15348
rect 14700 15308 14706 15320
rect 14921 15317 14933 15320
rect 14967 15317 14979 15351
rect 14921 15311 14979 15317
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 4798 15144 4804 15156
rect 4759 15116 4804 15144
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 6086 15144 6092 15156
rect 6047 15116 6092 15144
rect 6086 15104 6092 15116
rect 6144 15104 6150 15156
rect 7742 15144 7748 15156
rect 7703 15116 7748 15144
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 14734 15144 14740 15156
rect 14608 15116 14740 15144
rect 14608 15104 14614 15116
rect 14734 15104 14740 15116
rect 14792 15104 14798 15156
rect 20346 15144 20352 15156
rect 20307 15116 20352 15144
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 7558 15036 7564 15088
rect 7616 15076 7622 15088
rect 7616 15048 8432 15076
rect 7616 15036 7622 15048
rect 2498 14968 2504 15020
rect 2556 15008 2562 15020
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 2556 14980 4169 15008
rect 2556 14968 2562 14980
rect 4157 14977 4169 14980
rect 4203 14977 4215 15011
rect 8202 15008 8208 15020
rect 8163 14980 8208 15008
rect 4157 14971 4215 14977
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 14977 8355 15011
rect 8297 14971 8355 14977
rect 7466 14940 7472 14952
rect 7427 14912 7472 14940
rect 7466 14900 7472 14912
rect 7524 14900 7530 14952
rect 8312 14940 8340 14971
rect 8128 14912 8340 14940
rect 4433 14875 4491 14881
rect 4433 14841 4445 14875
rect 4479 14872 4491 14875
rect 5077 14875 5135 14881
rect 5077 14872 5089 14875
rect 4479 14844 5089 14872
rect 4479 14841 4491 14844
rect 4433 14835 4491 14841
rect 5077 14841 5089 14844
rect 5123 14841 5135 14875
rect 5077 14835 5135 14841
rect 7190 14832 7196 14884
rect 7248 14881 7254 14884
rect 7248 14872 7260 14881
rect 8128 14872 8156 14912
rect 7248 14844 8156 14872
rect 8404 14872 8432 15048
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 15008 12587 15011
rect 13998 15008 14004 15020
rect 12575 14980 14004 15008
rect 12575 14977 12587 14980
rect 12529 14971 12587 14977
rect 13998 14968 14004 14980
rect 14056 14968 14062 15020
rect 17126 14968 17132 15020
rect 17184 15008 17190 15020
rect 17773 15011 17831 15017
rect 17773 15008 17785 15011
rect 17184 14980 17785 15008
rect 17184 14968 17190 14980
rect 17773 14977 17785 14980
rect 17819 14977 17831 15011
rect 17773 14971 17831 14977
rect 9493 14943 9551 14949
rect 9493 14909 9505 14943
rect 9539 14940 9551 14943
rect 11054 14940 11060 14952
rect 9539 14912 11060 14940
rect 9539 14909 9551 14912
rect 9493 14903 9551 14909
rect 11054 14900 11060 14912
rect 11112 14900 11118 14952
rect 14550 14940 14556 14952
rect 14511 14912 14556 14940
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 20162 14940 20168 14952
rect 20123 14912 20168 14940
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 20530 14900 20536 14952
rect 20588 14940 20594 14952
rect 20625 14943 20683 14949
rect 20625 14940 20637 14943
rect 20588 14912 20637 14940
rect 20588 14900 20594 14912
rect 20625 14909 20637 14912
rect 20671 14909 20683 14943
rect 20625 14903 20683 14909
rect 17862 14872 17868 14884
rect 8404 14844 17868 14872
rect 7248 14835 7260 14844
rect 7248 14832 7254 14835
rect 17862 14832 17868 14844
rect 17920 14832 17926 14884
rect 17954 14832 17960 14884
rect 18012 14881 18018 14884
rect 18012 14875 18076 14881
rect 18012 14841 18030 14875
rect 18064 14841 18076 14875
rect 21177 14875 21235 14881
rect 21177 14872 21189 14875
rect 18012 14835 18076 14841
rect 20824 14844 21189 14872
rect 18012 14832 18018 14835
rect 4246 14764 4252 14816
rect 4304 14804 4310 14816
rect 4341 14807 4399 14813
rect 4341 14804 4353 14807
rect 4304 14776 4353 14804
rect 4304 14764 4310 14776
rect 4341 14773 4353 14776
rect 4387 14773 4399 14807
rect 4341 14767 4399 14773
rect 8113 14807 8171 14813
rect 8113 14773 8125 14807
rect 8159 14804 8171 14807
rect 8294 14804 8300 14816
rect 8159 14776 8300 14804
rect 8159 14773 8171 14776
rect 8113 14767 8171 14773
rect 8294 14764 8300 14776
rect 8352 14804 8358 14816
rect 9122 14804 9128 14816
rect 8352 14776 9128 14804
rect 8352 14764 8358 14776
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9306 14804 9312 14816
rect 9267 14776 9312 14804
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 12618 14804 12624 14816
rect 12579 14776 12624 14804
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 13078 14804 13084 14816
rect 12768 14776 12813 14804
rect 13039 14776 13084 14804
rect 12768 14764 12774 14776
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 13170 14764 13176 14816
rect 13228 14804 13234 14816
rect 18598 14804 18604 14816
rect 13228 14776 18604 14804
rect 13228 14764 13234 14776
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 19150 14804 19156 14816
rect 19111 14776 19156 14804
rect 19150 14764 19156 14776
rect 19208 14764 19214 14816
rect 20824 14813 20852 14844
rect 21177 14841 21189 14844
rect 21223 14841 21235 14875
rect 21358 14872 21364 14884
rect 21319 14844 21364 14872
rect 21177 14835 21235 14841
rect 21358 14832 21364 14844
rect 21416 14832 21422 14884
rect 20809 14807 20867 14813
rect 20809 14773 20821 14807
rect 20855 14773 20867 14807
rect 20809 14767 20867 14773
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 2498 14600 2504 14612
rect 2459 14572 2504 14600
rect 2498 14560 2504 14572
rect 2556 14560 2562 14612
rect 4246 14600 4252 14612
rect 4207 14572 4252 14600
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 4709 14603 4767 14609
rect 4709 14569 4721 14603
rect 4755 14600 4767 14603
rect 4982 14600 4988 14612
rect 4755 14572 4988 14600
rect 4755 14569 4767 14572
rect 4709 14563 4767 14569
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 8570 14600 8576 14612
rect 8531 14572 8576 14600
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 9677 14603 9735 14609
rect 9677 14569 9689 14603
rect 9723 14569 9735 14603
rect 9677 14563 9735 14569
rect 12161 14603 12219 14609
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 12250 14600 12256 14612
rect 12207 14572 12256 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 4617 14535 4675 14541
rect 4617 14501 4629 14535
rect 4663 14532 4675 14535
rect 5353 14535 5411 14541
rect 5353 14532 5365 14535
rect 4663 14504 5365 14532
rect 4663 14501 4675 14504
rect 4617 14495 4675 14501
rect 5353 14501 5365 14504
rect 5399 14532 5411 14535
rect 8294 14532 8300 14544
rect 5399 14504 8300 14532
rect 5399 14501 5411 14504
rect 5353 14495 5411 14501
rect 8294 14492 8300 14504
rect 8352 14492 8358 14544
rect 9692 14532 9720 14563
rect 12250 14560 12256 14572
rect 12308 14560 12314 14612
rect 12618 14600 12624 14612
rect 12579 14572 12624 14600
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 13078 14560 13084 14612
rect 13136 14600 13142 14612
rect 15565 14603 15623 14609
rect 15565 14600 15577 14603
rect 13136 14572 15577 14600
rect 13136 14560 13142 14572
rect 15565 14569 15577 14572
rect 15611 14569 15623 14603
rect 15565 14563 15623 14569
rect 17862 14560 17868 14612
rect 17920 14600 17926 14612
rect 17957 14603 18015 14609
rect 17957 14600 17969 14603
rect 17920 14572 17969 14600
rect 17920 14560 17926 14572
rect 17957 14569 17969 14572
rect 18003 14569 18015 14603
rect 17957 14563 18015 14569
rect 18417 14603 18475 14609
rect 18417 14569 18429 14603
rect 18463 14600 18475 14603
rect 18969 14603 19027 14609
rect 18969 14600 18981 14603
rect 18463 14572 18981 14600
rect 18463 14569 18475 14572
rect 18417 14563 18475 14569
rect 18969 14569 18981 14572
rect 19015 14569 19027 14603
rect 18969 14563 19027 14569
rect 20809 14603 20867 14609
rect 20809 14569 20821 14603
rect 20855 14600 20867 14603
rect 20898 14600 20904 14612
rect 20855 14572 20904 14600
rect 20855 14569 20867 14572
rect 20809 14563 20867 14569
rect 20898 14560 20904 14572
rect 20956 14560 20962 14612
rect 20162 14532 20168 14544
rect 9692 14504 20168 14532
rect 20162 14492 20168 14504
rect 20220 14492 20226 14544
rect 3625 14467 3683 14473
rect 3625 14433 3637 14467
rect 3671 14464 3683 14467
rect 4154 14464 4160 14476
rect 3671 14436 4160 14464
rect 3671 14433 3683 14436
rect 3625 14427 3683 14433
rect 4154 14424 4160 14436
rect 4212 14464 4218 14476
rect 8665 14467 8723 14473
rect 4212 14436 4844 14464
rect 4212 14424 4218 14436
rect 3878 14396 3884 14408
rect 3839 14368 3884 14396
rect 3878 14356 3884 14368
rect 3936 14356 3942 14408
rect 4816 14405 4844 14436
rect 8665 14433 8677 14467
rect 8711 14433 8723 14467
rect 9490 14464 9496 14476
rect 9451 14436 9496 14464
rect 8665 14427 8723 14433
rect 4801 14399 4859 14405
rect 4801 14365 4813 14399
rect 4847 14365 4859 14399
rect 8478 14396 8484 14408
rect 8439 14368 8484 14396
rect 4801 14359 4859 14365
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 8680 14396 8708 14427
rect 9490 14424 9496 14436
rect 9548 14424 9554 14476
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 12253 14467 12311 14473
rect 12253 14464 12265 14467
rect 9640 14436 12265 14464
rect 9640 14424 9646 14436
rect 12253 14433 12265 14436
rect 12299 14464 12311 14467
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12299 14436 12817 14464
rect 12299 14433 12311 14436
rect 12253 14427 12311 14433
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 13998 14424 14004 14476
rect 14056 14464 14062 14476
rect 14746 14467 14804 14473
rect 14746 14464 14758 14467
rect 14056 14436 14758 14464
rect 14056 14424 14062 14436
rect 14746 14433 14758 14436
rect 14792 14433 14804 14467
rect 14746 14427 14804 14433
rect 14918 14424 14924 14476
rect 14976 14464 14982 14476
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 14976 14436 15025 14464
rect 14976 14424 14982 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15654 14464 15660 14476
rect 15615 14436 15660 14464
rect 15013 14427 15071 14433
rect 15654 14424 15660 14436
rect 15712 14424 15718 14476
rect 18049 14467 18107 14473
rect 18049 14433 18061 14467
rect 18095 14464 18107 14467
rect 18598 14464 18604 14476
rect 18095 14436 18604 14464
rect 18095 14433 18107 14436
rect 18049 14427 18107 14433
rect 18598 14424 18604 14436
rect 18656 14424 18662 14476
rect 19061 14467 19119 14473
rect 19061 14433 19073 14467
rect 19107 14464 19119 14467
rect 19334 14464 19340 14476
rect 19107 14436 19340 14464
rect 19107 14433 19119 14436
rect 19061 14427 19119 14433
rect 19334 14424 19340 14436
rect 19392 14424 19398 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19444 14436 19993 14464
rect 9674 14396 9680 14408
rect 8680 14368 9680 14396
rect 9674 14356 9680 14368
rect 9732 14396 9738 14408
rect 9953 14399 10011 14405
rect 9953 14396 9965 14399
rect 9732 14368 9965 14396
rect 9732 14356 9738 14368
rect 9953 14365 9965 14368
rect 9999 14365 10011 14399
rect 9953 14359 10011 14365
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14396 12127 14399
rect 12158 14396 12164 14408
rect 12115 14368 12164 14396
rect 12115 14365 12127 14368
rect 12069 14359 12127 14365
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14365 15439 14399
rect 15381 14359 15439 14365
rect 17865 14399 17923 14405
rect 17865 14365 17877 14399
rect 17911 14365 17923 14399
rect 17865 14359 17923 14365
rect 12250 14288 12256 14340
rect 12308 14328 12314 14340
rect 12308 14300 13676 14328
rect 12308 14288 12314 14300
rect 9030 14260 9036 14272
rect 8991 14232 9036 14260
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 12805 14263 12863 14269
rect 12805 14229 12817 14263
rect 12851 14260 12863 14263
rect 12989 14263 13047 14269
rect 12989 14260 13001 14263
rect 12851 14232 13001 14260
rect 12851 14229 12863 14232
rect 12805 14223 12863 14229
rect 12989 14229 13001 14232
rect 13035 14260 13047 14263
rect 13354 14260 13360 14272
rect 13035 14232 13360 14260
rect 13035 14229 13047 14232
rect 12989 14223 13047 14229
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 13648 14269 13676 14300
rect 13633 14263 13691 14269
rect 13633 14229 13645 14263
rect 13679 14260 13691 14263
rect 15396 14260 15424 14359
rect 17880 14328 17908 14359
rect 18690 14356 18696 14408
rect 18748 14396 18754 14408
rect 18785 14399 18843 14405
rect 18785 14396 18797 14399
rect 18748 14368 18797 14396
rect 18748 14356 18754 14368
rect 18785 14365 18797 14368
rect 18831 14365 18843 14399
rect 18785 14359 18843 14365
rect 18046 14328 18052 14340
rect 17880 14300 18052 14328
rect 18046 14288 18052 14300
rect 18104 14328 18110 14340
rect 19150 14328 19156 14340
rect 18104 14300 19156 14328
rect 18104 14288 18110 14300
rect 19150 14288 19156 14300
rect 19208 14288 19214 14340
rect 19444 14337 19472 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 20625 14467 20683 14473
rect 20625 14464 20637 14467
rect 19981 14427 20039 14433
rect 20180 14436 20637 14464
rect 20180 14337 20208 14436
rect 20625 14433 20637 14436
rect 20671 14433 20683 14467
rect 20625 14427 20683 14433
rect 21085 14467 21143 14473
rect 21085 14433 21097 14467
rect 21131 14433 21143 14467
rect 21085 14427 21143 14433
rect 20438 14356 20444 14408
rect 20496 14396 20502 14408
rect 21100 14396 21128 14427
rect 20496 14368 21128 14396
rect 20496 14356 20502 14368
rect 19429 14331 19487 14337
rect 19429 14297 19441 14331
rect 19475 14297 19487 14331
rect 19429 14291 19487 14297
rect 20165 14331 20223 14337
rect 20165 14297 20177 14331
rect 20211 14297 20223 14331
rect 21266 14328 21272 14340
rect 21227 14300 21272 14328
rect 20165 14291 20223 14297
rect 21266 14288 21272 14300
rect 21324 14288 21330 14340
rect 13679 14232 15424 14260
rect 16025 14263 16083 14269
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 16025 14229 16037 14263
rect 16071 14260 16083 14263
rect 16390 14260 16396 14272
rect 16071 14232 16396 14260
rect 16071 14229 16083 14232
rect 16025 14223 16083 14229
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 4154 14056 4160 14068
rect 4115 14028 4160 14056
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 7285 14059 7343 14065
rect 7285 14056 7297 14059
rect 6886 14028 7297 14056
rect 6886 13920 6914 14028
rect 7285 14025 7297 14028
rect 7331 14056 7343 14059
rect 8662 14056 8668 14068
rect 7331 14028 8668 14056
rect 7331 14025 7343 14028
rect 7285 14019 7343 14025
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 11054 14056 11060 14068
rect 10967 14028 11060 14056
rect 11054 14016 11060 14028
rect 11112 14056 11118 14068
rect 12802 14056 12808 14068
rect 11112 14028 12808 14056
rect 11112 14016 11118 14028
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 13998 14056 14004 14068
rect 13959 14028 14004 14056
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 15654 14056 15660 14068
rect 15615 14028 15660 14056
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 16577 14059 16635 14065
rect 16577 14025 16589 14059
rect 16623 14056 16635 14059
rect 20530 14056 20536 14068
rect 16623 14028 20536 14056
rect 16623 14025 16635 14028
rect 16577 14019 16635 14025
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 5460 13892 6914 13920
rect 5281 13855 5339 13861
rect 5281 13821 5293 13855
rect 5327 13852 5339 13855
rect 5460 13852 5488 13892
rect 12158 13880 12164 13932
rect 12216 13920 12222 13932
rect 14016 13920 14044 14016
rect 15013 13923 15071 13929
rect 15013 13920 15025 13923
rect 12216 13892 12756 13920
rect 14016 13892 15025 13920
rect 12216 13880 12222 13892
rect 5327 13824 5488 13852
rect 5537 13855 5595 13861
rect 5327 13821 5339 13824
rect 5281 13815 5339 13821
rect 5537 13821 5549 13855
rect 5583 13852 5595 13855
rect 7466 13852 7472 13864
rect 5583 13824 7472 13852
rect 5583 13821 5595 13824
rect 5537 13815 5595 13821
rect 7466 13812 7472 13824
rect 7524 13852 7530 13864
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 7524 13824 8677 13852
rect 7524 13812 7530 13824
rect 8220 13796 8248 13824
rect 8665 13821 8677 13824
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 12345 13855 12403 13861
rect 12345 13821 12357 13855
rect 12391 13852 12403 13855
rect 12621 13855 12679 13861
rect 12391 13824 12572 13852
rect 12391 13821 12403 13824
rect 12345 13815 12403 13821
rect 8202 13744 8208 13796
rect 8260 13744 8266 13796
rect 8478 13793 8484 13796
rect 8420 13787 8484 13793
rect 8420 13784 8432 13787
rect 8391 13756 8432 13784
rect 8420 13753 8432 13756
rect 8466 13753 8484 13787
rect 8420 13747 8484 13753
rect 8478 13744 8484 13747
rect 8536 13784 8542 13796
rect 9582 13784 9588 13796
rect 8536 13756 9588 13784
rect 8536 13744 8542 13756
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 12544 13716 12572 13824
rect 12621 13821 12633 13855
rect 12667 13821 12679 13855
rect 12728 13852 12756 13892
rect 15013 13889 15025 13892
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 17313 13923 17371 13929
rect 17313 13920 17325 13923
rect 17184 13892 17325 13920
rect 17184 13880 17190 13892
rect 17313 13889 17325 13892
rect 17359 13889 17371 13923
rect 21358 13920 21364 13932
rect 21319 13892 21364 13920
rect 17313 13883 17371 13889
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 12877 13855 12935 13861
rect 12877 13852 12889 13855
rect 12728 13824 12889 13852
rect 12621 13815 12679 13821
rect 12877 13821 12889 13824
rect 12923 13821 12935 13855
rect 14734 13852 14740 13864
rect 12877 13815 12935 13821
rect 13004 13824 14740 13852
rect 12636 13784 12664 13815
rect 13004 13784 13032 13824
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 16390 13852 16396 13864
rect 16351 13824 16396 13852
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 17580 13855 17638 13861
rect 17580 13821 17592 13855
rect 17626 13852 17638 13855
rect 18046 13852 18052 13864
rect 17626 13824 18052 13852
rect 17626 13821 17638 13824
rect 17580 13815 17638 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18874 13812 18880 13864
rect 18932 13852 18938 13864
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 18932 13824 19625 13852
rect 18932 13812 18938 13824
rect 19613 13821 19625 13824
rect 19659 13821 19671 13855
rect 19613 13815 19671 13821
rect 20349 13855 20407 13861
rect 20349 13821 20361 13855
rect 20395 13852 20407 13855
rect 20530 13852 20536 13864
rect 20395 13824 20536 13852
rect 20395 13821 20407 13824
rect 20349 13815 20407 13821
rect 20530 13812 20536 13824
rect 20588 13852 20594 13864
rect 20809 13855 20867 13861
rect 20809 13852 20821 13855
rect 20588 13824 20821 13852
rect 20588 13812 20594 13824
rect 20809 13821 20821 13824
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 12636 13756 13032 13784
rect 18598 13744 18604 13796
rect 18656 13784 18662 13796
rect 18969 13787 19027 13793
rect 18969 13784 18981 13787
rect 18656 13756 18981 13784
rect 18656 13744 18662 13756
rect 18969 13753 18981 13756
rect 19015 13753 19027 13787
rect 21174 13784 21180 13796
rect 21135 13756 21180 13784
rect 18969 13747 19027 13753
rect 21174 13744 21180 13756
rect 21232 13744 21238 13796
rect 13170 13716 13176 13728
rect 12544 13688 13176 13716
rect 13170 13676 13176 13688
rect 13228 13676 13234 13728
rect 15194 13716 15200 13728
rect 15155 13688 15200 13716
rect 15194 13676 15200 13688
rect 15252 13676 15258 13728
rect 15289 13719 15347 13725
rect 15289 13685 15301 13719
rect 15335 13716 15347 13719
rect 15933 13719 15991 13725
rect 15933 13716 15945 13719
rect 15335 13688 15945 13716
rect 15335 13685 15347 13688
rect 15289 13679 15347 13685
rect 15933 13685 15945 13688
rect 15979 13685 15991 13719
rect 18690 13716 18696 13728
rect 18651 13688 18696 13716
rect 15933 13679 15991 13685
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 20622 13716 20628 13728
rect 20583 13688 20628 13716
rect 20622 13676 20628 13688
rect 20680 13676 20686 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 6641 13515 6699 13521
rect 6641 13481 6653 13515
rect 6687 13512 6699 13515
rect 7190 13512 7196 13524
rect 6687 13484 7196 13512
rect 6687 13481 6699 13484
rect 6641 13475 6699 13481
rect 7190 13472 7196 13484
rect 7248 13472 7254 13524
rect 8849 13515 8907 13521
rect 8849 13481 8861 13515
rect 8895 13512 8907 13515
rect 9030 13512 9036 13524
rect 8895 13484 9036 13512
rect 8895 13481 8907 13484
rect 8849 13475 8907 13481
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 9309 13515 9367 13521
rect 9309 13481 9321 13515
rect 9355 13512 9367 13515
rect 9490 13512 9496 13524
rect 9355 13484 9496 13512
rect 9355 13481 9367 13484
rect 9309 13475 9367 13481
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 12526 13512 12532 13524
rect 12487 13484 12532 13512
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 12989 13515 13047 13521
rect 12989 13512 13001 13515
rect 12768 13484 13001 13512
rect 12768 13472 12774 13484
rect 12989 13481 13001 13484
rect 13035 13481 13047 13515
rect 12989 13475 13047 13481
rect 13449 13515 13507 13521
rect 13449 13481 13461 13515
rect 13495 13512 13507 13515
rect 14550 13512 14556 13524
rect 13495 13484 14556 13512
rect 13495 13481 13507 13484
rect 13449 13475 13507 13481
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15746 13512 15752 13524
rect 15252 13484 15752 13512
rect 15252 13472 15258 13484
rect 15746 13472 15752 13484
rect 15804 13512 15810 13524
rect 15841 13515 15899 13521
rect 15841 13512 15853 13515
rect 15804 13484 15853 13512
rect 15804 13472 15810 13484
rect 15841 13481 15853 13484
rect 15887 13512 15899 13515
rect 16482 13512 16488 13524
rect 15887 13484 16488 13512
rect 15887 13481 15899 13484
rect 15841 13475 15899 13481
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 18874 13512 18880 13524
rect 18835 13484 18880 13512
rect 18874 13472 18880 13484
rect 18932 13512 18938 13524
rect 19150 13512 19156 13524
rect 18932 13484 19156 13512
rect 18932 13472 18938 13484
rect 19150 13472 19156 13484
rect 19208 13472 19214 13524
rect 19334 13512 19340 13524
rect 19295 13484 19340 13512
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 20346 13512 20352 13524
rect 20307 13484 20352 13512
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 7776 13447 7834 13453
rect 7776 13413 7788 13447
rect 7822 13444 7834 13447
rect 18690 13444 18696 13456
rect 7822 13416 18696 13444
rect 7822 13413 7834 13416
rect 7776 13407 7834 13413
rect 18690 13404 18696 13416
rect 18748 13404 18754 13456
rect 21358 13444 21364 13456
rect 21319 13416 21364 13444
rect 21358 13404 21364 13416
rect 21416 13404 21422 13456
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13376 8999 13379
rect 9766 13376 9772 13388
rect 8987 13348 9772 13376
rect 8987 13345 8999 13348
rect 8941 13339 8999 13345
rect 9766 13336 9772 13348
rect 9824 13336 9830 13388
rect 10709 13379 10767 13385
rect 10709 13345 10721 13379
rect 10755 13376 10767 13379
rect 12250 13376 12256 13388
rect 10755 13348 12256 13376
rect 10755 13345 10767 13348
rect 10709 13339 10767 13345
rect 12250 13336 12256 13348
rect 12308 13336 12314 13388
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 12492 13348 12633 13376
rect 12492 13336 12498 13348
rect 12621 13345 12633 13348
rect 12667 13345 12679 13379
rect 12621 13339 12679 13345
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13308 8079 13311
rect 8202 13308 8208 13320
rect 8067 13280 8208 13308
rect 8067 13277 8079 13280
rect 8021 13271 8079 13277
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 8662 13308 8668 13320
rect 8623 13280 8668 13308
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 10965 13311 11023 13317
rect 10965 13277 10977 13311
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 8220 13240 8248 13268
rect 8220 13212 10088 13240
rect 9582 13172 9588 13184
rect 9543 13144 9588 13172
rect 9582 13132 9588 13144
rect 9640 13132 9646 13184
rect 10060 13172 10088 13212
rect 10980 13172 11008 13271
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 12216 13280 12357 13308
rect 12216 13268 12222 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 10060 13144 11008 13172
rect 12636 13172 12664 13339
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 13265 13379 13323 13385
rect 13265 13376 13277 13379
rect 12860 13348 13277 13376
rect 12860 13336 12866 13348
rect 13265 13345 13277 13348
rect 13311 13345 13323 13379
rect 13265 13339 13323 13345
rect 18969 13379 19027 13385
rect 18969 13345 18981 13379
rect 19015 13376 19027 13379
rect 19613 13379 19671 13385
rect 19613 13376 19625 13379
rect 19015 13348 19625 13376
rect 19015 13345 19027 13348
rect 18969 13339 19027 13345
rect 19613 13345 19625 13348
rect 19659 13345 19671 13379
rect 19613 13339 19671 13345
rect 20165 13379 20223 13385
rect 20165 13345 20177 13379
rect 20211 13376 20223 13379
rect 20622 13376 20628 13388
rect 20211 13348 20628 13376
rect 20211 13345 20223 13348
rect 20165 13339 20223 13345
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 20809 13379 20867 13385
rect 20809 13345 20821 13379
rect 20855 13345 20867 13379
rect 20809 13339 20867 13345
rect 12710 13268 12716 13320
rect 12768 13308 12774 13320
rect 13630 13308 13636 13320
rect 12768 13280 13636 13308
rect 12768 13268 12774 13280
rect 13630 13268 13636 13280
rect 13688 13308 13694 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13688 13280 14105 13308
rect 13688 13268 13694 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 18046 13268 18052 13320
rect 18104 13308 18110 13320
rect 18693 13311 18751 13317
rect 18693 13308 18705 13311
rect 18104 13280 18705 13308
rect 18104 13268 18110 13280
rect 18693 13277 18705 13280
rect 18739 13277 18751 13311
rect 18693 13271 18751 13277
rect 20346 13268 20352 13320
rect 20404 13308 20410 13320
rect 20824 13308 20852 13339
rect 20898 13336 20904 13388
rect 20956 13376 20962 13388
rect 21177 13379 21235 13385
rect 21177 13376 21189 13379
rect 20956 13348 21189 13376
rect 20956 13336 20962 13348
rect 21177 13345 21189 13348
rect 21223 13345 21235 13379
rect 21177 13339 21235 13345
rect 20404 13280 20852 13308
rect 20404 13268 20410 13280
rect 20070 13200 20076 13252
rect 20128 13240 20134 13252
rect 20625 13243 20683 13249
rect 20625 13240 20637 13243
rect 20128 13212 20637 13240
rect 20128 13200 20134 13212
rect 20625 13209 20637 13212
rect 20671 13209 20683 13243
rect 20625 13203 20683 13209
rect 13538 13172 13544 13184
rect 12636 13144 13544 13172
rect 13538 13132 13544 13144
rect 13596 13172 13602 13184
rect 13725 13175 13783 13181
rect 13725 13172 13737 13175
rect 13596 13144 13737 13172
rect 13596 13132 13602 13144
rect 13725 13141 13737 13144
rect 13771 13141 13783 13175
rect 13725 13135 13783 13141
rect 16298 13132 16304 13184
rect 16356 13172 16362 13184
rect 17037 13175 17095 13181
rect 17037 13172 17049 13175
rect 16356 13144 17049 13172
rect 16356 13132 16362 13144
rect 17037 13141 17049 13144
rect 17083 13172 17095 13175
rect 18598 13172 18604 13184
rect 17083 13144 18604 13172
rect 17083 13141 17095 13144
rect 17037 13135 17095 13141
rect 18598 13132 18604 13144
rect 18656 13132 18662 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 9766 12968 9772 12980
rect 9727 12940 9772 12968
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 12158 12968 12164 12980
rect 12119 12940 12164 12968
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 13817 12971 13875 12977
rect 13817 12937 13829 12971
rect 13863 12968 13875 12971
rect 19981 12971 20039 12977
rect 13863 12940 19932 12968
rect 13863 12937 13875 12940
rect 13817 12931 13875 12937
rect 15286 12860 15292 12912
rect 15344 12900 15350 12912
rect 15344 12872 17080 12900
rect 15344 12860 15350 12872
rect 9582 12792 9588 12844
rect 9640 12832 9646 12844
rect 10321 12835 10379 12841
rect 10321 12832 10333 12835
rect 9640 12804 10333 12832
rect 9640 12792 9646 12804
rect 10321 12801 10333 12804
rect 10367 12801 10379 12835
rect 10321 12795 10379 12801
rect 16390 12792 16396 12844
rect 16448 12832 16454 12844
rect 17052 12841 17080 12872
rect 16577 12835 16635 12841
rect 16448 12804 16493 12832
rect 16448 12792 16454 12804
rect 16577 12801 16589 12835
rect 16623 12801 16635 12835
rect 16577 12795 16635 12801
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12764 10839 12767
rect 12434 12764 12440 12776
rect 10827 12736 12440 12764
rect 10827 12733 10839 12736
rect 10781 12727 10839 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 13906 12764 13912 12776
rect 13679 12736 13912 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 13906 12724 13912 12736
rect 13964 12724 13970 12776
rect 16298 12764 16304 12776
rect 16259 12736 16304 12764
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 16592 12764 16620 12795
rect 17126 12792 17132 12844
rect 17184 12832 17190 12844
rect 17221 12835 17279 12841
rect 17221 12832 17233 12835
rect 17184 12804 17233 12832
rect 17184 12792 17190 12804
rect 17221 12801 17233 12804
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17494 12832 17500 12844
rect 17368 12804 17500 12832
rect 17368 12792 17374 12804
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 19904 12832 19932 12940
rect 19981 12937 19993 12971
rect 20027 12968 20039 12971
rect 20346 12968 20352 12980
rect 20027 12940 20352 12968
rect 20027 12937 20039 12940
rect 19981 12931 20039 12937
rect 20346 12928 20352 12940
rect 20404 12928 20410 12980
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 21174 12968 21180 12980
rect 21135 12940 21180 12968
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 20438 12900 20444 12912
rect 20399 12872 20444 12900
rect 20438 12860 20444 12872
rect 20496 12860 20502 12912
rect 19904 12804 21404 12832
rect 17678 12764 17684 12776
rect 16592 12736 17684 12764
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 19245 12767 19303 12773
rect 19245 12733 19257 12767
rect 19291 12764 19303 12767
rect 19794 12764 19800 12776
rect 19291 12736 19800 12764
rect 19291 12733 19303 12736
rect 19245 12727 19303 12733
rect 19794 12724 19800 12736
rect 19852 12724 19858 12776
rect 20257 12767 20315 12773
rect 20257 12733 20269 12767
rect 20303 12733 20315 12767
rect 20257 12727 20315 12733
rect 11054 12705 11060 12708
rect 10137 12699 10195 12705
rect 10137 12665 10149 12699
rect 10183 12696 10195 12699
rect 10183 12668 11008 12696
rect 10183 12665 10195 12668
rect 10137 12659 10195 12665
rect 10229 12631 10287 12637
rect 10229 12597 10241 12631
rect 10275 12628 10287 12631
rect 10686 12628 10692 12640
rect 10275 12600 10692 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 10686 12588 10692 12600
rect 10744 12588 10750 12640
rect 10980 12628 11008 12668
rect 11048 12659 11060 12705
rect 11112 12696 11118 12708
rect 11112 12668 11148 12696
rect 11054 12656 11060 12659
rect 11112 12656 11118 12668
rect 15194 12656 15200 12708
rect 15252 12696 15258 12708
rect 15252 12668 16528 12696
rect 15252 12656 15258 12668
rect 11146 12628 11152 12640
rect 10980 12600 11152 12628
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 15930 12628 15936 12640
rect 15891 12600 15936 12628
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16500 12628 16528 12668
rect 16574 12656 16580 12708
rect 16632 12696 16638 12708
rect 17126 12696 17132 12708
rect 16632 12668 17132 12696
rect 16632 12656 16638 12668
rect 17126 12656 17132 12668
rect 17184 12656 17190 12708
rect 20272 12696 20300 12727
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 21376 12773 21404 12804
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 20496 12736 20729 12764
rect 20496 12724 20502 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12733 21419 12767
rect 21361 12727 21419 12733
rect 17236 12668 20300 12696
rect 17236 12628 17264 12668
rect 16500 12600 17264 12628
rect 17313 12631 17371 12637
rect 17313 12597 17325 12631
rect 17359 12628 17371 12631
rect 17494 12628 17500 12640
rect 17359 12600 17500 12628
rect 17359 12597 17371 12600
rect 17313 12591 17371 12597
rect 17494 12588 17500 12600
rect 17552 12588 17558 12640
rect 17681 12631 17739 12637
rect 17681 12597 17693 12631
rect 17727 12628 17739 12631
rect 18966 12628 18972 12640
rect 17727 12600 18972 12628
rect 17727 12597 17739 12600
rect 17681 12591 17739 12597
rect 18966 12588 18972 12600
rect 19024 12588 19030 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 10686 12424 10692 12436
rect 10647 12396 10692 12424
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 11057 12427 11115 12433
rect 11057 12393 11069 12427
rect 11103 12424 11115 12427
rect 11146 12424 11152 12436
rect 11103 12396 11152 12424
rect 11103 12393 11115 12396
rect 11057 12387 11115 12393
rect 11146 12384 11152 12396
rect 11204 12384 11210 12436
rect 12069 12427 12127 12433
rect 12069 12393 12081 12427
rect 12115 12424 12127 12427
rect 15194 12424 15200 12436
rect 12115 12396 15200 12424
rect 12115 12393 12127 12396
rect 12069 12387 12127 12393
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 15930 12384 15936 12436
rect 15988 12424 15994 12436
rect 16117 12427 16175 12433
rect 16117 12424 16129 12427
rect 15988 12396 16129 12424
rect 15988 12384 15994 12396
rect 16117 12393 16129 12396
rect 16163 12393 16175 12427
rect 16574 12424 16580 12436
rect 16535 12396 16580 12424
rect 16117 12387 16175 12393
rect 16574 12384 16580 12396
rect 16632 12384 16638 12436
rect 17129 12427 17187 12433
rect 17129 12393 17141 12427
rect 17175 12393 17187 12427
rect 17129 12387 17187 12393
rect 19521 12427 19579 12433
rect 19521 12393 19533 12427
rect 19567 12393 19579 12427
rect 19521 12387 19579 12393
rect 14216 12359 14274 12365
rect 14216 12325 14228 12359
rect 14262 12356 14274 12359
rect 15286 12356 15292 12368
rect 14262 12328 15292 12356
rect 14262 12325 14274 12328
rect 14216 12319 14274 12325
rect 15286 12316 15292 12328
rect 15344 12316 15350 12368
rect 16209 12359 16267 12365
rect 16209 12325 16221 12359
rect 16255 12356 16267 12359
rect 17144 12356 17172 12387
rect 16255 12328 17172 12356
rect 16255 12325 16267 12328
rect 16209 12319 16267 12325
rect 18966 12316 18972 12368
rect 19024 12356 19030 12368
rect 19536 12356 19564 12387
rect 20162 12384 20168 12436
rect 20220 12424 20226 12436
rect 20349 12427 20407 12433
rect 20349 12424 20361 12427
rect 20220 12396 20361 12424
rect 20220 12384 20226 12396
rect 20349 12393 20361 12396
rect 20395 12393 20407 12427
rect 20349 12387 20407 12393
rect 20622 12384 20628 12436
rect 20680 12424 20686 12436
rect 20809 12427 20867 12433
rect 20809 12424 20821 12427
rect 20680 12396 20821 12424
rect 20680 12384 20686 12396
rect 20809 12393 20821 12396
rect 20855 12393 20867 12427
rect 20809 12387 20867 12393
rect 19024 12328 19472 12356
rect 19536 12328 20576 12356
rect 19024 12316 19030 12328
rect 8665 12291 8723 12297
rect 8665 12257 8677 12291
rect 8711 12288 8723 12291
rect 9306 12288 9312 12300
rect 8711 12260 9312 12288
rect 8711 12257 8723 12260
rect 8665 12251 8723 12257
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 11885 12291 11943 12297
rect 11885 12288 11897 12291
rect 11756 12260 11897 12288
rect 11756 12248 11762 12260
rect 11885 12257 11897 12260
rect 11931 12257 11943 12291
rect 11885 12251 11943 12257
rect 12434 12248 12440 12300
rect 12492 12288 12498 12300
rect 14461 12291 14519 12297
rect 14461 12288 14473 12291
rect 12492 12260 14473 12288
rect 12492 12248 12498 12260
rect 14461 12257 14473 12260
rect 14507 12257 14519 12291
rect 17497 12291 17555 12297
rect 17497 12288 17509 12291
rect 14461 12251 14519 12257
rect 17144 12260 17509 12288
rect 15930 12220 15936 12232
rect 15891 12192 15936 12220
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 8938 12112 8944 12164
rect 8996 12152 9002 12164
rect 8996 12124 13584 12152
rect 8996 12112 9002 12124
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8481 12087 8539 12093
rect 8481 12084 8493 12087
rect 8260 12056 8493 12084
rect 8260 12044 8266 12056
rect 8481 12053 8493 12056
rect 8527 12053 8539 12087
rect 13078 12084 13084 12096
rect 13039 12056 13084 12084
rect 8481 12047 8539 12053
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 13556 12084 13584 12124
rect 17144 12084 17172 12260
rect 17497 12257 17509 12260
rect 17543 12288 17555 12291
rect 19061 12291 19119 12297
rect 17543 12260 18644 12288
rect 17543 12257 17555 12260
rect 17497 12251 17555 12257
rect 17586 12220 17592 12232
rect 17547 12192 17592 12220
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 17678 12180 17684 12232
rect 17736 12220 17742 12232
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 17736 12192 17785 12220
rect 17736 12180 17742 12192
rect 17773 12189 17785 12192
rect 17819 12220 17831 12223
rect 17862 12220 17868 12232
rect 17819 12192 17868 12220
rect 17819 12189 17831 12192
rect 17773 12183 17831 12189
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 17604 12152 17632 12180
rect 18141 12155 18199 12161
rect 18141 12152 18153 12155
rect 17604 12124 18153 12152
rect 18141 12121 18153 12124
rect 18187 12121 18199 12155
rect 18141 12115 18199 12121
rect 18616 12093 18644 12260
rect 19061 12257 19073 12291
rect 19107 12288 19119 12291
rect 19242 12288 19248 12300
rect 19107 12260 19248 12288
rect 19107 12257 19119 12260
rect 19061 12251 19119 12257
rect 19242 12248 19248 12260
rect 19300 12288 19306 12300
rect 19337 12291 19395 12297
rect 19337 12288 19349 12291
rect 19300 12260 19349 12288
rect 19300 12248 19306 12260
rect 19337 12257 19349 12260
rect 19383 12257 19395 12291
rect 19444 12288 19472 12328
rect 20548 12297 20576 12328
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 19444 12260 19809 12288
rect 19337 12251 19395 12257
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 20533 12291 20591 12297
rect 20533 12257 20545 12291
rect 20579 12257 20591 12291
rect 20533 12251 20591 12257
rect 20993 12291 21051 12297
rect 20993 12257 21005 12291
rect 21039 12257 21051 12291
rect 20993 12251 21051 12257
rect 20070 12180 20076 12232
rect 20128 12220 20134 12232
rect 21008 12220 21036 12251
rect 20128 12192 21036 12220
rect 20128 12180 20134 12192
rect 19981 12155 20039 12161
rect 19981 12121 19993 12155
rect 20027 12152 20039 12155
rect 20438 12152 20444 12164
rect 20027 12124 20444 12152
rect 20027 12121 20039 12124
rect 19981 12115 20039 12121
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 13556 12056 17172 12084
rect 18601 12087 18659 12093
rect 18601 12053 18613 12087
rect 18647 12084 18659 12087
rect 19334 12084 19340 12096
rect 18647 12056 19340 12084
rect 18647 12053 18659 12056
rect 18601 12047 18659 12053
rect 19334 12044 19340 12056
rect 19392 12044 19398 12096
rect 19610 12044 19616 12096
rect 19668 12084 19674 12096
rect 20622 12084 20628 12096
rect 19668 12056 20628 12084
rect 19668 12044 19674 12056
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 21358 12084 21364 12096
rect 21319 12056 21364 12084
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 11698 11880 11704 11892
rect 11659 11852 11704 11880
rect 11698 11840 11704 11852
rect 11756 11840 11762 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13630 11880 13636 11892
rect 13412 11852 13636 11880
rect 13412 11840 13418 11852
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 14829 11883 14887 11889
rect 14829 11849 14841 11883
rect 14875 11880 14887 11883
rect 15286 11880 15292 11892
rect 14875 11852 15292 11880
rect 14875 11849 14887 11852
rect 14829 11843 14887 11849
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 17405 11883 17463 11889
rect 17405 11880 17417 11883
rect 17368 11852 17417 11880
rect 17368 11840 17374 11852
rect 17405 11849 17417 11852
rect 17451 11849 17463 11883
rect 17405 11843 17463 11849
rect 18782 11840 18788 11892
rect 18840 11880 18846 11892
rect 19061 11883 19119 11889
rect 19061 11880 19073 11883
rect 18840 11852 19073 11880
rect 18840 11840 18846 11852
rect 19061 11849 19073 11852
rect 19107 11849 19119 11883
rect 20070 11880 20076 11892
rect 20031 11852 20076 11880
rect 19061 11843 19119 11849
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 20254 11840 20260 11892
rect 20312 11880 20318 11892
rect 20809 11883 20867 11889
rect 20809 11880 20821 11883
rect 20312 11852 20821 11880
rect 20312 11840 20318 11852
rect 20809 11849 20821 11852
rect 20855 11849 20867 11883
rect 20809 11843 20867 11849
rect 10689 11815 10747 11821
rect 10689 11781 10701 11815
rect 10735 11781 10747 11815
rect 10689 11775 10747 11781
rect 20533 11815 20591 11821
rect 20533 11781 20545 11815
rect 20579 11781 20591 11815
rect 20533 11775 20591 11781
rect 10704 11744 10732 11775
rect 11054 11744 11060 11756
rect 10704 11716 11060 11744
rect 11054 11704 11060 11716
rect 11112 11704 11118 11756
rect 13078 11704 13084 11756
rect 13136 11744 13142 11756
rect 13630 11744 13636 11756
rect 13136 11716 13636 11744
rect 13136 11704 13142 11716
rect 13630 11704 13636 11716
rect 13688 11744 13694 11756
rect 13725 11747 13783 11753
rect 13725 11744 13737 11747
rect 13688 11716 13737 11744
rect 13688 11704 13694 11716
rect 13725 11713 13737 11716
rect 13771 11713 13783 11747
rect 17957 11747 18015 11753
rect 17957 11744 17969 11747
rect 13725 11707 13783 11713
rect 16132 11716 17969 11744
rect 2314 11636 2320 11688
rect 2372 11676 2378 11688
rect 2372 11648 2774 11676
rect 2372 11636 2378 11648
rect 2746 11540 2774 11648
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 8260 11648 9321 11676
rect 8260 11636 8266 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 15930 11676 15936 11688
rect 15988 11685 15994 11688
rect 15988 11679 16011 11685
rect 15863 11648 15936 11676
rect 9309 11639 9367 11645
rect 15930 11636 15936 11648
rect 15999 11676 16011 11679
rect 16132 11676 16160 11716
rect 17957 11713 17969 11716
rect 18003 11713 18015 11747
rect 17957 11707 18015 11713
rect 15999 11648 16160 11676
rect 16209 11679 16267 11685
rect 15999 11645 16011 11648
rect 15988 11639 16011 11645
rect 16209 11645 16221 11679
rect 16255 11645 16267 11679
rect 18690 11676 18696 11688
rect 16209 11639 16267 11645
rect 16316 11648 18696 11676
rect 15988 11636 15994 11639
rect 9214 11568 9220 11620
rect 9272 11608 9278 11620
rect 9554 11611 9612 11617
rect 9554 11608 9566 11611
rect 9272 11580 9566 11608
rect 9272 11568 9278 11580
rect 9554 11577 9566 11580
rect 9600 11577 9612 11611
rect 12897 11611 12955 11617
rect 12897 11608 12909 11611
rect 9554 11571 9612 11577
rect 9692 11580 12909 11608
rect 9692 11540 9720 11580
rect 12897 11577 12909 11580
rect 12943 11608 12955 11611
rect 13633 11611 13691 11617
rect 13633 11608 13645 11611
rect 12943 11580 13645 11608
rect 12943 11577 12955 11580
rect 12897 11571 12955 11577
rect 13633 11577 13645 11580
rect 13679 11577 13691 11611
rect 13633 11571 13691 11577
rect 13722 11568 13728 11620
rect 13780 11608 13786 11620
rect 16224 11608 16252 11639
rect 13780 11580 16252 11608
rect 13780 11568 13786 11580
rect 2746 11512 9720 11540
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 9824 11512 11253 11540
rect 9824 11500 9830 11512
rect 11241 11509 11253 11512
rect 11287 11509 11299 11543
rect 11241 11503 11299 11509
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 13170 11540 13176 11552
rect 11388 11512 11433 11540
rect 13131 11512 13176 11540
rect 11388 11500 11394 11512
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 13446 11500 13452 11552
rect 13504 11540 13510 11552
rect 13541 11543 13599 11549
rect 13541 11540 13553 11543
rect 13504 11512 13553 11540
rect 13504 11500 13510 11512
rect 13541 11509 13553 11512
rect 13587 11540 13599 11543
rect 14461 11543 14519 11549
rect 14461 11540 14473 11543
rect 13587 11512 14473 11540
rect 13587 11509 13599 11512
rect 13541 11503 13599 11509
rect 14461 11509 14473 11512
rect 14507 11540 14519 11543
rect 16316 11540 16344 11648
rect 18690 11636 18696 11648
rect 18748 11636 18754 11688
rect 19058 11636 19064 11688
rect 19116 11676 19122 11688
rect 19245 11679 19303 11685
rect 19245 11676 19257 11679
rect 19116 11648 19257 11676
rect 19116 11636 19122 11648
rect 19245 11645 19257 11648
rect 19291 11645 19303 11679
rect 19245 11639 19303 11645
rect 19889 11679 19947 11685
rect 19889 11645 19901 11679
rect 19935 11645 19947 11679
rect 19889 11639 19947 11645
rect 20349 11679 20407 11685
rect 20349 11645 20361 11679
rect 20395 11645 20407 11679
rect 20548 11676 20576 11775
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20548 11648 21005 11676
rect 20349 11639 20407 11645
rect 20993 11645 21005 11648
rect 21039 11645 21051 11679
rect 20993 11639 21051 11645
rect 21085 11679 21143 11685
rect 21085 11645 21097 11679
rect 21131 11676 21143 11679
rect 21358 11676 21364 11688
rect 21131 11648 21364 11676
rect 21131 11645 21143 11648
rect 21085 11639 21143 11645
rect 17773 11611 17831 11617
rect 17773 11577 17785 11611
rect 17819 11608 17831 11611
rect 18417 11611 18475 11617
rect 18417 11608 18429 11611
rect 17819 11580 18429 11608
rect 17819 11577 17831 11580
rect 17773 11571 17831 11577
rect 18417 11577 18429 11580
rect 18463 11577 18475 11611
rect 18417 11571 18475 11577
rect 14507 11512 16344 11540
rect 17865 11543 17923 11549
rect 14507 11509 14519 11512
rect 14461 11503 14519 11509
rect 17865 11509 17877 11543
rect 17911 11540 17923 11543
rect 18046 11540 18052 11552
rect 17911 11512 18052 11540
rect 17911 11509 17923 11512
rect 17865 11503 17923 11509
rect 18046 11500 18052 11512
rect 18104 11500 18110 11552
rect 19904 11540 19932 11639
rect 20364 11608 20392 11639
rect 21358 11636 21364 11648
rect 21416 11636 21422 11688
rect 20364 11580 21404 11608
rect 21376 11552 21404 11580
rect 21085 11543 21143 11549
rect 21085 11540 21097 11543
rect 19904 11512 21097 11540
rect 21085 11509 21097 11512
rect 21131 11509 21143 11543
rect 21358 11540 21364 11552
rect 21319 11512 21364 11540
rect 21085 11503 21143 11509
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 8757 11339 8815 11345
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 9309 11339 9367 11345
rect 9309 11336 9321 11339
rect 8803 11308 9321 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 9309 11305 9321 11308
rect 9355 11305 9367 11339
rect 9766 11336 9772 11348
rect 9727 11308 9772 11336
rect 9309 11299 9367 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 11149 11339 11207 11345
rect 11149 11305 11161 11339
rect 11195 11336 11207 11339
rect 11330 11336 11336 11348
rect 11195 11308 11336 11336
rect 11195 11305 11207 11308
rect 11149 11299 11207 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 13906 11336 13912 11348
rect 13867 11308 13912 11336
rect 13906 11296 13912 11308
rect 13964 11296 13970 11348
rect 18046 11336 18052 11348
rect 18007 11308 18052 11336
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 19058 11336 19064 11348
rect 19019 11308 19064 11336
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 20073 11339 20131 11345
rect 20073 11305 20085 11339
rect 20119 11305 20131 11339
rect 20073 11299 20131 11305
rect 8297 11271 8355 11277
rect 8297 11237 8309 11271
rect 8343 11268 8355 11271
rect 8846 11268 8852 11280
rect 8343 11240 8852 11268
rect 8343 11237 8355 11240
rect 8297 11231 8355 11237
rect 8846 11228 8852 11240
rect 8904 11228 8910 11280
rect 9674 11268 9680 11280
rect 9232 11240 9680 11268
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 9232 11200 9260 11240
rect 9674 11228 9680 11240
rect 9732 11268 9738 11280
rect 10137 11271 10195 11277
rect 10137 11268 10149 11271
rect 9732 11240 10149 11268
rect 9732 11228 9738 11240
rect 10137 11237 10149 11240
rect 10183 11268 10195 11271
rect 16298 11268 16304 11280
rect 10183 11240 16304 11268
rect 10183 11237 10195 11240
rect 10137 11231 10195 11237
rect 16298 11228 16304 11240
rect 16356 11228 16362 11280
rect 18509 11271 18567 11277
rect 18509 11237 18521 11271
rect 18555 11268 18567 11271
rect 18966 11268 18972 11280
rect 18555 11240 18972 11268
rect 18555 11237 18567 11240
rect 18509 11231 18567 11237
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 20088 11268 20116 11299
rect 20622 11296 20628 11348
rect 20680 11336 20686 11348
rect 20809 11339 20867 11345
rect 20809 11336 20821 11339
rect 20680 11308 20821 11336
rect 20680 11296 20686 11308
rect 20809 11305 20821 11308
rect 20855 11305 20867 11339
rect 20809 11299 20867 11305
rect 20088 11240 21036 11268
rect 9398 11200 9404 11212
rect 8435 11172 9260 11200
rect 9359 11172 9404 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 10778 11200 10784 11212
rect 10739 11172 10784 11200
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 13541 11203 13599 11209
rect 13541 11169 13553 11203
rect 13587 11200 13599 11203
rect 14366 11200 14372 11212
rect 13587 11172 14372 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 14550 11200 14556 11212
rect 14511 11172 14556 11200
rect 14550 11160 14556 11172
rect 14608 11160 14614 11212
rect 16482 11160 16488 11212
rect 16540 11200 16546 11212
rect 17773 11203 17831 11209
rect 17773 11200 17785 11203
rect 16540 11172 17785 11200
rect 16540 11160 16546 11172
rect 17773 11169 17785 11172
rect 17819 11200 17831 11203
rect 18417 11203 18475 11209
rect 18417 11200 18429 11203
rect 17819 11172 18429 11200
rect 17819 11169 17831 11172
rect 17773 11163 17831 11169
rect 18417 11169 18429 11172
rect 18463 11200 18475 11203
rect 18782 11200 18788 11212
rect 18463 11172 18788 11200
rect 18463 11169 18475 11172
rect 18417 11163 18475 11169
rect 18782 11160 18788 11172
rect 18840 11200 18846 11212
rect 19150 11200 19156 11212
rect 18840 11172 19156 11200
rect 18840 11160 18846 11172
rect 19150 11160 19156 11172
rect 19208 11160 19214 11212
rect 19245 11203 19303 11209
rect 19245 11169 19257 11203
rect 19291 11200 19303 11203
rect 19794 11200 19800 11212
rect 19291 11172 19800 11200
rect 19291 11169 19303 11172
rect 19245 11163 19303 11169
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 19886 11160 19892 11212
rect 19944 11200 19950 11212
rect 21008 11209 21036 11240
rect 20533 11203 20591 11209
rect 19944 11172 19989 11200
rect 19944 11160 19950 11172
rect 20533 11169 20545 11203
rect 20579 11169 20591 11203
rect 20533 11163 20591 11169
rect 20993 11203 21051 11209
rect 20993 11169 21005 11203
rect 21039 11169 21051 11203
rect 20993 11163 21051 11169
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 8294 11132 8300 11144
rect 8251 11104 8300 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 9214 11132 9220 11144
rect 9175 11104 9220 11132
rect 9214 11092 9220 11104
rect 9272 11132 9278 11144
rect 10505 11135 10563 11141
rect 10505 11132 10517 11135
rect 9272 11104 10517 11132
rect 9272 11092 9278 11104
rect 10505 11101 10517 11104
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11132 10747 11135
rect 11054 11132 11060 11144
rect 10735 11104 11060 11132
rect 10735 11101 10747 11104
rect 10689 11095 10747 11101
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 13265 11135 13323 11141
rect 13265 11132 13277 11135
rect 11848 11104 13277 11132
rect 11848 11092 11854 11104
rect 13265 11101 13277 11104
rect 13311 11101 13323 11135
rect 13446 11132 13452 11144
rect 13407 11104 13452 11132
rect 13265 11095 13323 11101
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 18601 11135 18659 11141
rect 18601 11101 18613 11135
rect 18647 11101 18659 11135
rect 18601 11095 18659 11101
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11132 19671 11135
rect 19904 11132 19932 11160
rect 19659 11104 19932 11132
rect 20548 11132 20576 11163
rect 20548 11104 21404 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 14752 11036 16528 11064
rect 13722 10956 13728 11008
rect 13780 10996 13786 11008
rect 14752 11005 14780 11036
rect 14737 10999 14795 11005
rect 14737 10996 14749 10999
rect 13780 10968 14749 10996
rect 13780 10956 13786 10968
rect 14737 10965 14749 10968
rect 14783 10965 14795 10999
rect 16500 10996 16528 11036
rect 17862 11024 17868 11076
rect 17920 11064 17926 11076
rect 18616 11064 18644 11095
rect 21376 11076 21404 11104
rect 20346 11064 20352 11076
rect 17920 11036 18644 11064
rect 20307 11036 20352 11064
rect 17920 11024 17926 11036
rect 20346 11024 20352 11036
rect 20404 11024 20410 11076
rect 21358 11064 21364 11076
rect 21319 11036 21364 11064
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 18046 10996 18052 11008
rect 16500 10968 18052 10996
rect 14737 10959 14795 10965
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 8757 10795 8815 10801
rect 8757 10761 8769 10795
rect 8803 10792 8815 10795
rect 9398 10792 9404 10804
rect 8803 10764 9404 10792
rect 8803 10761 8815 10764
rect 8757 10755 8815 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 11054 10792 11060 10804
rect 11015 10764 11060 10792
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 11931 10764 12572 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 12544 10733 12572 10764
rect 13446 10752 13452 10804
rect 13504 10792 13510 10804
rect 13725 10795 13783 10801
rect 13725 10792 13737 10795
rect 13504 10764 13737 10792
rect 13504 10752 13510 10764
rect 13725 10761 13737 10764
rect 13771 10761 13783 10795
rect 13725 10755 13783 10761
rect 15930 10752 15936 10804
rect 15988 10792 15994 10804
rect 16117 10795 16175 10801
rect 16117 10792 16129 10795
rect 15988 10764 16129 10792
rect 15988 10752 15994 10764
rect 16117 10761 16129 10764
rect 16163 10761 16175 10795
rect 16117 10755 16175 10761
rect 16206 10752 16212 10804
rect 16264 10792 16270 10804
rect 19794 10792 19800 10804
rect 16264 10764 18552 10792
rect 19755 10764 19800 10792
rect 16264 10752 16270 10764
rect 10045 10727 10103 10733
rect 10045 10693 10057 10727
rect 10091 10724 10103 10727
rect 12529 10727 12587 10733
rect 10091 10696 12434 10724
rect 10091 10693 10103 10696
rect 10045 10687 10103 10693
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10656 8263 10659
rect 8294 10656 8300 10668
rect 8251 10628 8300 10656
rect 8251 10625 8263 10628
rect 8205 10619 8263 10625
rect 8294 10616 8300 10628
rect 8352 10656 8358 10668
rect 10778 10656 10784 10668
rect 8352 10628 9628 10656
rect 10739 10628 10784 10656
rect 8352 10616 8358 10628
rect 9600 10600 9628 10628
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 11609 10659 11667 10665
rect 11609 10625 11621 10659
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8938 10588 8944 10600
rect 8435 10560 8944 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 9582 10548 9588 10600
rect 9640 10588 9646 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9640 10560 9873 10588
rect 9640 10548 9646 10560
rect 9861 10557 9873 10560
rect 9907 10588 9919 10591
rect 11624 10588 11652 10619
rect 9907 10560 11652 10588
rect 12406 10588 12434 10696
rect 12529 10693 12541 10727
rect 12575 10724 12587 10727
rect 16482 10724 16488 10736
rect 12575 10696 16488 10724
rect 12575 10693 12587 10696
rect 12529 10687 12587 10693
rect 16482 10684 16488 10696
rect 16540 10684 16546 10736
rect 17681 10727 17739 10733
rect 17681 10693 17693 10727
rect 17727 10724 17739 10727
rect 17865 10727 17923 10733
rect 17865 10724 17877 10727
rect 17727 10696 17877 10724
rect 17727 10693 17739 10696
rect 17681 10687 17739 10693
rect 17865 10693 17877 10696
rect 17911 10693 17923 10727
rect 18524 10724 18552 10764
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 20809 10727 20867 10733
rect 20809 10724 20821 10727
rect 18524 10696 20821 10724
rect 17865 10687 17923 10693
rect 20809 10693 20821 10696
rect 20855 10693 20867 10727
rect 20809 10687 20867 10693
rect 12894 10616 12900 10668
rect 12952 10656 12958 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 12952 10628 13093 10656
rect 12952 10616 12958 10628
rect 13081 10625 13093 10628
rect 13127 10625 13139 10659
rect 13081 10619 13139 10625
rect 13170 10616 13176 10668
rect 13228 10656 13234 10668
rect 13265 10659 13323 10665
rect 13265 10656 13277 10659
rect 13228 10628 13277 10656
rect 13228 10616 13234 10628
rect 13265 10625 13277 10628
rect 13311 10625 13323 10659
rect 18046 10656 18052 10668
rect 13265 10619 13323 10625
rect 17696 10628 18052 10656
rect 16666 10588 16672 10600
rect 12406 10560 16672 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 17497 10591 17555 10597
rect 17497 10557 17509 10591
rect 17543 10588 17555 10591
rect 17696 10588 17724 10628
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 20070 10616 20076 10668
rect 20128 10656 20134 10668
rect 20349 10659 20407 10665
rect 20349 10656 20361 10659
rect 20128 10628 20361 10656
rect 20128 10616 20134 10628
rect 20349 10625 20361 10628
rect 20395 10625 20407 10659
rect 20349 10619 20407 10625
rect 17543 10560 17724 10588
rect 17543 10557 17555 10560
rect 17497 10551 17555 10557
rect 17862 10548 17868 10600
rect 17920 10588 17926 10600
rect 18325 10591 18383 10597
rect 18325 10588 18337 10591
rect 17920 10560 18337 10588
rect 17920 10548 17926 10560
rect 18325 10557 18337 10560
rect 18371 10557 18383 10591
rect 18325 10551 18383 10557
rect 20530 10548 20536 10600
rect 20588 10588 20594 10600
rect 20993 10591 21051 10597
rect 20993 10588 21005 10591
rect 20588 10560 21005 10588
rect 20588 10548 20594 10560
rect 20993 10557 21005 10560
rect 21039 10557 21051 10591
rect 20993 10551 21051 10557
rect 7650 10480 7656 10532
rect 7708 10520 7714 10532
rect 8297 10523 8355 10529
rect 8297 10520 8309 10523
rect 7708 10492 8309 10520
rect 7708 10480 7714 10492
rect 8297 10489 8309 10492
rect 8343 10520 8355 10523
rect 10045 10523 10103 10529
rect 10045 10520 10057 10523
rect 8343 10492 10057 10520
rect 8343 10489 8355 10492
rect 8297 10483 8355 10489
rect 10045 10489 10057 10492
rect 10091 10520 10103 10523
rect 10137 10523 10195 10529
rect 10137 10520 10149 10523
rect 10091 10492 10149 10520
rect 10091 10489 10103 10492
rect 10045 10483 10103 10489
rect 10137 10489 10149 10492
rect 10183 10489 10195 10523
rect 10137 10483 10195 10489
rect 10686 10480 10692 10532
rect 10744 10520 10750 10532
rect 11425 10523 11483 10529
rect 11425 10520 11437 10523
rect 10744 10492 11437 10520
rect 10744 10480 10750 10492
rect 11425 10489 11437 10492
rect 11471 10520 11483 10523
rect 11885 10523 11943 10529
rect 11885 10520 11897 10523
rect 11471 10492 11897 10520
rect 11471 10489 11483 10492
rect 11425 10483 11483 10489
rect 11885 10489 11897 10492
rect 11931 10489 11943 10523
rect 14642 10520 14648 10532
rect 11885 10483 11943 10489
rect 12406 10492 14648 10520
rect 9398 10452 9404 10464
rect 9359 10424 9404 10452
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 11517 10455 11575 10461
rect 11517 10421 11529 10455
rect 11563 10452 11575 10455
rect 12069 10455 12127 10461
rect 12069 10452 12081 10455
rect 11563 10424 12081 10452
rect 11563 10421 11575 10424
rect 11517 10415 11575 10421
rect 12069 10421 12081 10424
rect 12115 10452 12127 10455
rect 12406 10452 12434 10492
rect 14642 10480 14648 10492
rect 14700 10480 14706 10532
rect 17252 10523 17310 10529
rect 17252 10489 17264 10523
rect 17298 10520 17310 10523
rect 17681 10523 17739 10529
rect 17681 10520 17693 10523
rect 17298 10492 17693 10520
rect 17298 10489 17310 10492
rect 17252 10483 17310 10489
rect 17681 10489 17693 10492
rect 17727 10489 17739 10523
rect 17681 10483 17739 10489
rect 20165 10523 20223 10529
rect 20165 10489 20177 10523
rect 20211 10520 20223 10523
rect 20438 10520 20444 10532
rect 20211 10492 20444 10520
rect 20211 10489 20223 10492
rect 20165 10483 20223 10489
rect 20438 10480 20444 10492
rect 20496 10480 20502 10532
rect 12115 10424 12434 10452
rect 12115 10421 12127 10424
rect 12069 10415 12127 10421
rect 13078 10412 13084 10464
rect 13136 10452 13142 10464
rect 13357 10455 13415 10461
rect 13357 10452 13369 10455
rect 13136 10424 13369 10452
rect 13136 10412 13142 10424
rect 13357 10421 13369 10424
rect 13403 10421 13415 10455
rect 13357 10415 13415 10421
rect 13446 10412 13452 10464
rect 13504 10452 13510 10464
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 13504 10424 14473 10452
rect 13504 10412 13510 10424
rect 14461 10421 14473 10424
rect 14507 10452 14519 10455
rect 17954 10452 17960 10464
rect 14507 10424 17960 10452
rect 14507 10421 14519 10424
rect 14461 10415 14519 10421
rect 17954 10412 17960 10424
rect 18012 10412 18018 10464
rect 18966 10452 18972 10464
rect 18927 10424 18972 10452
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 20254 10452 20260 10464
rect 20215 10424 20260 10452
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 9953 10251 10011 10257
rect 9953 10248 9965 10251
rect 9640 10220 9965 10248
rect 9640 10208 9646 10220
rect 9953 10217 9965 10220
rect 9999 10217 10011 10251
rect 13078 10248 13084 10260
rect 13039 10220 13084 10248
rect 9953 10211 10011 10217
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 13354 10208 13360 10260
rect 13412 10248 13418 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 13412 10220 13553 10248
rect 13412 10208 13418 10220
rect 13541 10217 13553 10220
rect 13587 10217 13599 10251
rect 13541 10211 13599 10217
rect 14642 10208 14648 10260
rect 14700 10248 14706 10260
rect 18966 10248 18972 10260
rect 14700 10220 18972 10248
rect 14700 10208 14706 10220
rect 18966 10208 18972 10220
rect 19024 10208 19030 10260
rect 20438 10248 20444 10260
rect 20399 10220 20444 10248
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 20901 10251 20959 10257
rect 20901 10217 20913 10251
rect 20947 10248 20959 10251
rect 20990 10248 20996 10260
rect 20947 10220 20996 10248
rect 20947 10217 20959 10220
rect 20901 10211 20959 10217
rect 20990 10208 20996 10220
rect 21048 10208 21054 10260
rect 8288 10183 8346 10189
rect 8288 10149 8300 10183
rect 8334 10180 8346 10183
rect 9398 10180 9404 10192
rect 8334 10152 9404 10180
rect 8334 10149 8346 10152
rect 8288 10143 8346 10149
rect 9398 10140 9404 10152
rect 9456 10140 9462 10192
rect 11088 10183 11146 10189
rect 11088 10149 11100 10183
rect 11134 10180 11146 10183
rect 11790 10180 11796 10192
rect 11134 10152 11796 10180
rect 11134 10149 11146 10152
rect 11088 10143 11146 10149
rect 11790 10140 11796 10152
rect 11848 10140 11854 10192
rect 13446 10180 13452 10192
rect 13359 10152 13452 10180
rect 13446 10140 13452 10152
rect 13504 10180 13510 10192
rect 14458 10180 14464 10192
rect 13504 10152 14464 10180
rect 13504 10140 13510 10152
rect 14458 10140 14464 10152
rect 14516 10140 14522 10192
rect 16666 10140 16672 10192
rect 16724 10180 16730 10192
rect 17586 10180 17592 10192
rect 16724 10152 17592 10180
rect 16724 10140 16730 10152
rect 17586 10140 17592 10152
rect 17644 10140 17650 10192
rect 8021 10115 8079 10121
rect 8021 10081 8033 10115
rect 8067 10112 8079 10115
rect 8110 10112 8116 10124
rect 8067 10084 8116 10112
rect 8067 10081 8079 10084
rect 8021 10075 8079 10081
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 11333 10115 11391 10121
rect 11333 10081 11345 10115
rect 11379 10112 11391 10115
rect 12434 10112 12440 10124
rect 11379 10084 12440 10112
rect 11379 10081 11391 10084
rect 11333 10075 11391 10081
rect 12434 10072 12440 10084
rect 12492 10112 12498 10124
rect 13722 10112 13728 10124
rect 12492 10084 13728 10112
rect 12492 10072 12498 10084
rect 13722 10072 13728 10084
rect 13780 10112 13786 10124
rect 13780 10084 13860 10112
rect 13780 10072 13786 10084
rect 13630 10044 13636 10056
rect 13591 10016 13636 10044
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 13832 10044 13860 10084
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 14349 10115 14407 10121
rect 14349 10112 14361 10115
rect 13964 10084 14361 10112
rect 13964 10072 13970 10084
rect 14349 10081 14361 10084
rect 14395 10081 14407 10115
rect 14349 10075 14407 10081
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 18785 10115 18843 10121
rect 18785 10112 18797 10115
rect 18104 10084 18797 10112
rect 18104 10072 18110 10084
rect 18785 10081 18797 10084
rect 18831 10081 18843 10115
rect 18785 10075 18843 10081
rect 19052 10115 19110 10121
rect 19052 10081 19064 10115
rect 19098 10112 19110 10115
rect 19886 10112 19892 10124
rect 19098 10084 19892 10112
rect 19098 10081 19110 10084
rect 19052 10075 19110 10081
rect 19886 10072 19892 10084
rect 19944 10072 19950 10124
rect 20162 10072 20168 10124
rect 20220 10112 20226 10124
rect 21085 10115 21143 10121
rect 21085 10112 21097 10115
rect 20220 10084 21097 10112
rect 20220 10072 20226 10084
rect 21085 10081 21097 10084
rect 21131 10081 21143 10115
rect 21085 10075 21143 10081
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13832 10016 14105 10044
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 9214 9936 9220 9988
rect 9272 9976 9278 9988
rect 9401 9979 9459 9985
rect 9401 9976 9413 9979
rect 9272 9948 9413 9976
rect 9272 9936 9278 9948
rect 9401 9945 9413 9948
rect 9447 9945 9459 9979
rect 9401 9939 9459 9945
rect 15378 9868 15384 9920
rect 15436 9908 15442 9920
rect 15473 9911 15531 9917
rect 15473 9908 15485 9911
rect 15436 9880 15485 9908
rect 15436 9868 15442 9880
rect 15473 9877 15485 9880
rect 15519 9877 15531 9911
rect 15473 9871 15531 9877
rect 20070 9868 20076 9920
rect 20128 9908 20134 9920
rect 20165 9911 20223 9917
rect 20165 9908 20177 9911
rect 20128 9880 20177 9908
rect 20128 9868 20134 9880
rect 20165 9877 20177 9880
rect 20211 9877 20223 9911
rect 20165 9871 20223 9877
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 8938 9664 8944 9716
rect 8996 9704 9002 9716
rect 9125 9707 9183 9713
rect 9125 9704 9137 9707
rect 8996 9676 9137 9704
rect 8996 9664 9002 9676
rect 9125 9673 9137 9676
rect 9171 9673 9183 9707
rect 11790 9704 11796 9716
rect 11751 9676 11796 9704
rect 9125 9667 9183 9673
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 13906 9704 13912 9716
rect 13867 9676 13912 9704
rect 13906 9664 13912 9676
rect 13964 9664 13970 9716
rect 17221 9707 17279 9713
rect 17221 9673 17233 9707
rect 17267 9704 17279 9707
rect 17862 9704 17868 9716
rect 17267 9676 17868 9704
rect 17267 9673 17279 9676
rect 17221 9667 17279 9673
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 19797 9707 19855 9713
rect 19797 9673 19809 9707
rect 19843 9704 19855 9707
rect 20254 9704 20260 9716
rect 19843 9676 20260 9704
rect 19843 9673 19855 9676
rect 19797 9667 19855 9673
rect 20254 9664 20260 9676
rect 20312 9664 20318 9716
rect 14366 9596 14372 9648
rect 14424 9636 14430 9648
rect 14829 9639 14887 9645
rect 14829 9636 14841 9639
rect 14424 9608 14841 9636
rect 14424 9596 14430 9608
rect 14829 9605 14841 9608
rect 14875 9605 14887 9639
rect 14829 9599 14887 9605
rect 20809 9639 20867 9645
rect 20809 9605 20821 9639
rect 20855 9636 20867 9639
rect 21082 9636 21088 9648
rect 20855 9608 21088 9636
rect 20855 9605 20867 9608
rect 20809 9599 20867 9605
rect 21082 9596 21088 9608
rect 21140 9596 21146 9648
rect 22002 9636 22008 9648
rect 21963 9608 22008 9636
rect 22002 9596 22008 9608
rect 22060 9596 22066 9648
rect 15378 9568 15384 9580
rect 13096 9540 15384 9568
rect 12894 9460 12900 9512
rect 12952 9509 12958 9512
rect 12952 9500 12964 9509
rect 13096 9500 13124 9540
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 20349 9571 20407 9577
rect 20349 9568 20361 9571
rect 19944 9540 20361 9568
rect 19944 9528 19950 9540
rect 20349 9537 20361 9540
rect 20395 9537 20407 9571
rect 20349 9531 20407 9537
rect 12952 9472 13124 9500
rect 13173 9503 13231 9509
rect 12952 9463 12964 9472
rect 13173 9469 13185 9503
rect 13219 9469 13231 9503
rect 13173 9463 13231 9469
rect 13449 9503 13507 9509
rect 13449 9469 13461 9503
rect 13495 9500 13507 9503
rect 13630 9500 13636 9512
rect 13495 9472 13636 9500
rect 13495 9469 13507 9472
rect 13449 9463 13507 9469
rect 12952 9460 12958 9463
rect 12434 9392 12440 9444
rect 12492 9432 12498 9444
rect 13188 9432 13216 9463
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 18046 9460 18052 9512
rect 18104 9500 18110 9512
rect 18601 9503 18659 9509
rect 18601 9500 18613 9503
rect 18104 9472 18613 9500
rect 18104 9460 18110 9472
rect 18601 9469 18613 9472
rect 18647 9469 18659 9503
rect 20990 9500 20996 9512
rect 20951 9472 20996 9500
rect 18601 9463 18659 9469
rect 20990 9460 20996 9472
rect 21048 9460 21054 9512
rect 12492 9404 13216 9432
rect 15197 9435 15255 9441
rect 12492 9392 12498 9404
rect 15197 9401 15209 9435
rect 15243 9432 15255 9435
rect 15841 9435 15899 9441
rect 15841 9432 15853 9435
rect 15243 9404 15853 9432
rect 15243 9401 15255 9404
rect 15197 9395 15255 9401
rect 15841 9401 15853 9404
rect 15887 9401 15899 9435
rect 15841 9395 15899 9401
rect 18356 9435 18414 9441
rect 18356 9401 18368 9435
rect 18402 9432 18414 9435
rect 20070 9432 20076 9444
rect 18402 9404 20076 9432
rect 18402 9401 18414 9404
rect 18356 9395 18414 9401
rect 20070 9392 20076 9404
rect 20128 9392 20134 9444
rect 20165 9435 20223 9441
rect 20165 9401 20177 9435
rect 20211 9432 20223 9435
rect 20346 9432 20352 9444
rect 20211 9404 20352 9432
rect 20211 9401 20223 9404
rect 20165 9395 20223 9401
rect 20346 9392 20352 9404
rect 20404 9392 20410 9444
rect 14458 9364 14464 9376
rect 14419 9336 14464 9364
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 15289 9367 15347 9373
rect 15289 9333 15301 9367
rect 15335 9364 15347 9367
rect 15746 9364 15752 9376
rect 15335 9336 15752 9364
rect 15335 9333 15347 9336
rect 15289 9327 15347 9333
rect 15746 9324 15752 9336
rect 15804 9364 15810 9376
rect 16390 9364 16396 9376
rect 15804 9336 16396 9364
rect 15804 9324 15810 9336
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 19242 9364 19248 9376
rect 19155 9336 19248 9364
rect 19242 9324 19248 9336
rect 19300 9364 19306 9376
rect 20257 9367 20315 9373
rect 20257 9364 20269 9367
rect 19300 9336 20269 9364
rect 19300 9324 19306 9336
rect 20257 9333 20269 9336
rect 20303 9333 20315 9367
rect 20257 9327 20315 9333
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 11882 9120 11888 9172
rect 11940 9120 11946 9172
rect 12066 9160 12072 9172
rect 12027 9132 12072 9160
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 15749 9163 15807 9169
rect 15749 9160 15761 9163
rect 12406 9132 15761 9160
rect 11900 9092 11928 9120
rect 12406 9092 12434 9132
rect 15749 9129 15761 9132
rect 15795 9129 15807 9163
rect 15749 9123 15807 9129
rect 20073 9163 20131 9169
rect 20073 9129 20085 9163
rect 20119 9160 20131 9163
rect 20162 9160 20168 9172
rect 20119 9132 20168 9160
rect 20119 9129 20131 9132
rect 20073 9123 20131 9129
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 20533 9163 20591 9169
rect 20533 9129 20545 9163
rect 20579 9160 20591 9163
rect 20990 9160 20996 9172
rect 20579 9132 20996 9160
rect 20579 9129 20591 9132
rect 20533 9123 20591 9129
rect 20990 9120 20996 9132
rect 21048 9120 21054 9172
rect 11900 9064 12434 9092
rect 11882 9024 11888 9036
rect 11843 8996 11888 9024
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16206 9024 16212 9036
rect 15979 8996 16212 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16206 8984 16212 8996
rect 16264 8984 16270 9036
rect 19613 9027 19671 9033
rect 19613 8993 19625 9027
rect 19659 9024 19671 9027
rect 19886 9024 19892 9036
rect 19659 8996 19892 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 19886 8984 19892 8996
rect 19944 8984 19950 9036
rect 20349 9027 20407 9033
rect 20349 8993 20361 9027
rect 20395 8993 20407 9027
rect 20990 9024 20996 9036
rect 20951 8996 20996 9024
rect 20349 8987 20407 8993
rect 20364 8956 20392 8987
rect 20990 8984 20996 8996
rect 21048 8984 21054 9036
rect 21358 8956 21364 8968
rect 20364 8928 21364 8956
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 17770 8848 17776 8900
rect 17828 8888 17834 8900
rect 20809 8891 20867 8897
rect 20809 8888 20821 8891
rect 17828 8860 20821 8888
rect 17828 8848 17834 8860
rect 20809 8857 20821 8860
rect 20855 8857 20867 8891
rect 20809 8851 20867 8857
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 11425 8619 11483 8625
rect 11425 8585 11437 8619
rect 11471 8616 11483 8619
rect 11882 8616 11888 8628
rect 11471 8588 11888 8616
rect 11471 8585 11483 8588
rect 11425 8579 11483 8585
rect 11882 8576 11888 8588
rect 11940 8576 11946 8628
rect 13262 8616 13268 8628
rect 13223 8588 13268 8616
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 16206 8616 16212 8628
rect 16167 8588 16212 8616
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 20073 8619 20131 8625
rect 20073 8585 20085 8619
rect 20119 8616 20131 8619
rect 20990 8616 20996 8628
rect 20119 8588 20996 8616
rect 20119 8585 20131 8588
rect 20073 8579 20131 8585
rect 20990 8576 20996 8588
rect 21048 8576 21054 8628
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8616 21419 8619
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21407 8588 22017 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 13725 8551 13783 8557
rect 13725 8517 13737 8551
rect 13771 8517 13783 8551
rect 13725 8511 13783 8517
rect 14553 8551 14611 8557
rect 14553 8517 14565 8551
rect 14599 8517 14611 8551
rect 20530 8548 20536 8560
rect 20491 8520 20536 8548
rect 14553 8511 14611 8517
rect 11238 8412 11244 8424
rect 11199 8384 11244 8412
rect 11238 8372 11244 8384
rect 11296 8372 11302 8424
rect 13449 8415 13507 8421
rect 13449 8381 13461 8415
rect 13495 8412 13507 8415
rect 13740 8412 13768 8511
rect 13495 8384 13768 8412
rect 13909 8415 13967 8421
rect 13495 8381 13507 8384
rect 13449 8375 13507 8381
rect 13909 8381 13921 8415
rect 13955 8412 13967 8415
rect 14568 8412 14596 8511
rect 20530 8508 20536 8520
rect 20588 8508 20594 8560
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 14700 8452 15117 8480
rect 14700 8440 14706 8452
rect 15105 8449 15117 8452
rect 15151 8449 15163 8483
rect 21376 8480 21404 8579
rect 15105 8443 15163 8449
rect 20364 8452 21404 8480
rect 13955 8384 14596 8412
rect 16393 8415 16451 8421
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 16393 8381 16405 8415
rect 16439 8412 16451 8415
rect 17126 8412 17132 8424
rect 16439 8384 17132 8412
rect 16439 8381 16451 8384
rect 16393 8375 16451 8381
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 19245 8415 19303 8421
rect 19245 8381 19257 8415
rect 19291 8412 19303 8415
rect 19886 8412 19892 8424
rect 19291 8384 19892 8412
rect 19291 8381 19303 8384
rect 19245 8375 19303 8381
rect 19886 8372 19892 8384
rect 19944 8372 19950 8424
rect 20364 8421 20392 8452
rect 20349 8415 20407 8421
rect 20349 8381 20361 8415
rect 20395 8381 20407 8415
rect 20349 8375 20407 8381
rect 20438 8372 20444 8424
rect 20496 8412 20502 8424
rect 20993 8415 21051 8421
rect 20993 8412 21005 8415
rect 20496 8384 21005 8412
rect 20496 8372 20502 8384
rect 20993 8381 21005 8384
rect 21039 8381 21051 8415
rect 20993 8375 21051 8381
rect 15013 8347 15071 8353
rect 15013 8313 15025 8347
rect 15059 8344 15071 8347
rect 15194 8344 15200 8356
rect 15059 8316 15200 8344
rect 15059 8313 15071 8316
rect 15013 8307 15071 8313
rect 15194 8304 15200 8316
rect 15252 8304 15258 8356
rect 17402 8304 17408 8356
rect 17460 8344 17466 8356
rect 17460 8316 20852 8344
rect 17460 8304 17466 8316
rect 14734 8236 14740 8288
rect 14792 8276 14798 8288
rect 14921 8279 14979 8285
rect 14921 8276 14933 8279
rect 14792 8248 14933 8276
rect 14792 8236 14798 8248
rect 14921 8245 14933 8248
rect 14967 8245 14979 8279
rect 17494 8276 17500 8288
rect 17455 8248 17500 8276
rect 14921 8239 14979 8245
rect 17494 8236 17500 8248
rect 17552 8236 17558 8288
rect 20824 8285 20852 8316
rect 20809 8279 20867 8285
rect 20809 8245 20821 8279
rect 20855 8245 20867 8279
rect 20809 8239 20867 8245
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 11885 8075 11943 8081
rect 11885 8072 11897 8075
rect 11296 8044 11897 8072
rect 11296 8032 11302 8044
rect 11885 8041 11897 8044
rect 11931 8041 11943 8075
rect 17126 8072 17132 8084
rect 17087 8044 17132 8072
rect 11885 8035 11943 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 17494 8072 17500 8084
rect 17455 8044 17500 8072
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 19613 8075 19671 8081
rect 19613 8041 19625 8075
rect 19659 8072 19671 8075
rect 19794 8072 19800 8084
rect 19659 8044 19800 8072
rect 19659 8041 19671 8044
rect 19613 8035 19671 8041
rect 19794 8032 19800 8044
rect 19852 8032 19858 8084
rect 20073 8075 20131 8081
rect 20073 8041 20085 8075
rect 20119 8072 20131 8075
rect 20438 8072 20444 8084
rect 20119 8044 20444 8072
rect 20119 8041 20131 8044
rect 20073 8035 20131 8041
rect 20438 8032 20444 8044
rect 20496 8032 20502 8084
rect 20533 8075 20591 8081
rect 20533 8041 20545 8075
rect 20579 8041 20591 8075
rect 20533 8035 20591 8041
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 12253 7939 12311 7945
rect 12253 7936 12265 7939
rect 11756 7908 12265 7936
rect 11756 7896 11762 7908
rect 12253 7905 12265 7908
rect 12299 7905 12311 7939
rect 12253 7899 12311 7905
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 13722 7936 13728 7948
rect 13679 7908 13728 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 13906 7945 13912 7948
rect 13900 7936 13912 7945
rect 13867 7908 13912 7936
rect 13900 7899 13912 7908
rect 13906 7896 13912 7899
rect 13964 7896 13970 7948
rect 18138 7936 18144 7948
rect 17788 7908 18144 7936
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 12345 7871 12403 7877
rect 12345 7868 12357 7871
rect 11940 7840 12357 7868
rect 11940 7828 11946 7840
rect 12345 7837 12357 7840
rect 12391 7837 12403 7871
rect 12345 7831 12403 7837
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7837 12495 7871
rect 17586 7868 17592 7880
rect 17547 7840 17592 7868
rect 12437 7831 12495 7837
rect 12158 7760 12164 7812
rect 12216 7800 12222 7812
rect 12452 7800 12480 7831
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 17788 7877 17816 7908
rect 18138 7896 18144 7908
rect 18196 7936 18202 7948
rect 18489 7939 18547 7945
rect 18489 7936 18501 7939
rect 18196 7908 18501 7936
rect 18196 7896 18202 7908
rect 18489 7905 18501 7908
rect 18535 7905 18547 7939
rect 19886 7936 19892 7948
rect 19847 7908 19892 7936
rect 18489 7899 18547 7905
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 20349 7939 20407 7945
rect 20349 7905 20361 7939
rect 20395 7905 20407 7939
rect 20548 7936 20576 8035
rect 20993 7939 21051 7945
rect 20993 7936 21005 7939
rect 20548 7908 21005 7936
rect 20349 7899 20407 7905
rect 20993 7905 21005 7908
rect 21039 7905 21051 7939
rect 20993 7899 21051 7905
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7837 17831 7871
rect 17773 7831 17831 7837
rect 18046 7828 18052 7880
rect 18104 7868 18110 7880
rect 18233 7871 18291 7877
rect 18233 7868 18245 7871
rect 18104 7840 18245 7868
rect 18104 7828 18110 7840
rect 18233 7837 18245 7840
rect 18279 7837 18291 7871
rect 20364 7868 20392 7899
rect 20364 7840 21404 7868
rect 18233 7831 18291 7837
rect 12216 7772 12480 7800
rect 12216 7760 12222 7772
rect 21376 7744 21404 7840
rect 14642 7692 14648 7744
rect 14700 7732 14706 7744
rect 15010 7732 15016 7744
rect 14700 7704 15016 7732
rect 14700 7692 14706 7704
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 20809 7735 20867 7741
rect 20809 7732 20821 7735
rect 16080 7704 20821 7732
rect 16080 7692 16086 7704
rect 20809 7701 20821 7704
rect 20855 7701 20867 7735
rect 21358 7732 21364 7744
rect 21319 7704 21364 7732
rect 20809 7695 20867 7701
rect 21358 7692 21364 7704
rect 21416 7692 21422 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 15562 7488 15568 7540
rect 15620 7528 15626 7540
rect 15620 7500 18092 7528
rect 15620 7488 15626 7500
rect 18064 7460 18092 7500
rect 18138 7488 18144 7540
rect 18196 7528 18202 7540
rect 18417 7531 18475 7537
rect 18417 7528 18429 7531
rect 18196 7500 18429 7528
rect 18196 7488 18202 7500
rect 18417 7497 18429 7500
rect 18463 7497 18475 7531
rect 18417 7491 18475 7497
rect 19886 7488 19892 7540
rect 19944 7528 19950 7540
rect 19981 7531 20039 7537
rect 19981 7528 19993 7531
rect 19944 7500 19993 7528
rect 19944 7488 19950 7500
rect 19981 7497 19993 7500
rect 20027 7497 20039 7531
rect 20809 7531 20867 7537
rect 20809 7528 20821 7531
rect 19981 7491 20039 7497
rect 20088 7500 20821 7528
rect 20088 7460 20116 7500
rect 20809 7497 20821 7500
rect 20855 7497 20867 7531
rect 20809 7491 20867 7497
rect 18064 7432 20116 7460
rect 20533 7463 20591 7469
rect 20533 7429 20545 7463
rect 20579 7429 20591 7463
rect 20533 7423 20591 7429
rect 11609 7395 11667 7401
rect 11609 7361 11621 7395
rect 11655 7392 11667 7395
rect 11698 7392 11704 7404
rect 11655 7364 11704 7392
rect 11655 7361 11667 7364
rect 11609 7355 11667 7361
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 14734 7392 14740 7404
rect 14695 7364 14740 7392
rect 14734 7352 14740 7364
rect 14792 7352 14798 7404
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 8260 7296 9689 7324
rect 8260 7284 8266 7296
rect 9677 7293 9689 7296
rect 9723 7293 9735 7327
rect 9677 7287 9735 7293
rect 11885 7327 11943 7333
rect 11885 7293 11897 7327
rect 11931 7324 11943 7327
rect 11931 7296 12434 7324
rect 11931 7293 11943 7296
rect 11885 7287 11943 7293
rect 9950 7265 9956 7268
rect 9944 7256 9956 7265
rect 9911 7228 9956 7256
rect 9944 7219 9956 7228
rect 9950 7216 9956 7219
rect 10008 7216 10014 7268
rect 12158 7265 12164 7268
rect 12130 7259 12164 7265
rect 12130 7256 12142 7259
rect 11072 7228 12142 7256
rect 11072 7197 11100 7228
rect 12130 7225 12142 7228
rect 12216 7256 12222 7268
rect 12406 7256 12434 7296
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 15381 7327 15439 7333
rect 15381 7324 15393 7327
rect 13780 7296 15393 7324
rect 13780 7284 13786 7296
rect 15381 7293 15393 7296
rect 15427 7324 15439 7327
rect 17037 7327 17095 7333
rect 17037 7324 17049 7327
rect 15427 7296 17049 7324
rect 15427 7293 15439 7296
rect 15381 7287 15439 7293
rect 17037 7293 17049 7296
rect 17083 7293 17095 7327
rect 17037 7287 17095 7293
rect 20349 7327 20407 7333
rect 20349 7293 20361 7327
rect 20395 7293 20407 7327
rect 20548 7324 20576 7423
rect 20993 7327 21051 7333
rect 20993 7324 21005 7327
rect 20548 7296 21005 7324
rect 20349 7287 20407 7293
rect 20993 7293 21005 7296
rect 21039 7293 21051 7327
rect 20993 7287 21051 7293
rect 13740 7256 13768 7284
rect 12216 7228 12278 7256
rect 12406 7228 13768 7256
rect 12130 7219 12164 7225
rect 12158 7216 12164 7219
rect 12216 7216 12222 7228
rect 15010 7216 15016 7268
rect 15068 7256 15074 7268
rect 15626 7259 15684 7265
rect 15626 7256 15638 7259
rect 15068 7228 15638 7256
rect 15068 7216 15074 7228
rect 15626 7225 15638 7228
rect 15672 7225 15684 7259
rect 17304 7259 17362 7265
rect 17304 7256 17316 7259
rect 15626 7219 15684 7225
rect 16776 7228 17316 7256
rect 11057 7191 11115 7197
rect 11057 7157 11069 7191
rect 11103 7157 11115 7191
rect 11057 7151 11115 7157
rect 13265 7191 13323 7197
rect 13265 7157 13277 7191
rect 13311 7188 13323 7191
rect 13906 7188 13912 7200
rect 13311 7160 13912 7188
rect 13311 7157 13323 7160
rect 13265 7151 13323 7157
rect 13906 7148 13912 7160
rect 13964 7188 13970 7200
rect 14550 7188 14556 7200
rect 13964 7160 14556 7188
rect 13964 7148 13970 7160
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 16776 7197 16804 7228
rect 17304 7225 17316 7228
rect 17350 7256 17362 7259
rect 18230 7256 18236 7268
rect 17350 7228 18236 7256
rect 17350 7225 17362 7228
rect 17304 7219 17362 7225
rect 18230 7216 18236 7228
rect 18288 7216 18294 7268
rect 20364 7256 20392 7287
rect 20364 7228 21404 7256
rect 21376 7200 21404 7228
rect 16761 7191 16819 7197
rect 16761 7157 16773 7191
rect 16807 7157 16819 7191
rect 21358 7188 21364 7200
rect 21319 7160 21364 7188
rect 16761 7151 16819 7157
rect 21358 7148 21364 7160
rect 21416 7148 21422 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 11882 6984 11888 6996
rect 11843 6956 11888 6984
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12253 6987 12311 6993
rect 12253 6953 12265 6987
rect 12299 6984 12311 6987
rect 12299 6956 17540 6984
rect 12299 6953 12311 6956
rect 12253 6947 12311 6953
rect 14829 6919 14887 6925
rect 14829 6885 14841 6919
rect 14875 6916 14887 6919
rect 16482 6916 16488 6928
rect 14875 6888 16488 6916
rect 14875 6885 14887 6888
rect 14829 6879 14887 6885
rect 16482 6876 16488 6888
rect 16540 6876 16546 6928
rect 17512 6916 17540 6956
rect 17586 6944 17592 6996
rect 17644 6984 17650 6996
rect 17681 6987 17739 6993
rect 17681 6984 17693 6987
rect 17644 6956 17693 6984
rect 17644 6944 17650 6956
rect 17681 6953 17693 6956
rect 17727 6953 17739 6987
rect 17681 6947 17739 6953
rect 18049 6987 18107 6993
rect 18049 6953 18061 6987
rect 18095 6984 18107 6987
rect 20349 6987 20407 6993
rect 20349 6984 20361 6987
rect 18095 6956 20361 6984
rect 18095 6953 18107 6956
rect 18049 6947 18107 6953
rect 20349 6953 20361 6956
rect 20395 6953 20407 6987
rect 20349 6947 20407 6953
rect 21174 6916 21180 6928
rect 17512 6888 21180 6916
rect 21174 6876 21180 6888
rect 21232 6876 21238 6928
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 8461 6851 8519 6857
rect 8461 6848 8473 6851
rect 5684 6820 8473 6848
rect 5684 6808 5690 6820
rect 8461 6817 8473 6820
rect 8507 6817 8519 6851
rect 8461 6811 8519 6817
rect 11333 6851 11391 6857
rect 11333 6817 11345 6851
rect 11379 6848 11391 6851
rect 12342 6848 12348 6860
rect 11379 6820 12348 6848
rect 11379 6817 11391 6820
rect 11333 6811 11391 6817
rect 12342 6808 12348 6820
rect 12400 6848 12406 6860
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 12400 6820 14197 6848
rect 12400 6808 12406 6820
rect 14185 6817 14197 6820
rect 14231 6848 14243 6851
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 14231 6820 14749 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 14737 6817 14749 6820
rect 14783 6848 14795 6851
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 14783 6820 17417 6848
rect 14783 6817 14795 6820
rect 14737 6811 14795 6817
rect 17405 6817 17417 6820
rect 17451 6848 17463 6851
rect 18141 6851 18199 6857
rect 18141 6848 18153 6851
rect 17451 6820 18153 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 18141 6817 18153 6820
rect 18187 6848 18199 6851
rect 19242 6848 19248 6860
rect 18187 6820 19248 6848
rect 18187 6817 18199 6820
rect 18141 6811 18199 6817
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 20073 6851 20131 6857
rect 20073 6817 20085 6851
rect 20119 6848 20131 6851
rect 20530 6848 20536 6860
rect 20119 6820 20536 6848
rect 20119 6817 20131 6820
rect 20073 6811 20131 6817
rect 20530 6808 20536 6820
rect 20588 6808 20594 6860
rect 20898 6808 20904 6860
rect 20956 6848 20962 6860
rect 20993 6851 21051 6857
rect 20993 6848 21005 6851
rect 20956 6820 21005 6848
rect 20956 6808 20962 6820
rect 20993 6817 21005 6820
rect 21039 6817 21051 6851
rect 20993 6811 21051 6817
rect 8202 6780 8208 6792
rect 8163 6752 8208 6780
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6749 12495 6783
rect 14550 6780 14556 6792
rect 14511 6752 14556 6780
rect 12437 6743 12495 6749
rect 9585 6715 9643 6721
rect 9585 6681 9597 6715
rect 9631 6712 9643 6715
rect 9950 6712 9956 6724
rect 9631 6684 9956 6712
rect 9631 6681 9643 6684
rect 9585 6675 9643 6681
rect 9950 6672 9956 6684
rect 10008 6712 10014 6724
rect 12452 6712 12480 6743
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 18230 6780 18236 6792
rect 18191 6752 18236 6780
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 15194 6712 15200 6724
rect 10008 6684 12480 6712
rect 15155 6684 15200 6712
rect 10008 6672 10014 6684
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 20809 6647 20867 6653
rect 20809 6644 20821 6647
rect 14332 6616 20821 6644
rect 14332 6604 14338 6616
rect 20809 6613 20821 6616
rect 20855 6613 20867 6647
rect 21358 6644 21364 6656
rect 21319 6616 21364 6644
rect 20809 6607 20867 6613
rect 21358 6604 21364 6616
rect 21416 6604 21422 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 20898 6440 20904 6452
rect 20859 6412 20904 6440
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 16482 6332 16488 6384
rect 16540 6372 16546 6384
rect 21177 6375 21235 6381
rect 21177 6372 21189 6375
rect 16540 6344 21189 6372
rect 16540 6332 16546 6344
rect 21177 6341 21189 6344
rect 21223 6341 21235 6375
rect 21177 6335 21235 6341
rect 20441 6239 20499 6245
rect 20441 6205 20453 6239
rect 20487 6236 20499 6239
rect 20714 6236 20720 6248
rect 20487 6208 20720 6236
rect 20487 6205 20499 6208
rect 20441 6199 20499 6205
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 21358 6236 21364 6248
rect 21319 6208 21364 6236
rect 21358 6196 21364 6208
rect 21416 6196 21422 6248
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1765 5899 1823 5905
rect 1765 5865 1777 5899
rect 1811 5896 1823 5899
rect 5626 5896 5632 5908
rect 1811 5868 5632 5896
rect 1811 5865 1823 5868
rect 1765 5859 1823 5865
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 12986 5788 12992 5840
rect 13044 5828 13050 5840
rect 20809 5831 20867 5837
rect 20809 5828 20821 5831
rect 13044 5800 20821 5828
rect 13044 5788 13050 5800
rect 20809 5797 20821 5800
rect 20855 5797 20867 5831
rect 20809 5791 20867 5797
rect 1578 5760 1584 5772
rect 1539 5732 1584 5760
rect 1578 5720 1584 5732
rect 1636 5760 1642 5772
rect 2041 5763 2099 5769
rect 2041 5760 2053 5763
rect 1636 5732 2053 5760
rect 1636 5720 1642 5732
rect 2041 5729 2053 5732
rect 2087 5729 2099 5763
rect 20990 5760 20996 5772
rect 20951 5732 20996 5760
rect 2041 5723 2099 5729
rect 20990 5720 20996 5732
rect 21048 5720 21054 5772
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 20901 5355 20959 5361
rect 20901 5321 20913 5355
rect 20947 5352 20959 5355
rect 20990 5352 20996 5364
rect 20947 5324 20996 5352
rect 20947 5321 20959 5324
rect 20901 5315 20959 5321
rect 20990 5312 20996 5324
rect 21048 5312 21054 5364
rect 21174 5352 21180 5364
rect 21135 5324 21180 5352
rect 21174 5312 21180 5324
rect 21232 5312 21238 5364
rect 20441 5151 20499 5157
rect 20441 5117 20453 5151
rect 20487 5148 20499 5151
rect 20714 5148 20720 5160
rect 20487 5120 20720 5148
rect 20487 5117 20499 5120
rect 20441 5111 20499 5117
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 21358 5148 21364 5160
rect 21319 5120 21364 5148
rect 21358 5108 21364 5120
rect 21416 5108 21422 5160
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 19978 4768 19984 4820
rect 20036 4808 20042 4820
rect 20809 4811 20867 4817
rect 20809 4808 20821 4811
rect 20036 4780 20821 4808
rect 20036 4768 20042 4780
rect 20809 4777 20821 4780
rect 20855 4777 20867 4811
rect 20809 4771 20867 4777
rect 21358 4740 21364 4752
rect 21319 4712 21364 4740
rect 21358 4700 21364 4712
rect 21416 4700 21422 4752
rect 20990 4672 20996 4684
rect 20951 4644 20996 4672
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 20809 4267 20867 4273
rect 20809 4233 20821 4267
rect 20855 4264 20867 4267
rect 20990 4264 20996 4276
rect 20855 4236 20996 4264
rect 20855 4233 20867 4236
rect 20809 4227 20867 4233
rect 20990 4224 20996 4236
rect 21048 4224 21054 4276
rect 18782 4088 18788 4140
rect 18840 4128 18846 4140
rect 21085 4131 21143 4137
rect 21085 4128 21097 4131
rect 18840 4100 21097 4128
rect 18840 4088 18846 4100
rect 21085 4097 21097 4100
rect 21131 4097 21143 4131
rect 21085 4091 21143 4097
rect 20349 4063 20407 4069
rect 20349 4029 20361 4063
rect 20395 4060 20407 4063
rect 20622 4060 20628 4072
rect 20395 4032 20628 4060
rect 20395 4029 20407 4032
rect 20349 4023 20407 4029
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 19981 3995 20039 4001
rect 19981 3961 19993 3995
rect 20027 3992 20039 3995
rect 21266 3992 21272 4004
rect 20027 3964 21272 3992
rect 20027 3961 20039 3964
rect 19981 3955 20039 3961
rect 21266 3952 21272 3964
rect 21324 3952 21330 4004
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 20625 3723 20683 3729
rect 20625 3720 20637 3723
rect 18012 3692 20637 3720
rect 18012 3680 18018 3692
rect 20625 3689 20637 3692
rect 20671 3689 20683 3723
rect 20625 3683 20683 3689
rect 16390 3612 16396 3664
rect 16448 3652 16454 3664
rect 21085 3655 21143 3661
rect 21085 3652 21097 3655
rect 16448 3624 21097 3652
rect 16448 3612 16454 3624
rect 21085 3621 21097 3624
rect 21131 3621 21143 3655
rect 21085 3615 21143 3621
rect 19337 3587 19395 3593
rect 19337 3553 19349 3587
rect 19383 3584 19395 3587
rect 20622 3584 20628 3596
rect 19383 3556 20628 3584
rect 19383 3553 19395 3556
rect 19337 3547 19395 3553
rect 20622 3544 20628 3556
rect 20680 3584 20686 3596
rect 20717 3587 20775 3593
rect 20717 3584 20729 3587
rect 20680 3556 20729 3584
rect 20680 3544 20686 3556
rect 20717 3553 20729 3556
rect 20763 3553 20775 3587
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 20717 3547 20775 3553
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3516 20315 3519
rect 21284 3516 21312 3544
rect 20303 3488 21312 3516
rect 20303 3485 20315 3488
rect 20257 3479 20315 3485
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19613 3383 19671 3389
rect 19613 3380 19625 3383
rect 19484 3352 19625 3380
rect 19484 3340 19490 3352
rect 19613 3349 19625 3352
rect 19659 3349 19671 3383
rect 19613 3343 19671 3349
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 18690 3136 18696 3188
rect 18748 3176 18754 3188
rect 20625 3179 20683 3185
rect 20625 3176 20637 3179
rect 18748 3148 20637 3176
rect 18748 3136 18754 3148
rect 20625 3145 20637 3148
rect 20671 3145 20683 3179
rect 20625 3139 20683 3145
rect 19334 3068 19340 3120
rect 19392 3108 19398 3120
rect 19981 3111 20039 3117
rect 19981 3108 19993 3111
rect 19392 3080 19993 3108
rect 19392 3068 19398 3080
rect 19981 3077 19993 3080
rect 20027 3077 20039 3111
rect 19981 3071 20039 3077
rect 19245 3043 19303 3049
rect 19245 3009 19257 3043
rect 19291 3040 19303 3043
rect 20901 3043 20959 3049
rect 20901 3040 20913 3043
rect 19291 3012 20913 3040
rect 19291 3009 19303 3012
rect 19245 3003 19303 3009
rect 20901 3009 20913 3012
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 19705 2975 19763 2981
rect 19705 2941 19717 2975
rect 19751 2972 19763 2975
rect 19751 2944 21312 2972
rect 19751 2941 19763 2944
rect 19705 2935 19763 2941
rect 21284 2916 21312 2944
rect 18877 2907 18935 2913
rect 18877 2873 18889 2907
rect 18923 2904 18935 2907
rect 20162 2904 20168 2916
rect 18923 2876 20168 2904
rect 18923 2873 18935 2876
rect 18877 2867 18935 2873
rect 20162 2864 20168 2876
rect 20220 2864 20226 2916
rect 20714 2904 20720 2916
rect 20627 2876 20720 2904
rect 20714 2864 20720 2876
rect 20772 2904 20778 2916
rect 20901 2907 20959 2913
rect 20901 2904 20913 2907
rect 20772 2876 20913 2904
rect 20772 2864 20778 2876
rect 20901 2873 20913 2876
rect 20947 2873 20959 2907
rect 21266 2904 21272 2916
rect 21227 2876 21272 2904
rect 20901 2867 20959 2873
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 18966 2796 18972 2848
rect 19024 2836 19030 2848
rect 21177 2839 21235 2845
rect 21177 2836 21189 2839
rect 19024 2808 21189 2836
rect 19024 2796 19030 2808
rect 21177 2805 21189 2808
rect 21223 2805 21235 2839
rect 21177 2799 21235 2805
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 18598 2592 18604 2644
rect 18656 2632 18662 2644
rect 20625 2635 20683 2641
rect 20625 2632 20637 2635
rect 18656 2604 20637 2632
rect 18656 2592 18662 2604
rect 20625 2601 20637 2604
rect 20671 2601 20683 2635
rect 20625 2595 20683 2601
rect 18969 2567 19027 2573
rect 18969 2533 18981 2567
rect 19015 2564 19027 2567
rect 20717 2567 20775 2573
rect 20717 2564 20729 2567
rect 19015 2536 20729 2564
rect 19015 2533 19027 2536
rect 18969 2527 19027 2533
rect 20717 2533 20729 2536
rect 20763 2564 20775 2567
rect 22005 2567 22063 2573
rect 22005 2564 22017 2567
rect 20763 2536 22017 2564
rect 20763 2533 20775 2536
rect 20717 2527 20775 2533
rect 22005 2533 22017 2536
rect 22051 2533 22063 2567
rect 22005 2527 22063 2533
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 19245 2499 19303 2505
rect 19245 2496 19257 2499
rect 17460 2468 19257 2496
rect 17460 2456 17466 2468
rect 19245 2465 19257 2468
rect 19291 2465 19303 2499
rect 19426 2496 19432 2508
rect 19387 2468 19432 2496
rect 19245 2459 19303 2465
rect 19426 2456 19432 2468
rect 19484 2456 19490 2508
rect 21266 2496 21272 2508
rect 21227 2468 21272 2496
rect 21266 2456 21272 2468
rect 21324 2456 21330 2508
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2428 20315 2431
rect 21284 2428 21312 2456
rect 20303 2400 21312 2428
rect 20303 2397 20315 2400
rect 20257 2391 20315 2397
rect 14458 2320 14464 2372
rect 14516 2360 14522 2372
rect 21085 2363 21143 2369
rect 21085 2360 21097 2363
rect 14516 2332 21097 2360
rect 14516 2320 14522 2332
rect 21085 2329 21097 2332
rect 21131 2329 21143 2363
rect 21085 2323 21143 2329
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 22002 1408 22008 1420
rect 21963 1380 22008 1408
rect 22002 1368 22008 1380
rect 22060 1368 22066 1420
<< via1 >>
rect 3056 20816 3108 20868
rect 4252 20816 4304 20868
rect 4712 20816 4764 20868
rect 5448 20816 5500 20868
rect 4160 20748 4212 20800
rect 5540 20748 5592 20800
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 6736 20544 6788 20596
rect 6920 20544 6972 20596
rect 8852 20544 8904 20596
rect 14280 20544 14332 20596
rect 18144 20544 18196 20596
rect 19432 20544 19484 20596
rect 20996 20544 21048 20596
rect 1400 20476 1452 20528
rect 848 20408 900 20460
rect 296 20340 348 20392
rect 1308 20340 1360 20392
rect 2044 20340 2096 20392
rect 2504 20340 2556 20392
rect 3608 20476 3660 20528
rect 5172 20476 5224 20528
rect 7748 20476 7800 20528
rect 8208 20476 8260 20528
rect 11796 20476 11848 20528
rect 12072 20519 12124 20528
rect 12072 20485 12081 20519
rect 12081 20485 12115 20519
rect 12115 20485 12124 20519
rect 12072 20476 12124 20485
rect 12624 20519 12676 20528
rect 12624 20485 12633 20519
rect 12633 20485 12667 20519
rect 12667 20485 12676 20519
rect 12624 20476 12676 20485
rect 13176 20519 13228 20528
rect 13176 20485 13185 20519
rect 13185 20485 13219 20519
rect 13219 20485 13228 20519
rect 13176 20476 13228 20485
rect 13728 20519 13780 20528
rect 13728 20485 13737 20519
rect 13737 20485 13771 20519
rect 13771 20485 13780 20519
rect 13728 20476 13780 20485
rect 17684 20476 17736 20528
rect 17960 20476 18012 20528
rect 18604 20476 18656 20528
rect 18788 20476 18840 20528
rect 18972 20519 19024 20528
rect 18972 20485 18981 20519
rect 18981 20485 19015 20519
rect 19015 20485 19024 20519
rect 18972 20476 19024 20485
rect 19524 20519 19576 20528
rect 19524 20485 19533 20519
rect 19533 20485 19567 20519
rect 19567 20485 19576 20519
rect 19524 20476 19576 20485
rect 2780 20408 2832 20460
rect 3792 20408 3844 20460
rect 4160 20408 4212 20460
rect 1952 20272 2004 20324
rect 2872 20272 2924 20324
rect 4252 20340 4304 20392
rect 5080 20340 5132 20392
rect 5448 20408 5500 20460
rect 5356 20340 5408 20392
rect 5540 20340 5592 20392
rect 6828 20408 6880 20460
rect 12256 20408 12308 20460
rect 6460 20340 6512 20392
rect 6920 20340 6972 20392
rect 7104 20340 7156 20392
rect 7564 20340 7616 20392
rect 8300 20383 8352 20392
rect 8300 20349 8309 20383
rect 8309 20349 8343 20383
rect 8343 20349 8352 20383
rect 8300 20340 8352 20349
rect 8668 20340 8720 20392
rect 9128 20340 9180 20392
rect 9220 20340 9272 20392
rect 9772 20340 9824 20392
rect 10324 20383 10376 20392
rect 10324 20349 10333 20383
rect 10333 20349 10367 20383
rect 10367 20349 10376 20383
rect 10324 20340 10376 20349
rect 10876 20340 10928 20392
rect 15844 20340 15896 20392
rect 16212 20340 16264 20392
rect 1768 20247 1820 20256
rect 1768 20213 1777 20247
rect 1777 20213 1811 20247
rect 1811 20213 1820 20247
rect 1768 20204 1820 20213
rect 2320 20247 2372 20256
rect 2320 20213 2329 20247
rect 2329 20213 2363 20247
rect 2363 20213 2372 20247
rect 2320 20204 2372 20213
rect 4620 20204 4672 20256
rect 4896 20204 4948 20256
rect 5448 20247 5500 20256
rect 5448 20213 5457 20247
rect 5457 20213 5491 20247
rect 5491 20213 5500 20247
rect 5448 20204 5500 20213
rect 6092 20247 6144 20256
rect 6092 20213 6101 20247
rect 6101 20213 6135 20247
rect 6135 20213 6144 20247
rect 6092 20204 6144 20213
rect 11244 20272 11296 20324
rect 11888 20272 11940 20324
rect 12164 20272 12216 20324
rect 12900 20272 12952 20324
rect 13268 20272 13320 20324
rect 7472 20204 7524 20256
rect 7656 20204 7708 20256
rect 8668 20247 8720 20256
rect 8668 20213 8677 20247
rect 8677 20213 8711 20247
rect 8711 20213 8720 20247
rect 8668 20204 8720 20213
rect 9588 20247 9640 20256
rect 9588 20213 9597 20247
rect 9597 20213 9631 20247
rect 9631 20213 9640 20247
rect 9588 20204 9640 20213
rect 10876 20204 10928 20256
rect 14188 20204 14240 20256
rect 14372 20204 14424 20256
rect 17592 20272 17644 20324
rect 18144 20272 18196 20324
rect 18604 20272 18656 20324
rect 19524 20340 19576 20392
rect 20260 20383 20312 20392
rect 20260 20349 20269 20383
rect 20269 20349 20303 20383
rect 20303 20349 20312 20383
rect 20260 20340 20312 20349
rect 20536 20340 20588 20392
rect 18880 20272 18932 20324
rect 19432 20204 19484 20256
rect 20168 20272 20220 20324
rect 20812 20315 20864 20324
rect 20812 20281 20821 20315
rect 20821 20281 20855 20315
rect 20855 20281 20864 20315
rect 20812 20272 20864 20281
rect 21364 20315 21416 20324
rect 21364 20281 21373 20315
rect 21373 20281 21407 20315
rect 21407 20281 21416 20315
rect 21364 20272 21416 20281
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 1308 20000 1360 20052
rect 2044 20043 2096 20052
rect 2044 20009 2053 20043
rect 2053 20009 2087 20043
rect 2087 20009 2096 20043
rect 2044 20000 2096 20009
rect 2504 20043 2556 20052
rect 2504 20009 2513 20043
rect 2513 20009 2547 20043
rect 2547 20009 2556 20043
rect 2504 20000 2556 20009
rect 2872 20043 2924 20052
rect 2872 20009 2881 20043
rect 2881 20009 2915 20043
rect 2915 20009 2924 20043
rect 2872 20000 2924 20009
rect 3792 20043 3844 20052
rect 3792 20009 3801 20043
rect 3801 20009 3835 20043
rect 3835 20009 3844 20043
rect 3792 20000 3844 20009
rect 5448 20000 5500 20052
rect 6828 20043 6880 20052
rect 6828 20009 6837 20043
rect 6837 20009 6871 20043
rect 6871 20009 6880 20043
rect 6828 20000 6880 20009
rect 8300 20000 8352 20052
rect 10324 20000 10376 20052
rect 16304 20000 16356 20052
rect 16580 20000 16632 20052
rect 19340 20000 19392 20052
rect 4712 19932 4764 19984
rect 5080 19932 5132 19984
rect 5356 19932 5408 19984
rect 5816 19932 5868 19984
rect 1768 19864 1820 19916
rect 4252 19839 4304 19848
rect 4252 19805 4261 19839
rect 4261 19805 4295 19839
rect 4295 19805 4304 19839
rect 4252 19796 4304 19805
rect 4804 19864 4856 19916
rect 5264 19864 5316 19916
rect 5724 19864 5776 19916
rect 6460 19932 6512 19984
rect 6736 19864 6788 19916
rect 7840 19907 7892 19916
rect 5172 19796 5224 19848
rect 4620 19728 4672 19780
rect 4896 19703 4948 19712
rect 4896 19669 4905 19703
rect 4905 19669 4939 19703
rect 4939 19669 4948 19703
rect 4896 19660 4948 19669
rect 7840 19873 7874 19907
rect 7874 19873 7892 19907
rect 7840 19864 7892 19873
rect 7196 19796 7248 19848
rect 8576 19660 8628 19712
rect 8944 19703 8996 19712
rect 8944 19669 8953 19703
rect 8953 19669 8987 19703
rect 8987 19669 8996 19703
rect 8944 19660 8996 19669
rect 9772 19932 9824 19984
rect 10876 19932 10928 19984
rect 15200 19932 15252 19984
rect 15384 19932 15436 19984
rect 15936 19932 15988 19984
rect 9220 19864 9272 19916
rect 11704 19864 11756 19916
rect 14648 19907 14700 19916
rect 14648 19873 14657 19907
rect 14657 19873 14691 19907
rect 14691 19873 14700 19907
rect 14648 19864 14700 19873
rect 15568 19864 15620 19916
rect 16028 19907 16080 19916
rect 16028 19873 16037 19907
rect 16037 19873 16071 19907
rect 16071 19873 16080 19907
rect 16028 19864 16080 19873
rect 17408 19864 17460 19916
rect 17776 19864 17828 19916
rect 19708 19932 19760 19984
rect 20352 19932 20404 19984
rect 19616 19864 19668 19916
rect 20628 19864 20680 19916
rect 9680 19796 9732 19848
rect 10968 19796 11020 19848
rect 14832 19796 14884 19848
rect 16580 19839 16632 19848
rect 16580 19805 16589 19839
rect 16589 19805 16623 19839
rect 16623 19805 16632 19839
rect 16580 19796 16632 19805
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 18696 19796 18748 19805
rect 19892 19796 19944 19848
rect 9128 19728 9180 19780
rect 11244 19728 11296 19780
rect 11152 19660 11204 19712
rect 12900 19660 12952 19712
rect 16672 19728 16724 19780
rect 21364 19771 21416 19780
rect 21364 19737 21373 19771
rect 21373 19737 21407 19771
rect 21407 19737 21416 19771
rect 21364 19728 21416 19737
rect 16764 19660 16816 19712
rect 17592 19660 17644 19712
rect 20996 19660 21048 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 7104 19456 7156 19508
rect 7748 19456 7800 19508
rect 12348 19456 12400 19508
rect 7840 19388 7892 19440
rect 14280 19456 14332 19508
rect 18604 19499 18656 19508
rect 18604 19465 18613 19499
rect 18613 19465 18647 19499
rect 18647 19465 18656 19499
rect 18604 19456 18656 19465
rect 20536 19456 20588 19508
rect 6920 19320 6972 19372
rect 3884 19252 3936 19304
rect 4804 19252 4856 19304
rect 5908 19295 5960 19304
rect 4252 19184 4304 19236
rect 4804 19116 4856 19168
rect 5908 19261 5917 19295
rect 5917 19261 5951 19295
rect 5951 19261 5960 19295
rect 5908 19252 5960 19261
rect 7196 19252 7248 19304
rect 8668 19320 8720 19372
rect 8944 19320 8996 19372
rect 9404 19363 9456 19372
rect 9404 19329 9413 19363
rect 9413 19329 9447 19363
rect 9447 19329 9456 19363
rect 9404 19320 9456 19329
rect 9680 19295 9732 19304
rect 9680 19261 9689 19295
rect 9689 19261 9723 19295
rect 9723 19261 9732 19295
rect 9680 19252 9732 19261
rect 6644 19184 6696 19236
rect 8944 19184 8996 19236
rect 10876 19252 10928 19304
rect 15844 19388 15896 19440
rect 13176 19252 13228 19304
rect 14556 19295 14608 19304
rect 14556 19261 14565 19295
rect 14565 19261 14599 19295
rect 14599 19261 14608 19295
rect 14556 19252 14608 19261
rect 14832 19295 14884 19304
rect 14832 19261 14866 19295
rect 14866 19261 14884 19295
rect 14832 19252 14884 19261
rect 16672 19320 16724 19372
rect 20168 19388 20220 19440
rect 19892 19320 19944 19372
rect 16580 19295 16632 19304
rect 11336 19184 11388 19236
rect 11980 19116 12032 19168
rect 12072 19116 12124 19168
rect 13820 19159 13872 19168
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 15844 19116 15896 19168
rect 16580 19261 16589 19295
rect 16589 19261 16623 19295
rect 16623 19261 16632 19295
rect 16580 19252 16632 19261
rect 17040 19252 17092 19304
rect 17500 19252 17552 19304
rect 19064 19295 19116 19304
rect 17316 19184 17368 19236
rect 19064 19261 19073 19295
rect 19073 19261 19107 19295
rect 19107 19261 19116 19295
rect 19064 19252 19116 19261
rect 20076 19252 20128 19304
rect 20444 19295 20496 19304
rect 20444 19261 20453 19295
rect 20453 19261 20487 19295
rect 20487 19261 20496 19295
rect 20444 19252 20496 19261
rect 16948 19159 17000 19168
rect 16948 19125 16957 19159
rect 16957 19125 16991 19159
rect 16991 19125 17000 19159
rect 16948 19116 17000 19125
rect 17040 19116 17092 19168
rect 20536 19184 20588 19236
rect 20904 19184 20956 19236
rect 21364 19227 21416 19236
rect 21364 19193 21373 19227
rect 21373 19193 21407 19227
rect 21407 19193 21416 19227
rect 21364 19184 21416 19193
rect 21548 19116 21600 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 4252 18912 4304 18964
rect 4896 18912 4948 18964
rect 5540 18912 5592 18964
rect 7564 18912 7616 18964
rect 11336 18955 11388 18964
rect 11336 18921 11345 18955
rect 11345 18921 11379 18955
rect 11379 18921 11388 18955
rect 11336 18912 11388 18921
rect 11980 18912 12032 18964
rect 14740 18955 14792 18964
rect 6736 18844 6788 18896
rect 1768 18776 1820 18828
rect 7196 18819 7248 18828
rect 7196 18785 7205 18819
rect 7205 18785 7239 18819
rect 7239 18785 7248 18819
rect 7196 18776 7248 18785
rect 10232 18819 10284 18828
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 7288 18708 7340 18760
rect 10232 18785 10266 18819
rect 10266 18785 10284 18819
rect 10232 18776 10284 18785
rect 11796 18776 11848 18828
rect 12440 18776 12492 18828
rect 13176 18776 13228 18828
rect 13820 18844 13872 18896
rect 14740 18921 14749 18955
rect 14749 18921 14783 18955
rect 14783 18921 14792 18955
rect 14740 18912 14792 18921
rect 17040 18912 17092 18964
rect 17500 18955 17552 18964
rect 17500 18921 17509 18955
rect 17509 18921 17543 18955
rect 17543 18921 17552 18955
rect 17500 18912 17552 18921
rect 18144 18912 18196 18964
rect 19524 18955 19576 18964
rect 19524 18921 19533 18955
rect 19533 18921 19567 18955
rect 19567 18921 19576 18955
rect 19524 18912 19576 18921
rect 22652 18912 22704 18964
rect 12072 18751 12124 18760
rect 3884 18572 3936 18624
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 8944 18615 8996 18624
rect 8944 18581 8953 18615
rect 8953 18581 8987 18615
rect 8987 18581 8996 18615
rect 8944 18572 8996 18581
rect 12072 18717 12081 18751
rect 12081 18717 12115 18751
rect 12115 18717 12124 18751
rect 12072 18708 12124 18717
rect 13084 18751 13136 18760
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 13084 18708 13136 18717
rect 16948 18776 17000 18828
rect 22100 18844 22152 18896
rect 18052 18819 18104 18828
rect 18052 18785 18061 18819
rect 18061 18785 18095 18819
rect 18095 18785 18104 18819
rect 18052 18776 18104 18785
rect 19064 18776 19116 18828
rect 19248 18819 19300 18828
rect 19248 18785 19257 18819
rect 19257 18785 19291 18819
rect 19291 18785 19300 18819
rect 19248 18776 19300 18785
rect 19708 18819 19760 18828
rect 19708 18785 19717 18819
rect 19717 18785 19751 18819
rect 19751 18785 19760 18819
rect 19708 18776 19760 18785
rect 19984 18776 20036 18828
rect 20444 18776 20496 18828
rect 21180 18819 21232 18828
rect 21180 18785 21189 18819
rect 21189 18785 21223 18819
rect 21223 18785 21232 18819
rect 21180 18776 21232 18785
rect 18604 18708 18656 18760
rect 20260 18640 20312 18692
rect 21364 18683 21416 18692
rect 21364 18649 21373 18683
rect 21373 18649 21407 18683
rect 21407 18649 21416 18683
rect 21364 18640 21416 18649
rect 10968 18572 11020 18624
rect 13360 18572 13412 18624
rect 14648 18572 14700 18624
rect 17316 18572 17368 18624
rect 21088 18572 21140 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 6644 18411 6696 18420
rect 6644 18377 6653 18411
rect 6653 18377 6687 18411
rect 6687 18377 6696 18411
rect 6644 18368 6696 18377
rect 7196 18368 7248 18420
rect 8944 18368 8996 18420
rect 18052 18368 18104 18420
rect 19800 18368 19852 18420
rect 20628 18368 20680 18420
rect 21180 18368 21232 18420
rect 12716 18300 12768 18352
rect 11244 18232 11296 18284
rect 13820 18300 13872 18352
rect 13360 18275 13412 18284
rect 13360 18241 13369 18275
rect 13369 18241 13403 18275
rect 13403 18241 13412 18275
rect 13360 18232 13412 18241
rect 14556 18232 14608 18284
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 18328 18275 18380 18284
rect 18328 18241 18337 18275
rect 18337 18241 18371 18275
rect 18371 18241 18380 18275
rect 18328 18232 18380 18241
rect 19340 18232 19392 18284
rect 5264 18207 5316 18216
rect 5264 18173 5273 18207
rect 5273 18173 5307 18207
rect 5307 18173 5316 18207
rect 5264 18164 5316 18173
rect 5908 18164 5960 18216
rect 7288 18207 7340 18216
rect 7288 18173 7297 18207
rect 7297 18173 7331 18207
rect 7331 18173 7340 18207
rect 7288 18164 7340 18173
rect 5540 18139 5592 18148
rect 5540 18105 5574 18139
rect 5574 18105 5592 18139
rect 5540 18096 5592 18105
rect 9404 18164 9456 18216
rect 13084 18164 13136 18216
rect 15844 18207 15896 18216
rect 15844 18173 15878 18207
rect 15878 18173 15896 18207
rect 18604 18207 18656 18216
rect 15844 18164 15896 18173
rect 18604 18173 18613 18207
rect 18613 18173 18647 18207
rect 18647 18173 18656 18207
rect 18604 18164 18656 18173
rect 20168 18207 20220 18216
rect 20168 18173 20177 18207
rect 20177 18173 20211 18207
rect 20211 18173 20220 18207
rect 20168 18164 20220 18173
rect 10968 18096 11020 18148
rect 14188 18096 14240 18148
rect 20260 18096 20312 18148
rect 21364 18139 21416 18148
rect 21364 18105 21373 18139
rect 21373 18105 21407 18139
rect 21407 18105 21416 18139
rect 21364 18096 21416 18105
rect 7380 18071 7432 18080
rect 7380 18037 7389 18071
rect 7389 18037 7423 18071
rect 7423 18037 7432 18071
rect 7380 18028 7432 18037
rect 9772 18028 9824 18080
rect 10232 18028 10284 18080
rect 11244 18071 11296 18080
rect 11244 18037 11253 18071
rect 11253 18037 11287 18071
rect 11287 18037 11296 18071
rect 11244 18028 11296 18037
rect 12440 18028 12492 18080
rect 16488 18028 16540 18080
rect 17592 18071 17644 18080
rect 17592 18037 17601 18071
rect 17601 18037 17635 18071
rect 17635 18037 17644 18071
rect 17592 18028 17644 18037
rect 19064 18028 19116 18080
rect 19800 18028 19852 18080
rect 19984 18028 20036 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 3608 17867 3660 17876
rect 3608 17833 3617 17867
rect 3617 17833 3651 17867
rect 3651 17833 3660 17867
rect 3608 17824 3660 17833
rect 5724 17867 5776 17876
rect 5724 17833 5733 17867
rect 5733 17833 5767 17867
rect 5767 17833 5776 17867
rect 5724 17824 5776 17833
rect 7380 17824 7432 17876
rect 9588 17824 9640 17876
rect 11244 17824 11296 17876
rect 7748 17688 7800 17740
rect 8484 17688 8536 17740
rect 9128 17688 9180 17740
rect 18328 17824 18380 17876
rect 19708 17824 19760 17876
rect 20260 17867 20312 17876
rect 20260 17833 20269 17867
rect 20269 17833 20303 17867
rect 20303 17833 20312 17867
rect 20260 17824 20312 17833
rect 17316 17756 17368 17808
rect 17592 17756 17644 17808
rect 16488 17688 16540 17740
rect 3700 17663 3752 17672
rect 3700 17629 3709 17663
rect 3709 17629 3743 17663
rect 3743 17629 3752 17663
rect 3700 17620 3752 17629
rect 5540 17620 5592 17672
rect 7656 17620 7708 17672
rect 9772 17663 9824 17672
rect 9772 17629 9781 17663
rect 9781 17629 9815 17663
rect 9815 17629 9824 17663
rect 9772 17620 9824 17629
rect 17132 17663 17184 17672
rect 17132 17629 17141 17663
rect 17141 17629 17175 17663
rect 17175 17629 17184 17663
rect 17132 17620 17184 17629
rect 18144 17620 18196 17672
rect 12440 17552 12492 17604
rect 20628 17731 20680 17740
rect 20628 17697 20637 17731
rect 20637 17697 20671 17731
rect 20671 17697 20680 17731
rect 20628 17688 20680 17697
rect 20720 17688 20772 17740
rect 20812 17595 20864 17604
rect 20812 17561 20821 17595
rect 20821 17561 20855 17595
rect 20855 17561 20864 17595
rect 20812 17552 20864 17561
rect 21364 17595 21416 17604
rect 21364 17561 21373 17595
rect 21373 17561 21407 17595
rect 21407 17561 21416 17595
rect 21364 17552 21416 17561
rect 1676 17527 1728 17536
rect 1676 17493 1685 17527
rect 1685 17493 1719 17527
rect 1719 17493 1728 17527
rect 1676 17484 1728 17493
rect 3056 17484 3108 17536
rect 7748 17484 7800 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 1768 17323 1820 17332
rect 1768 17289 1777 17323
rect 1777 17289 1811 17323
rect 1811 17289 1820 17323
rect 1768 17280 1820 17289
rect 3516 17280 3568 17332
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 7472 17144 7524 17153
rect 8484 17187 8536 17196
rect 8484 17153 8493 17187
rect 8493 17153 8527 17187
rect 8527 17153 8536 17187
rect 8484 17144 8536 17153
rect 11244 17144 11296 17196
rect 12532 17144 12584 17196
rect 3884 17076 3936 17128
rect 4252 17076 4304 17128
rect 6092 17076 6144 17128
rect 11152 17076 11204 17128
rect 2872 17051 2924 17060
rect 2872 17017 2912 17051
rect 2912 17017 2924 17051
rect 2872 17008 2924 17017
rect 3700 17008 3752 17060
rect 12440 17008 12492 17060
rect 15200 17144 15252 17196
rect 18144 17280 18196 17332
rect 19248 17323 19300 17332
rect 19248 17289 19257 17323
rect 19257 17289 19291 17323
rect 19291 17289 19300 17323
rect 19248 17280 19300 17289
rect 20628 17323 20680 17332
rect 20628 17289 20637 17323
rect 20637 17289 20671 17323
rect 20671 17289 20680 17323
rect 20628 17280 20680 17289
rect 19708 17144 19760 17196
rect 19064 17119 19116 17128
rect 8300 16940 8352 16992
rect 12624 16983 12676 16992
rect 12624 16949 12633 16983
rect 12633 16949 12667 16983
rect 12667 16949 12676 16983
rect 12624 16940 12676 16949
rect 14740 16940 14792 16992
rect 19064 17085 19073 17119
rect 19073 17085 19107 17119
rect 19107 17085 19116 17119
rect 19064 17076 19116 17085
rect 19432 16940 19484 16992
rect 21180 17051 21232 17060
rect 21180 17017 21189 17051
rect 21189 17017 21223 17051
rect 21223 17017 21232 17051
rect 21180 17008 21232 17017
rect 21456 17008 21508 17060
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 3056 16779 3108 16788
rect 3056 16745 3065 16779
rect 3065 16745 3099 16779
rect 3099 16745 3108 16779
rect 3056 16736 3108 16745
rect 3516 16779 3568 16788
rect 3516 16745 3525 16779
rect 3525 16745 3559 16779
rect 3559 16745 3568 16779
rect 3516 16736 3568 16745
rect 4804 16711 4856 16720
rect 4804 16677 4838 16711
rect 4838 16677 4856 16711
rect 8300 16736 8352 16788
rect 4804 16668 4856 16677
rect 7472 16668 7524 16720
rect 3884 16600 3936 16652
rect 5264 16600 5316 16652
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 12624 16736 12676 16788
rect 14280 16736 14332 16788
rect 14740 16736 14792 16788
rect 19340 16736 19392 16788
rect 19432 16736 19484 16788
rect 20720 16736 20772 16788
rect 21180 16736 21232 16788
rect 1768 16532 1820 16584
rect 9404 16532 9456 16584
rect 12532 16600 12584 16652
rect 14648 16600 14700 16652
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 14556 16532 14608 16584
rect 15292 16600 15344 16652
rect 15936 16600 15988 16652
rect 18696 16643 18748 16652
rect 18696 16609 18705 16643
rect 18705 16609 18739 16643
rect 18739 16609 18748 16643
rect 18696 16600 18748 16609
rect 19708 16643 19760 16652
rect 19708 16609 19717 16643
rect 19717 16609 19751 16643
rect 19751 16609 19760 16643
rect 19708 16600 19760 16609
rect 21180 16643 21232 16652
rect 21180 16609 21189 16643
rect 21189 16609 21223 16643
rect 21223 16609 21232 16643
rect 21180 16600 21232 16609
rect 21364 16643 21416 16652
rect 21364 16609 21373 16643
rect 21373 16609 21407 16643
rect 21407 16609 21416 16643
rect 21364 16600 21416 16609
rect 14556 16396 14608 16448
rect 16580 16439 16632 16448
rect 16580 16405 16589 16439
rect 16589 16405 16623 16439
rect 16623 16405 16632 16439
rect 16580 16396 16632 16405
rect 20260 16396 20312 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 5540 16192 5592 16244
rect 11244 16192 11296 16244
rect 12532 16192 12584 16244
rect 15936 16235 15988 16244
rect 15936 16201 15945 16235
rect 15945 16201 15979 16235
rect 15979 16201 15988 16235
rect 15936 16192 15988 16201
rect 16672 16192 16724 16244
rect 17592 16192 17644 16244
rect 18696 16192 18748 16244
rect 20168 16192 20220 16244
rect 21180 16192 21232 16244
rect 7288 16056 7340 16108
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 16580 16056 16632 16108
rect 17960 16099 18012 16108
rect 17960 16065 17969 16099
rect 17969 16065 18003 16099
rect 18003 16065 18012 16099
rect 17960 16056 18012 16065
rect 7472 15988 7524 16040
rect 9404 15988 9456 16040
rect 11244 16031 11296 16040
rect 11244 15997 11278 16031
rect 11278 15997 11296 16031
rect 11244 15988 11296 15997
rect 16120 15988 16172 16040
rect 20260 15988 20312 16040
rect 6092 15920 6144 15972
rect 14280 15920 14332 15972
rect 16764 15920 16816 15972
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 20812 15920 20864 15972
rect 21364 15963 21416 15972
rect 21364 15929 21373 15963
rect 21373 15929 21407 15963
rect 21407 15929 21416 15963
rect 21364 15920 21416 15929
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 2872 15648 2924 15700
rect 16120 15648 16172 15700
rect 17960 15648 18012 15700
rect 20812 15691 20864 15700
rect 20812 15657 20821 15691
rect 20821 15657 20855 15691
rect 20855 15657 20864 15691
rect 20812 15648 20864 15657
rect 3884 15580 3936 15632
rect 10968 15580 11020 15632
rect 2504 15512 2556 15564
rect 9312 15512 9364 15564
rect 6092 15444 6144 15496
rect 7748 15444 7800 15496
rect 4804 15376 4856 15428
rect 16580 15512 16632 15564
rect 20352 15580 20404 15632
rect 14556 15444 14608 15496
rect 17132 15487 17184 15496
rect 17132 15453 17141 15487
rect 17141 15453 17175 15487
rect 17175 15453 17184 15487
rect 17132 15444 17184 15453
rect 21364 15419 21416 15428
rect 21364 15385 21373 15419
rect 21373 15385 21407 15419
rect 21407 15385 21416 15419
rect 21364 15376 21416 15385
rect 7288 15308 7340 15360
rect 9128 15351 9180 15360
rect 9128 15317 9137 15351
rect 9137 15317 9171 15351
rect 9171 15317 9180 15351
rect 9128 15308 9180 15317
rect 9588 15308 9640 15360
rect 14648 15308 14700 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 4804 15147 4856 15156
rect 4804 15113 4813 15147
rect 4813 15113 4847 15147
rect 4847 15113 4856 15147
rect 4804 15104 4856 15113
rect 6092 15147 6144 15156
rect 6092 15113 6101 15147
rect 6101 15113 6135 15147
rect 6135 15113 6144 15147
rect 6092 15104 6144 15113
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 14556 15104 14608 15156
rect 14740 15147 14792 15156
rect 14740 15113 14749 15147
rect 14749 15113 14783 15147
rect 14783 15113 14792 15147
rect 14740 15104 14792 15113
rect 20352 15147 20404 15156
rect 20352 15113 20361 15147
rect 20361 15113 20395 15147
rect 20395 15113 20404 15147
rect 20352 15104 20404 15113
rect 7564 15036 7616 15088
rect 2504 14968 2556 15020
rect 8208 15011 8260 15020
rect 8208 14977 8217 15011
rect 8217 14977 8251 15011
rect 8251 14977 8260 15011
rect 8208 14968 8260 14977
rect 7472 14943 7524 14952
rect 7472 14909 7481 14943
rect 7481 14909 7515 14943
rect 7515 14909 7524 14943
rect 7472 14900 7524 14909
rect 7196 14875 7248 14884
rect 7196 14841 7214 14875
rect 7214 14841 7248 14875
rect 14004 14968 14056 15020
rect 17132 14968 17184 15020
rect 11060 14900 11112 14952
rect 14556 14943 14608 14952
rect 14556 14909 14565 14943
rect 14565 14909 14599 14943
rect 14599 14909 14608 14943
rect 14556 14900 14608 14909
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 20536 14900 20588 14952
rect 7196 14832 7248 14841
rect 17868 14832 17920 14884
rect 17960 14832 18012 14884
rect 4252 14764 4304 14816
rect 8300 14764 8352 14816
rect 9128 14764 9180 14816
rect 9312 14807 9364 14816
rect 9312 14773 9321 14807
rect 9321 14773 9355 14807
rect 9355 14773 9364 14807
rect 9312 14764 9364 14773
rect 12624 14807 12676 14816
rect 12624 14773 12633 14807
rect 12633 14773 12667 14807
rect 12667 14773 12676 14807
rect 12624 14764 12676 14773
rect 12716 14807 12768 14816
rect 12716 14773 12725 14807
rect 12725 14773 12759 14807
rect 12759 14773 12768 14807
rect 13084 14807 13136 14816
rect 12716 14764 12768 14773
rect 13084 14773 13093 14807
rect 13093 14773 13127 14807
rect 13127 14773 13136 14807
rect 13084 14764 13136 14773
rect 13176 14764 13228 14816
rect 18604 14764 18656 14816
rect 19156 14807 19208 14816
rect 19156 14773 19165 14807
rect 19165 14773 19199 14807
rect 19199 14773 19208 14807
rect 19156 14764 19208 14773
rect 21364 14875 21416 14884
rect 21364 14841 21373 14875
rect 21373 14841 21407 14875
rect 21407 14841 21416 14875
rect 21364 14832 21416 14841
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 2504 14603 2556 14612
rect 2504 14569 2513 14603
rect 2513 14569 2547 14603
rect 2547 14569 2556 14603
rect 2504 14560 2556 14569
rect 4252 14603 4304 14612
rect 4252 14569 4261 14603
rect 4261 14569 4295 14603
rect 4295 14569 4304 14603
rect 4252 14560 4304 14569
rect 4988 14560 5040 14612
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 8300 14492 8352 14544
rect 12256 14560 12308 14612
rect 12624 14603 12676 14612
rect 12624 14569 12633 14603
rect 12633 14569 12667 14603
rect 12667 14569 12676 14603
rect 12624 14560 12676 14569
rect 13084 14560 13136 14612
rect 17868 14560 17920 14612
rect 20904 14560 20956 14612
rect 20168 14492 20220 14544
rect 4160 14424 4212 14476
rect 3884 14399 3936 14408
rect 3884 14365 3893 14399
rect 3893 14365 3927 14399
rect 3927 14365 3936 14399
rect 3884 14356 3936 14365
rect 9496 14467 9548 14476
rect 8484 14399 8536 14408
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 8484 14356 8536 14365
rect 9496 14433 9505 14467
rect 9505 14433 9539 14467
rect 9539 14433 9548 14467
rect 9496 14424 9548 14433
rect 9588 14424 9640 14476
rect 14004 14424 14056 14476
rect 14924 14424 14976 14476
rect 15660 14467 15712 14476
rect 15660 14433 15669 14467
rect 15669 14433 15703 14467
rect 15703 14433 15712 14467
rect 15660 14424 15712 14433
rect 18604 14424 18656 14476
rect 19340 14424 19392 14476
rect 9680 14356 9732 14408
rect 12164 14356 12216 14408
rect 12256 14288 12308 14340
rect 9036 14263 9088 14272
rect 9036 14229 9045 14263
rect 9045 14229 9079 14263
rect 9079 14229 9088 14263
rect 9036 14220 9088 14229
rect 13360 14220 13412 14272
rect 18696 14356 18748 14408
rect 18052 14288 18104 14340
rect 19156 14288 19208 14340
rect 20444 14356 20496 14408
rect 21272 14331 21324 14340
rect 21272 14297 21281 14331
rect 21281 14297 21315 14331
rect 21315 14297 21324 14331
rect 21272 14288 21324 14297
rect 16396 14220 16448 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 4160 14059 4212 14068
rect 4160 14025 4169 14059
rect 4169 14025 4203 14059
rect 4203 14025 4212 14059
rect 4160 14016 4212 14025
rect 8668 14016 8720 14068
rect 11060 14059 11112 14068
rect 11060 14025 11069 14059
rect 11069 14025 11103 14059
rect 11103 14025 11112 14059
rect 11060 14016 11112 14025
rect 12808 14016 12860 14068
rect 14004 14059 14056 14068
rect 14004 14025 14013 14059
rect 14013 14025 14047 14059
rect 14047 14025 14056 14059
rect 14004 14016 14056 14025
rect 15660 14059 15712 14068
rect 15660 14025 15669 14059
rect 15669 14025 15703 14059
rect 15703 14025 15712 14059
rect 15660 14016 15712 14025
rect 20536 14016 20588 14068
rect 12164 13880 12216 13932
rect 7472 13812 7524 13864
rect 8208 13744 8260 13796
rect 8484 13744 8536 13796
rect 9588 13744 9640 13796
rect 17132 13880 17184 13932
rect 21364 13923 21416 13932
rect 21364 13889 21373 13923
rect 21373 13889 21407 13923
rect 21407 13889 21416 13923
rect 21364 13880 21416 13889
rect 14740 13812 14792 13864
rect 16396 13855 16448 13864
rect 16396 13821 16405 13855
rect 16405 13821 16439 13855
rect 16439 13821 16448 13855
rect 16396 13812 16448 13821
rect 18052 13812 18104 13864
rect 18880 13812 18932 13864
rect 20536 13812 20588 13864
rect 18604 13744 18656 13796
rect 21180 13787 21232 13796
rect 21180 13753 21189 13787
rect 21189 13753 21223 13787
rect 21223 13753 21232 13787
rect 21180 13744 21232 13753
rect 13176 13676 13228 13728
rect 15200 13719 15252 13728
rect 15200 13685 15209 13719
rect 15209 13685 15243 13719
rect 15243 13685 15252 13719
rect 15200 13676 15252 13685
rect 18696 13719 18748 13728
rect 18696 13685 18705 13719
rect 18705 13685 18739 13719
rect 18739 13685 18748 13719
rect 18696 13676 18748 13685
rect 20628 13719 20680 13728
rect 20628 13685 20637 13719
rect 20637 13685 20671 13719
rect 20671 13685 20680 13719
rect 20628 13676 20680 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 7196 13472 7248 13524
rect 9036 13472 9088 13524
rect 9496 13472 9548 13524
rect 12532 13515 12584 13524
rect 12532 13481 12541 13515
rect 12541 13481 12575 13515
rect 12575 13481 12584 13515
rect 12532 13472 12584 13481
rect 12716 13472 12768 13524
rect 14556 13472 14608 13524
rect 15200 13472 15252 13524
rect 15752 13472 15804 13524
rect 16488 13472 16540 13524
rect 18880 13515 18932 13524
rect 18880 13481 18889 13515
rect 18889 13481 18923 13515
rect 18923 13481 18932 13515
rect 18880 13472 18932 13481
rect 19156 13472 19208 13524
rect 19340 13515 19392 13524
rect 19340 13481 19349 13515
rect 19349 13481 19383 13515
rect 19383 13481 19392 13515
rect 19340 13472 19392 13481
rect 20352 13515 20404 13524
rect 20352 13481 20361 13515
rect 20361 13481 20395 13515
rect 20395 13481 20404 13515
rect 20352 13472 20404 13481
rect 18696 13404 18748 13456
rect 21364 13447 21416 13456
rect 21364 13413 21373 13447
rect 21373 13413 21407 13447
rect 21407 13413 21416 13447
rect 21364 13404 21416 13413
rect 9772 13336 9824 13388
rect 12256 13336 12308 13388
rect 12440 13336 12492 13388
rect 8208 13268 8260 13320
rect 8668 13311 8720 13320
rect 8668 13277 8677 13311
rect 8677 13277 8711 13311
rect 8711 13277 8720 13311
rect 8668 13268 8720 13277
rect 9588 13175 9640 13184
rect 9588 13141 9597 13175
rect 9597 13141 9631 13175
rect 9631 13141 9640 13175
rect 9588 13132 9640 13141
rect 12164 13268 12216 13320
rect 12808 13336 12860 13388
rect 20628 13336 20680 13388
rect 12716 13268 12768 13320
rect 13636 13268 13688 13320
rect 18052 13268 18104 13320
rect 20352 13268 20404 13320
rect 20904 13336 20956 13388
rect 20076 13200 20128 13252
rect 13544 13132 13596 13184
rect 16304 13132 16356 13184
rect 18604 13132 18656 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 9772 12971 9824 12980
rect 9772 12937 9781 12971
rect 9781 12937 9815 12971
rect 9815 12937 9824 12971
rect 9772 12928 9824 12937
rect 12164 12971 12216 12980
rect 12164 12937 12173 12971
rect 12173 12937 12207 12971
rect 12207 12937 12216 12971
rect 12164 12928 12216 12937
rect 15292 12860 15344 12912
rect 9588 12792 9640 12844
rect 16396 12835 16448 12844
rect 16396 12801 16405 12835
rect 16405 12801 16439 12835
rect 16439 12801 16448 12835
rect 16396 12792 16448 12801
rect 12440 12724 12492 12776
rect 13912 12724 13964 12776
rect 16304 12767 16356 12776
rect 16304 12733 16313 12767
rect 16313 12733 16347 12767
rect 16347 12733 16356 12767
rect 16304 12724 16356 12733
rect 17132 12792 17184 12844
rect 17316 12792 17368 12844
rect 17500 12792 17552 12844
rect 20352 12928 20404 12980
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 21180 12971 21232 12980
rect 21180 12937 21189 12971
rect 21189 12937 21223 12971
rect 21223 12937 21232 12971
rect 21180 12928 21232 12937
rect 20444 12903 20496 12912
rect 20444 12869 20453 12903
rect 20453 12869 20487 12903
rect 20487 12869 20496 12903
rect 20444 12860 20496 12869
rect 17684 12724 17736 12776
rect 19800 12767 19852 12776
rect 19800 12733 19809 12767
rect 19809 12733 19843 12767
rect 19843 12733 19852 12767
rect 19800 12724 19852 12733
rect 10692 12588 10744 12640
rect 11060 12699 11112 12708
rect 11060 12665 11094 12699
rect 11094 12665 11112 12699
rect 11060 12656 11112 12665
rect 15200 12656 15252 12708
rect 11152 12588 11204 12640
rect 15936 12631 15988 12640
rect 15936 12597 15945 12631
rect 15945 12597 15979 12631
rect 15979 12597 15988 12631
rect 15936 12588 15988 12597
rect 16580 12656 16632 12708
rect 17132 12656 17184 12708
rect 20444 12724 20496 12776
rect 17500 12588 17552 12640
rect 18972 12588 19024 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 10692 12427 10744 12436
rect 10692 12393 10701 12427
rect 10701 12393 10735 12427
rect 10735 12393 10744 12427
rect 10692 12384 10744 12393
rect 11152 12384 11204 12436
rect 15200 12384 15252 12436
rect 15936 12384 15988 12436
rect 16580 12427 16632 12436
rect 16580 12393 16589 12427
rect 16589 12393 16623 12427
rect 16623 12393 16632 12427
rect 16580 12384 16632 12393
rect 15292 12316 15344 12368
rect 18972 12316 19024 12368
rect 20168 12384 20220 12436
rect 20628 12384 20680 12436
rect 9312 12248 9364 12300
rect 11704 12248 11756 12300
rect 12440 12248 12492 12300
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 8944 12112 8996 12164
rect 8208 12044 8260 12096
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 17592 12223 17644 12232
rect 17592 12189 17601 12223
rect 17601 12189 17635 12223
rect 17635 12189 17644 12223
rect 17592 12180 17644 12189
rect 17684 12180 17736 12232
rect 17868 12180 17920 12232
rect 19248 12248 19300 12300
rect 20076 12180 20128 12232
rect 20444 12112 20496 12164
rect 19340 12044 19392 12096
rect 19616 12044 19668 12096
rect 20628 12044 20680 12096
rect 21364 12087 21416 12096
rect 21364 12053 21373 12087
rect 21373 12053 21407 12087
rect 21407 12053 21416 12087
rect 21364 12044 21416 12053
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 11704 11883 11756 11892
rect 11704 11849 11713 11883
rect 11713 11849 11747 11883
rect 11747 11849 11756 11883
rect 11704 11840 11756 11849
rect 13360 11840 13412 11892
rect 13636 11840 13688 11892
rect 15292 11840 15344 11892
rect 17316 11840 17368 11892
rect 18788 11840 18840 11892
rect 20076 11883 20128 11892
rect 20076 11849 20085 11883
rect 20085 11849 20119 11883
rect 20119 11849 20128 11883
rect 20076 11840 20128 11849
rect 20260 11840 20312 11892
rect 11060 11747 11112 11756
rect 11060 11713 11069 11747
rect 11069 11713 11103 11747
rect 11103 11713 11112 11747
rect 11060 11704 11112 11713
rect 13084 11704 13136 11756
rect 13636 11704 13688 11756
rect 2320 11636 2372 11688
rect 8208 11636 8260 11688
rect 15936 11679 15988 11688
rect 15936 11645 15965 11679
rect 15965 11645 15988 11679
rect 15936 11636 15988 11645
rect 9220 11568 9272 11620
rect 13728 11568 13780 11620
rect 9772 11500 9824 11552
rect 11336 11543 11388 11552
rect 11336 11509 11345 11543
rect 11345 11509 11379 11543
rect 11379 11509 11388 11543
rect 13176 11543 13228 11552
rect 11336 11500 11388 11509
rect 13176 11509 13185 11543
rect 13185 11509 13219 11543
rect 13219 11509 13228 11543
rect 13176 11500 13228 11509
rect 13452 11500 13504 11552
rect 18696 11636 18748 11688
rect 19064 11636 19116 11688
rect 18052 11500 18104 11552
rect 21364 11636 21416 11688
rect 21364 11543 21416 11552
rect 21364 11509 21373 11543
rect 21373 11509 21407 11543
rect 21407 11509 21416 11543
rect 21364 11500 21416 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 9772 11339 9824 11348
rect 9772 11305 9781 11339
rect 9781 11305 9815 11339
rect 9815 11305 9824 11339
rect 9772 11296 9824 11305
rect 11336 11296 11388 11348
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 19064 11339 19116 11348
rect 19064 11305 19073 11339
rect 19073 11305 19107 11339
rect 19107 11305 19116 11339
rect 19064 11296 19116 11305
rect 8852 11228 8904 11280
rect 9680 11228 9732 11280
rect 16304 11228 16356 11280
rect 18972 11228 19024 11280
rect 20628 11296 20680 11348
rect 9404 11203 9456 11212
rect 9404 11169 9413 11203
rect 9413 11169 9447 11203
rect 9447 11169 9456 11203
rect 9404 11160 9456 11169
rect 10784 11203 10836 11212
rect 10784 11169 10793 11203
rect 10793 11169 10827 11203
rect 10827 11169 10836 11203
rect 10784 11160 10836 11169
rect 14372 11160 14424 11212
rect 14556 11203 14608 11212
rect 14556 11169 14565 11203
rect 14565 11169 14599 11203
rect 14599 11169 14608 11203
rect 14556 11160 14608 11169
rect 16488 11160 16540 11212
rect 18788 11160 18840 11212
rect 19156 11160 19208 11212
rect 19800 11160 19852 11212
rect 19892 11203 19944 11212
rect 19892 11169 19901 11203
rect 19901 11169 19935 11203
rect 19935 11169 19944 11203
rect 19892 11160 19944 11169
rect 8300 11092 8352 11144
rect 9220 11135 9272 11144
rect 9220 11101 9229 11135
rect 9229 11101 9263 11135
rect 9263 11101 9272 11135
rect 9220 11092 9272 11101
rect 11060 11092 11112 11144
rect 11796 11092 11848 11144
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 13728 10956 13780 11008
rect 17868 11024 17920 11076
rect 20352 11067 20404 11076
rect 20352 11033 20361 11067
rect 20361 11033 20395 11067
rect 20395 11033 20404 11067
rect 20352 11024 20404 11033
rect 21364 11067 21416 11076
rect 21364 11033 21373 11067
rect 21373 11033 21407 11067
rect 21407 11033 21416 11067
rect 21364 11024 21416 11033
rect 18052 10956 18104 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 9404 10752 9456 10804
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 13452 10752 13504 10804
rect 15936 10752 15988 10804
rect 16212 10752 16264 10804
rect 19800 10795 19852 10804
rect 8300 10616 8352 10668
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 8944 10548 8996 10600
rect 9588 10548 9640 10600
rect 16488 10684 16540 10736
rect 19800 10761 19809 10795
rect 19809 10761 19843 10795
rect 19843 10761 19852 10795
rect 19800 10752 19852 10761
rect 12900 10616 12952 10668
rect 13176 10616 13228 10668
rect 16672 10548 16724 10600
rect 18052 10616 18104 10668
rect 20076 10616 20128 10668
rect 17868 10548 17920 10600
rect 20536 10548 20588 10600
rect 7656 10480 7708 10532
rect 10692 10480 10744 10532
rect 9404 10455 9456 10464
rect 9404 10421 9413 10455
rect 9413 10421 9447 10455
rect 9447 10421 9456 10455
rect 9404 10412 9456 10421
rect 14648 10480 14700 10532
rect 20444 10480 20496 10532
rect 13084 10412 13136 10464
rect 13452 10412 13504 10464
rect 17960 10412 18012 10464
rect 18972 10455 19024 10464
rect 18972 10421 18981 10455
rect 18981 10421 19015 10455
rect 19015 10421 19024 10455
rect 18972 10412 19024 10421
rect 20260 10455 20312 10464
rect 20260 10421 20269 10455
rect 20269 10421 20303 10455
rect 20303 10421 20312 10455
rect 20260 10412 20312 10421
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 9588 10208 9640 10260
rect 13084 10251 13136 10260
rect 13084 10217 13093 10251
rect 13093 10217 13127 10251
rect 13127 10217 13136 10251
rect 13084 10208 13136 10217
rect 13360 10208 13412 10260
rect 14648 10208 14700 10260
rect 18972 10208 19024 10260
rect 20444 10251 20496 10260
rect 20444 10217 20453 10251
rect 20453 10217 20487 10251
rect 20487 10217 20496 10251
rect 20444 10208 20496 10217
rect 20996 10208 21048 10260
rect 9404 10140 9456 10192
rect 11796 10140 11848 10192
rect 13452 10183 13504 10192
rect 13452 10149 13461 10183
rect 13461 10149 13495 10183
rect 13495 10149 13504 10183
rect 13452 10140 13504 10149
rect 14464 10140 14516 10192
rect 16672 10140 16724 10192
rect 17592 10140 17644 10192
rect 8116 10072 8168 10124
rect 12440 10072 12492 10124
rect 13728 10072 13780 10124
rect 13636 10047 13688 10056
rect 13636 10013 13645 10047
rect 13645 10013 13679 10047
rect 13679 10013 13688 10047
rect 13636 10004 13688 10013
rect 13912 10072 13964 10124
rect 18052 10072 18104 10124
rect 19892 10072 19944 10124
rect 20168 10072 20220 10124
rect 9220 9936 9272 9988
rect 15384 9868 15436 9920
rect 20076 9868 20128 9920
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 8944 9664 8996 9716
rect 11796 9707 11848 9716
rect 11796 9673 11805 9707
rect 11805 9673 11839 9707
rect 11839 9673 11848 9707
rect 11796 9664 11848 9673
rect 13912 9707 13964 9716
rect 13912 9673 13921 9707
rect 13921 9673 13955 9707
rect 13955 9673 13964 9707
rect 13912 9664 13964 9673
rect 17868 9664 17920 9716
rect 20260 9664 20312 9716
rect 14372 9596 14424 9648
rect 21088 9596 21140 9648
rect 22008 9639 22060 9648
rect 22008 9605 22017 9639
rect 22017 9605 22051 9639
rect 22051 9605 22060 9639
rect 22008 9596 22060 9605
rect 15384 9571 15436 9580
rect 12900 9503 12952 9512
rect 12900 9469 12918 9503
rect 12918 9469 12952 9503
rect 15384 9537 15393 9571
rect 15393 9537 15427 9571
rect 15427 9537 15436 9571
rect 15384 9528 15436 9537
rect 19892 9528 19944 9580
rect 12900 9460 12952 9469
rect 12440 9392 12492 9444
rect 13636 9460 13688 9512
rect 18052 9460 18104 9512
rect 20996 9503 21048 9512
rect 20996 9469 21005 9503
rect 21005 9469 21039 9503
rect 21039 9469 21048 9503
rect 20996 9460 21048 9469
rect 20076 9392 20128 9444
rect 20352 9392 20404 9444
rect 14464 9367 14516 9376
rect 14464 9333 14473 9367
rect 14473 9333 14507 9367
rect 14507 9333 14516 9367
rect 14464 9324 14516 9333
rect 15752 9324 15804 9376
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 19248 9367 19300 9376
rect 19248 9333 19257 9367
rect 19257 9333 19291 9367
rect 19291 9333 19300 9367
rect 19248 9324 19300 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 11888 9120 11940 9172
rect 12072 9163 12124 9172
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 20168 9120 20220 9172
rect 20996 9120 21048 9172
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 16212 8984 16264 9036
rect 19892 9027 19944 9036
rect 19892 8993 19901 9027
rect 19901 8993 19935 9027
rect 19935 8993 19944 9027
rect 19892 8984 19944 8993
rect 20996 9027 21048 9036
rect 20996 8993 21005 9027
rect 21005 8993 21039 9027
rect 21039 8993 21048 9027
rect 20996 8984 21048 8993
rect 21364 8959 21416 8968
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 17776 8848 17828 8900
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 11888 8576 11940 8628
rect 13268 8619 13320 8628
rect 13268 8585 13277 8619
rect 13277 8585 13311 8619
rect 13311 8585 13320 8619
rect 13268 8576 13320 8585
rect 16212 8619 16264 8628
rect 16212 8585 16221 8619
rect 16221 8585 16255 8619
rect 16255 8585 16264 8619
rect 16212 8576 16264 8585
rect 20996 8576 21048 8628
rect 20536 8551 20588 8560
rect 11244 8415 11296 8424
rect 11244 8381 11253 8415
rect 11253 8381 11287 8415
rect 11287 8381 11296 8415
rect 11244 8372 11296 8381
rect 20536 8517 20545 8551
rect 20545 8517 20579 8551
rect 20579 8517 20588 8551
rect 20536 8508 20588 8517
rect 14648 8440 14700 8492
rect 17132 8372 17184 8424
rect 19892 8415 19944 8424
rect 19892 8381 19901 8415
rect 19901 8381 19935 8415
rect 19935 8381 19944 8415
rect 19892 8372 19944 8381
rect 20444 8372 20496 8424
rect 15200 8304 15252 8356
rect 17408 8304 17460 8356
rect 14740 8236 14792 8288
rect 17500 8279 17552 8288
rect 17500 8245 17509 8279
rect 17509 8245 17543 8279
rect 17543 8245 17552 8279
rect 17500 8236 17552 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 11244 8032 11296 8084
rect 17132 8075 17184 8084
rect 17132 8041 17141 8075
rect 17141 8041 17175 8075
rect 17175 8041 17184 8075
rect 17132 8032 17184 8041
rect 17500 8075 17552 8084
rect 17500 8041 17509 8075
rect 17509 8041 17543 8075
rect 17543 8041 17552 8075
rect 17500 8032 17552 8041
rect 19800 8032 19852 8084
rect 20444 8032 20496 8084
rect 11704 7896 11756 7948
rect 13728 7896 13780 7948
rect 13912 7939 13964 7948
rect 13912 7905 13946 7939
rect 13946 7905 13964 7939
rect 13912 7896 13964 7905
rect 11888 7828 11940 7880
rect 17592 7871 17644 7880
rect 12164 7760 12216 7812
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 18144 7896 18196 7948
rect 19892 7939 19944 7948
rect 19892 7905 19901 7939
rect 19901 7905 19935 7939
rect 19935 7905 19944 7939
rect 19892 7896 19944 7905
rect 18052 7828 18104 7880
rect 14648 7692 14700 7744
rect 15016 7735 15068 7744
rect 15016 7701 15025 7735
rect 15025 7701 15059 7735
rect 15059 7701 15068 7735
rect 15016 7692 15068 7701
rect 16028 7692 16080 7744
rect 21364 7735 21416 7744
rect 21364 7701 21373 7735
rect 21373 7701 21407 7735
rect 21407 7701 21416 7735
rect 21364 7692 21416 7701
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 15568 7488 15620 7540
rect 18144 7488 18196 7540
rect 19892 7488 19944 7540
rect 11704 7352 11756 7404
rect 14740 7395 14792 7404
rect 14740 7361 14749 7395
rect 14749 7361 14783 7395
rect 14783 7361 14792 7395
rect 14740 7352 14792 7361
rect 8208 7284 8260 7336
rect 9956 7259 10008 7268
rect 9956 7225 9990 7259
rect 9990 7225 10008 7259
rect 9956 7216 10008 7225
rect 12164 7259 12216 7268
rect 12164 7225 12176 7259
rect 12176 7225 12216 7259
rect 13728 7284 13780 7336
rect 12164 7216 12216 7225
rect 15016 7216 15068 7268
rect 13912 7148 13964 7200
rect 14556 7148 14608 7200
rect 18236 7216 18288 7268
rect 21364 7191 21416 7200
rect 21364 7157 21373 7191
rect 21373 7157 21407 7191
rect 21407 7157 21416 7191
rect 21364 7148 21416 7157
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 11888 6987 11940 6996
rect 11888 6953 11897 6987
rect 11897 6953 11931 6987
rect 11931 6953 11940 6987
rect 11888 6944 11940 6953
rect 16488 6876 16540 6928
rect 17592 6944 17644 6996
rect 21180 6876 21232 6928
rect 5632 6808 5684 6860
rect 12348 6851 12400 6860
rect 12348 6817 12357 6851
rect 12357 6817 12391 6851
rect 12391 6817 12400 6851
rect 12348 6808 12400 6817
rect 19248 6808 19300 6860
rect 20536 6851 20588 6860
rect 20536 6817 20545 6851
rect 20545 6817 20579 6851
rect 20579 6817 20588 6851
rect 20536 6808 20588 6817
rect 20904 6808 20956 6860
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 14556 6783 14608 6792
rect 9956 6672 10008 6724
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 15200 6715 15252 6724
rect 15200 6681 15209 6715
rect 15209 6681 15243 6715
rect 15243 6681 15252 6715
rect 15200 6672 15252 6681
rect 14280 6604 14332 6656
rect 21364 6647 21416 6656
rect 21364 6613 21373 6647
rect 21373 6613 21407 6647
rect 21407 6613 21416 6647
rect 21364 6604 21416 6613
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 20904 6443 20956 6452
rect 20904 6409 20913 6443
rect 20913 6409 20947 6443
rect 20947 6409 20956 6443
rect 20904 6400 20956 6409
rect 16488 6332 16540 6384
rect 20720 6239 20772 6248
rect 20720 6205 20729 6239
rect 20729 6205 20763 6239
rect 20763 6205 20772 6239
rect 20720 6196 20772 6205
rect 21364 6239 21416 6248
rect 21364 6205 21373 6239
rect 21373 6205 21407 6239
rect 21407 6205 21416 6239
rect 21364 6196 21416 6205
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 5632 5856 5684 5908
rect 12992 5788 13044 5840
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 20996 5763 21048 5772
rect 20996 5729 21005 5763
rect 21005 5729 21039 5763
rect 21039 5729 21048 5763
rect 20996 5720 21048 5729
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 20996 5312 21048 5364
rect 21180 5355 21232 5364
rect 21180 5321 21189 5355
rect 21189 5321 21223 5355
rect 21223 5321 21232 5355
rect 21180 5312 21232 5321
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 20720 5108 20772 5117
rect 21364 5151 21416 5160
rect 21364 5117 21373 5151
rect 21373 5117 21407 5151
rect 21407 5117 21416 5151
rect 21364 5108 21416 5117
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 19984 4768 20036 4820
rect 21364 4743 21416 4752
rect 21364 4709 21373 4743
rect 21373 4709 21407 4743
rect 21407 4709 21416 4743
rect 21364 4700 21416 4709
rect 20996 4675 21048 4684
rect 20996 4641 21005 4675
rect 21005 4641 21039 4675
rect 21039 4641 21048 4675
rect 20996 4632 21048 4641
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 20996 4224 21048 4276
rect 18788 4088 18840 4140
rect 20628 4063 20680 4072
rect 20628 4029 20637 4063
rect 20637 4029 20671 4063
rect 20671 4029 20680 4063
rect 20628 4020 20680 4029
rect 21272 3995 21324 4004
rect 21272 3961 21281 3995
rect 21281 3961 21315 3995
rect 21315 3961 21324 3995
rect 21272 3952 21324 3961
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 17960 3680 18012 3732
rect 16396 3612 16448 3664
rect 20628 3544 20680 3596
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 19432 3340 19484 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 18696 3136 18748 3188
rect 19340 3068 19392 3120
rect 20168 2907 20220 2916
rect 20168 2873 20177 2907
rect 20177 2873 20211 2907
rect 20211 2873 20220 2907
rect 20168 2864 20220 2873
rect 20720 2907 20772 2916
rect 20720 2873 20729 2907
rect 20729 2873 20763 2907
rect 20763 2873 20772 2907
rect 20720 2864 20772 2873
rect 21272 2907 21324 2916
rect 21272 2873 21281 2907
rect 21281 2873 21315 2907
rect 21315 2873 21324 2907
rect 21272 2864 21324 2873
rect 18972 2796 19024 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 18604 2592 18656 2644
rect 17408 2456 17460 2508
rect 19432 2499 19484 2508
rect 19432 2465 19441 2499
rect 19441 2465 19475 2499
rect 19475 2465 19484 2499
rect 19432 2456 19484 2465
rect 21272 2499 21324 2508
rect 21272 2465 21281 2499
rect 21281 2465 21315 2499
rect 21315 2465 21324 2499
rect 21272 2456 21324 2465
rect 14464 2320 14516 2372
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 22008 1411 22060 1420
rect 22008 1377 22017 1411
rect 22017 1377 22051 1411
rect 22051 1377 22060 1411
rect 22008 1368 22060 1377
<< metal2 >>
rect 294 22200 350 23000
rect 846 22200 902 23000
rect 1398 22200 1454 23000
rect 1950 22200 2006 23000
rect 2502 22200 2558 23000
rect 3054 22200 3110 23000
rect 3606 22200 3662 23000
rect 4158 22200 4214 23000
rect 4710 22200 4766 23000
rect 5262 22200 5318 23000
rect 5814 22200 5870 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 12070 22200 12126 23000
rect 12622 22200 12678 23000
rect 13174 22200 13230 23000
rect 13726 22200 13782 23000
rect 14278 22200 14334 23000
rect 14830 22200 14886 23000
rect 15382 22200 15438 23000
rect 15934 22200 15990 23000
rect 16486 22200 16542 23000
rect 17038 22200 17094 23000
rect 17682 22200 17738 23000
rect 17958 22264 18014 22273
rect 308 20398 336 22200
rect 860 20466 888 22200
rect 1412 20534 1440 22200
rect 1400 20528 1452 20534
rect 1400 20470 1452 20476
rect 848 20460 900 20466
rect 848 20402 900 20408
rect 296 20392 348 20398
rect 296 20334 348 20340
rect 1308 20392 1360 20398
rect 1308 20334 1360 20340
rect 1320 20058 1348 20334
rect 1964 20330 1992 22200
rect 2516 20482 2544 22200
rect 3068 20874 3096 22200
rect 3056 20868 3108 20874
rect 3056 20810 3108 20816
rect 3620 20618 3648 22200
rect 4172 20806 4200 22200
rect 4724 20890 4752 22200
rect 4724 20874 4844 20890
rect 4252 20868 4304 20874
rect 4252 20810 4304 20816
rect 4712 20868 4844 20874
rect 4764 20862 4844 20868
rect 4712 20810 4764 20816
rect 4160 20800 4212 20806
rect 4160 20742 4212 20748
rect 3620 20590 4200 20618
rect 3608 20528 3660 20534
rect 2516 20466 2820 20482
rect 3608 20470 3660 20476
rect 2516 20460 2832 20466
rect 2516 20454 2780 20460
rect 2780 20402 2832 20408
rect 2044 20392 2096 20398
rect 2044 20334 2096 20340
rect 2504 20392 2556 20398
rect 2504 20334 2556 20340
rect 1952 20324 2004 20330
rect 1952 20266 2004 20272
rect 1768 20256 1820 20262
rect 1768 20198 1820 20204
rect 1308 20052 1360 20058
rect 1308 19994 1360 20000
rect 1780 19922 1808 20198
rect 2056 20058 2084 20334
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2044 20052 2096 20058
rect 2044 19994 2096 20000
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1768 18828 1820 18834
rect 1768 18770 1820 18776
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1688 17241 1716 17478
rect 1780 17338 1808 18770
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1674 17232 1730 17241
rect 1674 17167 1730 17176
rect 1780 16590 1808 17274
rect 1768 16584 1820 16590
rect 1768 16526 1820 16532
rect 2332 11694 2360 20198
rect 2516 20058 2544 20334
rect 2872 20324 2924 20330
rect 2872 20266 2924 20272
rect 2884 20058 2912 20266
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 3620 17882 3648 20470
rect 4172 20466 4200 20590
rect 3792 20460 3844 20466
rect 3792 20402 3844 20408
rect 4160 20460 4212 20466
rect 4160 20402 4212 20408
rect 3804 20058 3832 20402
rect 4264 20398 4292 20810
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 3896 18630 3924 19246
rect 4264 19242 4292 19790
rect 4632 19786 4660 20198
rect 4816 20074 4844 20862
rect 5172 20528 5224 20534
rect 5172 20470 5224 20476
rect 5080 20392 5132 20398
rect 5080 20334 5132 20340
rect 4896 20256 4948 20262
rect 4948 20216 5028 20244
rect 4896 20198 4948 20204
rect 4724 20046 4844 20074
rect 4724 19990 4752 20046
rect 4712 19984 4764 19990
rect 4712 19926 4764 19932
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4816 19310 4844 19858
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 4264 18970 4292 19178
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4816 18766 4844 19110
rect 4908 18970 4936 19654
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 3608 17876 3660 17882
rect 3608 17818 3660 17824
rect 3700 17672 3752 17678
rect 3700 17614 3752 17620
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 2884 15706 2912 17002
rect 3068 16794 3096 17478
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3528 16794 3556 17274
rect 3712 17066 3740 17614
rect 3896 17134 3924 18566
rect 4264 17134 4292 18566
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 3700 17060 3752 17066
rect 3700 17002 3752 17008
rect 3056 16788 3108 16794
rect 3056 16730 3108 16736
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3896 16658 3924 17070
rect 4816 16726 4844 18702
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 3896 15638 3924 16594
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 3884 15632 3936 15638
rect 3884 15574 3936 15580
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2516 15026 2544 15506
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2516 14618 2544 14962
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 3896 14414 3924 15574
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4816 15162 4844 15370
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4264 14618 4292 14758
rect 5000 14618 5028 20216
rect 5092 19990 5120 20334
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 5184 19854 5212 20470
rect 5276 19922 5304 22200
rect 5448 20868 5500 20874
rect 5448 20810 5500 20816
rect 5460 20466 5488 20810
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5552 20398 5580 20742
rect 5356 20392 5408 20398
rect 5356 20334 5408 20340
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5368 19990 5396 20334
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5460 20058 5488 20198
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5552 18970 5580 20334
rect 5828 19990 5856 22200
rect 6472 20398 6500 22200
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6748 20505 6776 20538
rect 6932 20505 6960 20538
rect 6734 20496 6790 20505
rect 6918 20496 6974 20505
rect 6734 20431 6790 20440
rect 6828 20460 6880 20466
rect 6918 20431 6974 20440
rect 6828 20402 6880 20408
rect 6460 20392 6512 20398
rect 6460 20334 6512 20340
rect 6092 20256 6144 20262
rect 6092 20198 6144 20204
rect 5816 19984 5868 19990
rect 5816 19926 5868 19932
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5276 16658 5304 18158
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5552 17678 5580 18090
rect 5736 17882 5764 19858
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5920 18222 5948 19246
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5552 16250 5580 17614
rect 6104 17134 6132 20198
rect 6472 19990 6500 20334
rect 6840 20058 6868 20402
rect 6920 20392 6972 20398
rect 7024 20380 7052 22200
rect 7576 20398 7604 22200
rect 8128 20618 8156 22200
rect 8128 20590 8340 20618
rect 7748 20528 7800 20534
rect 7748 20470 7800 20476
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 7104 20392 7156 20398
rect 7024 20352 7104 20380
rect 6920 20334 6972 20340
rect 7104 20334 7156 20340
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6460 19984 6512 19990
rect 6460 19926 6512 19932
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6656 18426 6684 19178
rect 6748 18902 6776 19858
rect 6932 19378 6960 20334
rect 7116 19514 7144 20334
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7208 19310 7236 19790
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 6736 18896 6788 18902
rect 6736 18838 6788 18844
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7208 18426 7236 18770
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7300 18222 7328 18702
rect 7484 18408 7512 20198
rect 7576 18970 7604 20334
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7484 18380 7604 18408
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 7392 17882 7420 18022
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 7484 16726 7512 17138
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 7300 16114 7328 16594
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6104 15502 6132 15914
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6104 15162 6132 15438
rect 7300 15366 7328 16050
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 7484 14958 7512 15982
rect 7576 15094 7604 18380
rect 7668 17678 7696 20198
rect 7760 19514 7788 20470
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7852 19446 7880 19858
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7760 17542 7788 17682
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7760 16574 7788 17478
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7668 16546 7788 16574
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 4172 14074 4200 14418
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 7208 13530 7236 14826
rect 7484 13870 7512 14894
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 2320 11688 2372 11694
rect 2320 11630 2372 11636
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 7668 10538 7696 16546
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7760 15162 7788 15438
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 8220 15026 8248 20470
rect 8312 20398 8340 20590
rect 8680 20398 8708 22200
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8312 20058 8340 20334
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8496 17202 8524 17682
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 8312 16794 8340 16934
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 8312 14550 8340 14758
rect 8588 14618 8616 19654
rect 8680 19378 8708 20198
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8496 13802 8524 14350
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 8220 13326 8248 13738
rect 8680 13326 8708 14010
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8220 12102 8248 13262
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11694 8248 12038
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7656 10532 7708 10538
rect 7656 10474 7708 10480
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 8116 10124 8168 10130
rect 8220 10112 8248 11630
rect 8864 11286 8892 20538
rect 9232 20398 9260 22200
rect 9784 20398 9812 22200
rect 10336 20398 10364 22200
rect 10888 20398 10916 22200
rect 11440 20890 11468 22200
rect 11440 20862 11744 20890
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 9220 20392 9272 20398
rect 9220 20334 9272 20340
rect 9772 20392 9824 20398
rect 9772 20334 9824 20340
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10876 20392 10928 20398
rect 10928 20352 11008 20380
rect 10876 20334 10928 20340
rect 9140 19786 9168 20334
rect 9232 19922 9260 20334
rect 9588 20256 9640 20262
rect 9588 20198 9640 20204
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8956 19378 8984 19654
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 8944 19236 8996 19242
rect 8944 19178 8996 19184
rect 8956 18630 8984 19178
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8956 18426 8984 18566
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 9416 18222 9444 19314
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9600 17882 9628 20198
rect 9784 19990 9812 20334
rect 10336 20058 10364 20334
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10324 20052 10376 20058
rect 10324 19994 10376 20000
rect 10888 19990 10916 20198
rect 9772 19984 9824 19990
rect 9772 19926 9824 19932
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 10980 19854 11008 20352
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 9692 19310 9720 19790
rect 11256 19786 11284 20266
rect 11716 19922 11744 20862
rect 12084 20534 12112 22200
rect 12636 20534 12664 22200
rect 13188 20534 13216 22200
rect 13740 20534 13768 22200
rect 14292 20602 14320 22200
rect 14844 20754 14872 22200
rect 14844 20726 15148 20754
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 12072 20528 12124 20534
rect 12072 20470 12124 20476
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 13176 20528 13228 20534
rect 13176 20470 13228 20476
rect 13728 20528 13780 20534
rect 13728 20470 13780 20476
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 10876 19304 10928 19310
rect 10928 19264 11008 19292
rect 10876 19246 10928 19252
rect 10232 18828 10284 18834
rect 10232 18770 10284 18776
rect 10244 18086 10272 18770
rect 10980 18630 11008 19264
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 10980 18154 11008 18566
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9140 16574 9168 17682
rect 9784 17678 9812 18022
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 8956 16546 9168 16574
rect 9404 16584 9456 16590
rect 8956 12170 8984 16546
rect 9404 16526 9456 16532
rect 9416 16046 9444 16526
rect 10980 16114 11008 18090
rect 11164 17134 11192 19654
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11336 19236 11388 19242
rect 11336 19178 11388 19184
rect 11348 18970 11376 19178
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11348 18714 11376 18906
rect 11808 18834 11836 20470
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 11888 20324 11940 20330
rect 11888 20266 11940 20272
rect 12164 20324 12216 20330
rect 12164 20266 12216 20272
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11256 18686 11376 18714
rect 11256 18290 11284 18686
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 11244 18080 11296 18086
rect 11244 18022 11296 18028
rect 11256 17882 11284 18022
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 11256 16250 11284 17138
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 10980 15638 11008 16050
rect 11256 16046 11284 16186
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 10968 15632 11020 15638
rect 10968 15574 11020 15580
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9140 14822 9168 15302
rect 9324 14822 9352 15506
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 13530 9076 14214
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9324 12306 9352 14758
rect 9600 14482 9628 15302
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 9496 14476 9548 14482
rect 9496 14418 9548 14424
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9508 13530 9536 14418
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9600 13190 9628 13738
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12850 9628 13126
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 8944 12164 8996 12170
rect 8944 12106 8996 12112
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8312 10674 8340 11086
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8956 10606 8984 12106
rect 9220 11620 9272 11626
rect 9220 11562 9272 11568
rect 9232 11150 9260 11562
rect 9692 11286 9720 14350
rect 11072 14074 11100 14894
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9784 12986 9812 13330
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10704 12442 10732 12582
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11354 9812 11494
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8168 10084 8248 10112
rect 8116 10066 8168 10072
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 8220 7342 8248 10084
rect 8956 9722 8984 10542
rect 9232 9994 9260 11086
rect 9416 10810 9444 11154
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 10198 9444 10406
rect 9600 10266 9628 10542
rect 10704 10538 10732 12378
rect 11072 11762 11100 12650
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11164 12442 11192 12582
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11716 11898 11744 12242
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11348 11354 11376 11494
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10796 10674 10824 11154
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11072 10810 11100 11086
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 11808 10198 11836 11086
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11808 9722 11836 10134
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11900 9178 11928 20266
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11992 18970 12020 19110
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 12084 18766 12112 19110
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12176 18442 12204 20266
rect 12084 18414 12204 18442
rect 12084 9178 12112 18414
rect 12268 14618 12296 20402
rect 12900 20324 12952 20330
rect 12900 20266 12952 20272
rect 13268 20324 13320 20330
rect 15120 20312 15148 20726
rect 15120 20284 15240 20312
rect 13268 20266 13320 20272
rect 12912 19718 12940 20266
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12348 19508 12400 19514
rect 12348 19450 12400 19456
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12176 13938 12204 14350
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12176 13326 12204 13874
rect 12268 13394 12296 14282
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12176 12986 12204 13262
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11900 8634 11928 8978
rect 11888 8628 11940 8634
rect 11888 8570 11940 8576
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11256 8090 11284 8366
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11716 7410 11744 7890
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 5644 5914 5672 6802
rect 8220 6798 8248 7278
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 9968 6730 9996 7210
rect 11900 7002 11928 7822
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12176 7274 12204 7754
rect 12164 7268 12216 7274
rect 12164 7210 12216 7216
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 12360 6866 12388 19450
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12452 18086 12480 18770
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 17610 12480 18022
rect 12440 17604 12492 17610
rect 12440 17546 12492 17552
rect 12452 17066 12480 17546
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12452 13394 12480 17002
rect 12544 16658 12572 17138
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12636 16794 12664 16934
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12544 16250 12572 16594
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12728 14906 12756 18294
rect 12544 14878 12756 14906
rect 12544 13530 12572 14878
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12636 14618 12664 14758
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12728 13530 12756 14758
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12544 13308 12572 13466
rect 12820 13394 12848 14010
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12716 13320 12768 13326
rect 12544 13280 12716 13308
rect 12716 13262 12768 13268
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12306 12480 12718
rect 12912 12434 12940 19654
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 13188 18834 13216 19246
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 13096 18222 13124 18702
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13096 14618 13124 14758
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13188 13734 13216 14758
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 12912 12406 13032 12434
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12452 10130 12480 12242
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 12440 10124 12492 10130
rect 12440 10066 12492 10072
rect 12452 9450 12480 10066
rect 12912 9518 12940 10610
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 12440 9444 12492 9450
rect 12440 9386 12492 9392
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 13004 5846 13032 12406
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 13096 11762 13124 12038
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13188 10674 13216 11494
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13096 10266 13124 10406
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13280 8634 13308 20266
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14372 20256 14424 20262
rect 14372 20198 14424 20204
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18902 13860 19110
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13372 18290 13400 18566
rect 13832 18358 13860 18838
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13360 18284 13412 18290
rect 13360 18226 13412 18232
rect 14200 18154 14228 20198
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14188 18148 14240 18154
rect 14188 18090 14240 18096
rect 14292 16794 14320 19450
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14292 15978 14320 16526
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14016 14482 14044 14962
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13372 12434 13400 14214
rect 14016 14074 14044 14418
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13372 12406 13492 12434
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13372 10282 13400 11834
rect 13464 11558 13492 12406
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13464 10810 13492 11086
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 10282 13492 10406
rect 13372 10266 13492 10282
rect 13360 10260 13492 10266
rect 13412 10254 13492 10260
rect 13360 10202 13412 10208
rect 13452 10192 13504 10198
rect 13556 10146 13584 13126
rect 13648 11898 13676 13262
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13504 10140 13584 10146
rect 13452 10134 13584 10140
rect 13464 10118 13584 10134
rect 13648 10062 13676 11698
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13740 11014 13768 11562
rect 13924 11354 13952 12718
rect 14384 12434 14412 20198
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15212 19990 15240 20284
rect 15396 19990 15424 22200
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15200 19984 15252 19990
rect 15200 19926 15252 19932
rect 15384 19984 15436 19990
rect 15384 19926 15436 19932
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 15568 19916 15620 19922
rect 15568 19858 15620 19864
rect 14556 19304 14608 19310
rect 14556 19246 14608 19252
rect 14568 18290 14596 19246
rect 14660 18630 14688 19858
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14844 19310 14872 19790
rect 14832 19304 14884 19310
rect 14752 19252 14832 19258
rect 14752 19246 14884 19252
rect 14752 19230 14872 19246
rect 14752 18970 14780 19230
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 14740 18964 14792 18970
rect 14740 18906 14792 18912
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14568 16590 14596 18226
rect 14660 16658 14688 18566
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15212 17082 15240 17138
rect 15212 17054 15332 17082
rect 14740 16992 14792 16998
rect 14740 16934 14792 16940
rect 14752 16794 14780 16934
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 15304 16658 15332 17054
rect 14648 16652 14700 16658
rect 14648 16594 14700 16600
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14568 16454 14596 16526
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14568 16114 14596 16390
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14568 15502 14596 16050
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 15162 14596 15438
rect 14660 15366 14688 16594
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 14648 15360 14700 15366
rect 14648 15302 14700 15308
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14568 13530 14596 14894
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14292 12406 14412 12434
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13740 10130 13768 10950
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13648 9518 13676 9998
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13740 7954 13768 10066
rect 13924 9722 13952 10066
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13740 7342 13768 7890
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13924 7206 13952 7890
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 14292 6662 14320 12406
rect 14568 11218 14596 13466
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14384 9654 14412 11154
rect 14660 10538 14688 15302
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14752 14498 14780 15098
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14752 14482 14964 14498
rect 14752 14476 14976 14482
rect 14752 14470 14924 14476
rect 14752 13870 14780 14470
rect 14924 14418 14976 14424
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 15212 13530 15240 13670
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15292 12912 15344 12918
rect 15292 12854 15344 12860
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15212 12442 15240 12650
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15304 12374 15332 12854
rect 15292 12368 15344 12374
rect 15292 12310 15344 12316
rect 15304 11898 15332 12310
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14660 10266 14688 10474
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 14648 10260 14700 10266
rect 14648 10202 14700 10208
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14476 9382 14504 10134
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 9586 15424 9862
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 12992 5840 13044 5846
rect 1582 5808 1638 5817
rect 12992 5782 13044 5788
rect 1582 5743 1584 5752
rect 1636 5743 1638 5752
rect 1584 5714 1636 5720
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 14476 2378 14504 9318
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14660 7750 14688 8434
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14752 7410 14780 8230
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 15028 7274 15056 7686
rect 15016 7268 15068 7274
rect 15016 7210 15068 7216
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 6798 14596 7142
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 15212 6730 15240 8298
rect 15580 7546 15608 19858
rect 15856 19446 15884 20334
rect 15948 19990 15976 22200
rect 16212 20392 16264 20398
rect 16212 20334 16264 20340
rect 15936 19984 15988 19990
rect 15936 19926 15988 19932
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15844 19440 15896 19446
rect 15844 19382 15896 19388
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18222 15884 19110
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15948 16250 15976 16594
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15660 14476 15712 14482
rect 15660 14418 15712 14424
rect 15672 14074 15700 14418
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15764 9382 15792 13466
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15948 12442 15976 12582
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15948 11694 15976 12174
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15948 10810 15976 11630
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 16040 7750 16068 19858
rect 16120 16040 16172 16046
rect 16120 15982 16172 15988
rect 16132 15706 16160 15982
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16224 10810 16252 20334
rect 16500 20074 16528 22200
rect 16500 20058 16620 20074
rect 16304 20052 16356 20058
rect 16500 20052 16632 20058
rect 16500 20046 16580 20052
rect 16304 19994 16356 20000
rect 16580 19994 16632 20000
rect 16316 13682 16344 19994
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16592 19310 16620 19790
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16684 19378 16712 19722
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 17746 16528 18022
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16592 16114 16620 16390
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16592 15570 16620 16050
rect 16684 15910 16712 16186
rect 16776 15978 16804 19654
rect 17052 19310 17080 22200
rect 17696 20534 17724 22200
rect 17958 22199 18014 22208
rect 18234 22200 18290 23000
rect 18786 22200 18842 23000
rect 19338 22200 19394 23000
rect 19706 22672 19762 22681
rect 19706 22607 19762 22616
rect 17972 20534 18000 22199
rect 18248 20890 18276 22200
rect 18602 21720 18658 21729
rect 18602 21655 18658 21664
rect 18156 20862 18276 20890
rect 18156 20602 18184 20862
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18616 20534 18644 21655
rect 18800 20534 18828 22200
rect 18970 21312 19026 21321
rect 18970 21247 19026 21256
rect 18984 20534 19012 21247
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 17960 20528 18012 20534
rect 17960 20470 18012 20476
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 17592 20324 17644 20330
rect 17592 20266 17644 20272
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 18604 20324 18656 20330
rect 18604 20266 18656 20272
rect 18880 20324 18932 20330
rect 18880 20266 18932 20272
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 16960 18834 16988 19110
rect 17052 18970 17080 19110
rect 17040 18964 17092 18970
rect 17040 18906 17092 18912
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 17328 18630 17356 19178
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17328 17814 17356 18226
rect 17316 17808 17368 17814
rect 17316 17750 17368 17756
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 13870 16436 14214
rect 16684 13920 16712 15846
rect 17144 15502 17172 17614
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 17144 15026 17172 15438
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17144 13938 17172 14962
rect 16500 13892 16712 13920
rect 17132 13932 17184 13938
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16316 13654 16436 13682
rect 16304 13184 16356 13190
rect 16304 13126 16356 13132
rect 16316 12782 16344 13126
rect 16408 12850 16436 13654
rect 16500 13530 16528 13892
rect 17132 13874 17184 13880
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16316 11286 16344 12718
rect 17144 12714 17172 12786
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 16592 12442 16620 12650
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 17328 11898 17356 12786
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16500 10742 16528 11154
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16684 10198 16712 10542
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16224 8634 16252 8978
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 16408 3670 16436 9318
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 17144 8090 17172 8366
rect 17420 8362 17448 19858
rect 17604 19718 17632 20266
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17512 18970 17540 19246
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17604 17814 17632 18022
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17604 16250 17632 17750
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17512 12646 17540 12786
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17696 12238 17724 12718
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17604 10198 17632 12174
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17408 8356 17460 8362
rect 17408 8298 17460 8304
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17512 8090 17540 8230
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17604 7970 17632 10134
rect 17788 8906 17816 19858
rect 18156 18970 18184 20266
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18616 19514 18644 20266
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 18064 18426 18092 18770
rect 18604 18760 18656 18766
rect 18604 18702 18656 18708
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18340 17882 18368 18226
rect 18616 18222 18644 18702
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18156 17338 18184 17614
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 18708 16810 18736 19790
rect 18616 16782 18736 16810
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17972 15706 18000 16050
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 17972 14890 18000 15642
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 17868 14884 17920 14890
rect 17868 14826 17920 14832
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17880 14618 17908 14826
rect 18616 14822 18644 16782
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18708 16250 18736 16594
rect 18892 16402 18920 20266
rect 19352 20058 19380 22200
rect 19522 20904 19578 20913
rect 19522 20839 19578 20848
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19444 20262 19472 20538
rect 19536 20534 19564 20839
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19076 18834 19104 19246
rect 19536 18970 19564 20334
rect 19720 19990 19748 22607
rect 19890 22200 19946 23000
rect 20442 22200 20498 23000
rect 20994 22200 21050 23000
rect 21546 22200 21602 23000
rect 22098 22200 22154 23000
rect 22650 22200 22706 23000
rect 19708 19984 19760 19990
rect 19708 19926 19760 19932
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 19076 17134 19104 18022
rect 19260 17338 19288 18770
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 19352 16794 19380 18226
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19444 16794 19472 16934
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 18800 16374 18920 16402
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 18604 14476 18656 14482
rect 18604 14418 18656 14424
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 18064 13870 18092 14282
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 13326 18092 13806
rect 18616 13802 18644 14418
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18616 13190 18644 13738
rect 18708 13734 18736 14350
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18708 13462 18736 13670
rect 18696 13456 18748 13462
rect 18696 13398 18748 13404
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17880 11082 17908 12174
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 11354 18092 11494
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17880 10606 17908 11018
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 10674 18092 10950
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17880 9722 17908 10542
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 17420 7942 17632 7970
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16500 6390 16528 6870
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 16396 3664 16448 3670
rect 16396 3606 16448 3612
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 17420 2514 17448 7942
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7002 17632 7822
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17972 3738 18000 10406
rect 18064 10130 18092 10610
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18064 9518 18092 10066
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 7886 18092 9454
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 18156 7546 18184 7890
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18236 7268 18288 7274
rect 18236 7210 18288 7216
rect 18248 6798 18276 7210
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 2650 18644 13126
rect 18800 11898 18828 16374
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19168 14346 19196 14758
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18892 13530 18920 13806
rect 19352 13530 19380 14418
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18984 12374 19012 12582
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 18708 3194 18736 11630
rect 19076 11354 19104 11630
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 18800 4146 18828 11154
rect 18984 10470 19012 11222
rect 19168 11218 19196 13466
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19260 12073 19288 12242
rect 19628 12102 19656 19858
rect 19720 18986 19748 19926
rect 19904 19854 19932 22200
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 20180 19446 20208 20266
rect 20168 19440 20220 19446
rect 20168 19382 20220 19388
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19720 18958 19840 18986
rect 19708 18828 19760 18834
rect 19708 18770 19760 18776
rect 19720 17882 19748 18770
rect 19812 18426 19840 18958
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19708 17876 19760 17882
rect 19708 17818 19760 17824
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19720 16658 19748 17138
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19812 12866 19840 18022
rect 19904 13002 19932 19314
rect 20076 19304 20128 19310
rect 20076 19246 20128 19252
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19996 18086 20024 18770
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 20088 13258 20116 19246
rect 20272 18698 20300 20334
rect 20352 19984 20404 19990
rect 20352 19926 20404 19932
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 20180 16250 20208 18158
rect 20260 18148 20312 18154
rect 20260 18090 20312 18096
rect 20272 17882 20300 18090
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20272 16046 20300 16390
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20364 15858 20392 19926
rect 20456 19310 20484 22200
rect 21008 20602 21036 22200
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20810 20360 20866 20369
rect 20548 19514 20576 20334
rect 20810 20295 20812 20304
rect 20864 20295 20866 20304
rect 21364 20324 21416 20330
rect 20812 20266 20864 20272
rect 21364 20266 21416 20272
rect 21376 19961 21404 20266
rect 21362 19952 21418 19961
rect 20628 19916 20680 19922
rect 21362 19887 21418 19896
rect 20628 19858 20680 19864
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20444 19304 20496 19310
rect 20444 19246 20496 19252
rect 20536 19236 20588 19242
rect 20536 19178 20588 19184
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20272 15830 20392 15858
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20180 14550 20208 14894
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 20076 13252 20128 13258
rect 20076 13194 20128 13200
rect 19904 12974 20208 13002
rect 19812 12838 19932 12866
rect 19800 12776 19852 12782
rect 19800 12718 19852 12724
rect 19812 12617 19840 12718
rect 19798 12608 19854 12617
rect 19798 12543 19854 12552
rect 19904 12434 19932 12838
rect 20180 12442 20208 12974
rect 20168 12436 20220 12442
rect 19904 12406 20024 12434
rect 19340 12096 19392 12102
rect 19246 12064 19302 12073
rect 19340 12038 19392 12044
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19246 11999 19302 12008
rect 19156 11212 19208 11218
rect 19156 11154 19208 11160
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18984 10266 19012 10406
rect 18972 10260 19024 10266
rect 18972 10202 19024 10208
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18984 2854 19012 10202
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19260 6866 19288 9318
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19352 3126 19380 12038
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19812 10810 19840 11154
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19904 10713 19932 11154
rect 19890 10704 19946 10713
rect 19890 10639 19946 10648
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19904 9586 19932 10066
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19904 9466 19932 9522
rect 19812 9438 19932 9466
rect 19812 8090 19840 9438
rect 19890 9344 19946 9353
rect 19890 9279 19946 9288
rect 19904 9042 19932 9279
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 19892 8424 19944 8430
rect 19890 8392 19892 8401
rect 19944 8392 19946 8401
rect 19890 8327 19946 8336
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19890 7984 19946 7993
rect 19890 7919 19892 7928
rect 19944 7919 19946 7928
rect 19892 7890 19944 7896
rect 19904 7546 19932 7890
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19996 4826 20024 12406
rect 20168 12378 20220 12384
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20088 11898 20116 12174
rect 20272 11898 20300 15830
rect 20352 15632 20404 15638
rect 20352 15574 20404 15580
rect 20364 15162 20392 15574
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20456 15042 20484 18770
rect 20548 15858 20576 19178
rect 20640 18426 20668 19858
rect 21364 19780 21416 19786
rect 21364 19722 21416 19728
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 20904 19236 20956 19242
rect 20904 19178 20956 19184
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20640 17338 20668 17682
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20732 16794 20760 17682
rect 20810 17640 20866 17649
rect 20810 17575 20812 17584
rect 20864 17575 20866 17584
rect 20812 17546 20864 17552
rect 20720 16788 20772 16794
rect 20720 16730 20772 16736
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 20548 15830 20668 15858
rect 20364 15014 20484 15042
rect 20364 13530 20392 15014
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20364 12986 20392 13262
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20456 12918 20484 14350
rect 20548 14074 20576 14894
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20640 13818 20668 15830
rect 20824 15706 20852 15914
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20916 14618 20944 19178
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20548 13025 20576 13806
rect 20640 13790 20760 13818
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20640 13394 20668 13670
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20732 13274 20760 13790
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20640 13246 20760 13274
rect 20534 13016 20590 13025
rect 20534 12951 20590 12960
rect 20444 12912 20496 12918
rect 20444 12854 20496 12860
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 12170 20484 12718
rect 20640 12442 20668 13246
rect 20916 12986 20944 13330
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20640 11354 20668 12038
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20088 9926 20116 10610
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20168 10124 20220 10130
rect 20168 10066 20220 10072
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 20088 9450 20116 9862
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 20180 9178 20208 10066
rect 20272 9722 20300 10406
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 20364 9450 20392 11018
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20456 10266 20484 10474
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20548 8566 20576 10542
rect 21008 10266 21036 19654
rect 21376 19417 21404 19722
rect 21362 19408 21418 19417
rect 21362 19343 21418 19352
rect 21364 19236 21416 19242
rect 21364 19178 21416 19184
rect 21376 19009 21404 19178
rect 21560 19174 21588 22200
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21362 19000 21418 19009
rect 21362 18935 21418 18944
rect 22112 18902 22140 22200
rect 22664 18970 22692 22200
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 22100 18896 22152 18902
rect 22100 18838 22152 18844
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 21100 9654 21128 18566
rect 21192 18426 21220 18770
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21376 18601 21404 18634
rect 21362 18592 21418 18601
rect 21362 18527 21418 18536
rect 21180 18420 21232 18426
rect 21180 18362 21232 18368
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21376 18057 21404 18090
rect 21362 18048 21418 18057
rect 21362 17983 21418 17992
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21376 17241 21404 17546
rect 21362 17232 21418 17241
rect 21362 17167 21418 17176
rect 21180 17060 21232 17066
rect 21180 17002 21232 17008
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21192 16794 21220 17002
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21468 16697 21496 17002
rect 21454 16688 21510 16697
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21364 16652 21416 16658
rect 21454 16623 21510 16632
rect 21364 16594 21416 16600
rect 21192 16250 21220 16594
rect 21376 16289 21404 16594
rect 21362 16280 21418 16289
rect 21180 16244 21232 16250
rect 21362 16215 21418 16224
rect 21180 16186 21232 16192
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21376 15745 21404 15914
rect 21362 15736 21418 15745
rect 21362 15671 21418 15680
rect 21364 15428 21416 15434
rect 21364 15370 21416 15376
rect 21376 15337 21404 15370
rect 21362 15328 21418 15337
rect 21362 15263 21418 15272
rect 21362 14920 21418 14929
rect 21362 14855 21364 14864
rect 21416 14855 21418 14864
rect 21364 14826 21416 14832
rect 21270 14376 21326 14385
rect 21270 14311 21272 14320
rect 21324 14311 21326 14320
rect 21272 14282 21324 14288
rect 21362 13968 21418 13977
rect 21362 13903 21364 13912
rect 21416 13903 21418 13912
rect 21364 13874 21416 13880
rect 21180 13796 21232 13802
rect 21180 13738 21232 13744
rect 21192 12986 21220 13738
rect 21362 13560 21418 13569
rect 21362 13495 21418 13504
rect 21376 13462 21404 13495
rect 21364 13456 21416 13462
rect 21364 13398 21416 13404
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21376 11694 21404 12038
rect 21364 11688 21416 11694
rect 21362 11656 21364 11665
rect 21416 11656 21418 11665
rect 21362 11591 21418 11600
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 11257 21404 11494
rect 21362 11248 21418 11257
rect 21362 11183 21418 11192
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21376 10305 21404 11018
rect 21362 10296 21418 10305
rect 21362 10231 21418 10240
rect 22006 9752 22062 9761
rect 22006 9687 22062 9696
rect 22020 9654 22048 9687
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 22008 9648 22060 9654
rect 22008 9590 22060 9596
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 21008 9178 21036 9454
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 21008 8634 21036 8978
rect 21364 8968 21416 8974
rect 21362 8936 21364 8945
rect 21416 8936 21418 8945
rect 21362 8871 21418 8880
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20536 8560 20588 8566
rect 20536 8502 20588 8508
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20456 8090 20484 8366
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21376 7585 21404 7686
rect 21362 7576 21418 7585
rect 21362 7511 21418 7520
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21376 7041 21404 7142
rect 21362 7032 21418 7041
rect 21362 6967 21418 6976
rect 21180 6928 21232 6934
rect 21180 6870 21232 6876
rect 20536 6860 20588 6866
rect 20536 6802 20588 6808
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20548 6633 20576 6802
rect 20534 6624 20590 6633
rect 20534 6559 20590 6568
rect 20916 6458 20944 6802
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20732 6089 20760 6190
rect 20718 6080 20774 6089
rect 20718 6015 20774 6024
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 21008 5370 21036 5714
rect 21192 5370 21220 6870
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 21376 6254 21404 6598
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21376 5681 21404 6190
rect 21362 5672 21418 5681
rect 21362 5607 21418 5616
rect 20996 5364 21048 5370
rect 20996 5306 21048 5312
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 20718 5264 20774 5273
rect 20718 5199 20774 5208
rect 20732 5166 20760 5199
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 21376 4758 21404 5102
rect 21364 4752 21416 4758
rect 21362 4720 21364 4729
rect 21416 4720 21418 4729
rect 20996 4684 21048 4690
rect 21362 4655 21418 4664
rect 20996 4626 21048 4632
rect 20626 4312 20682 4321
rect 21008 4282 21036 4626
rect 20626 4247 20682 4256
rect 20996 4276 21048 4282
rect 20640 4078 20668 4247
rect 20996 4218 21048 4224
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 21272 4004 21324 4010
rect 21272 3946 21324 3952
rect 21284 3913 21312 3946
rect 21270 3904 21326 3913
rect 21270 3839 21326 3848
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 19444 2514 19472 3334
rect 20168 2916 20220 2922
rect 20168 2858 20220 2864
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 19432 2508 19484 2514
rect 19432 2450 19484 2456
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 19444 1057 19472 2450
rect 20180 2009 20208 2858
rect 20166 2000 20222 2009
rect 20166 1935 20222 1944
rect 20640 1601 20668 3538
rect 21284 3369 21312 3538
rect 21270 3360 21326 3369
rect 21270 3295 21326 3304
rect 21270 2952 21326 2961
rect 20720 2916 20772 2922
rect 21270 2887 21272 2896
rect 20720 2858 20772 2864
rect 21324 2887 21326 2896
rect 21272 2858 21324 2864
rect 20626 1592 20682 1601
rect 20626 1527 20682 1536
rect 19430 1048 19486 1057
rect 19430 983 19486 992
rect 20732 649 20760 2858
rect 21272 2508 21324 2514
rect 21272 2450 21324 2456
rect 21284 2417 21312 2450
rect 21270 2408 21326 2417
rect 21270 2343 21326 2352
rect 22008 1420 22060 1426
rect 22008 1362 22060 1368
rect 20718 640 20774 649
rect 20718 575 20774 584
rect 22020 241 22048 1362
rect 22006 232 22062 241
rect 22006 167 22062 176
<< via2 >>
rect 17958 22208 18014 22264
rect 1674 17176 1730 17232
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 6734 20440 6790 20496
rect 6918 20440 6974 20496
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 1582 5772 1638 5808
rect 1582 5752 1584 5772
rect 1584 5752 1636 5772
rect 1636 5752 1638 5772
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 19706 22616 19762 22672
rect 18602 21664 18658 21720
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18970 21256 19026 21312
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 19522 20848 19578 20904
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 20810 20324 20866 20360
rect 20810 20304 20812 20324
rect 20812 20304 20864 20324
rect 20864 20304 20866 20324
rect 21362 19896 21418 19952
rect 19798 12552 19854 12608
rect 19246 12008 19302 12064
rect 19890 10648 19946 10704
rect 19890 9288 19946 9344
rect 19890 8372 19892 8392
rect 19892 8372 19944 8392
rect 19944 8372 19946 8392
rect 19890 8336 19946 8372
rect 19890 7948 19946 7984
rect 19890 7928 19892 7948
rect 19892 7928 19944 7948
rect 19944 7928 19946 7948
rect 20810 17604 20866 17640
rect 20810 17584 20812 17604
rect 20812 17584 20864 17604
rect 20864 17584 20866 17604
rect 20534 12960 20590 13016
rect 21362 19352 21418 19408
rect 21362 18944 21418 19000
rect 21362 18536 21418 18592
rect 21362 17992 21418 18048
rect 21362 17176 21418 17232
rect 21454 16632 21510 16688
rect 21362 16224 21418 16280
rect 21362 15680 21418 15736
rect 21362 15272 21418 15328
rect 21362 14884 21418 14920
rect 21362 14864 21364 14884
rect 21364 14864 21416 14884
rect 21416 14864 21418 14884
rect 21270 14340 21326 14376
rect 21270 14320 21272 14340
rect 21272 14320 21324 14340
rect 21324 14320 21326 14340
rect 21362 13932 21418 13968
rect 21362 13912 21364 13932
rect 21364 13912 21416 13932
rect 21416 13912 21418 13932
rect 21362 13504 21418 13560
rect 21362 11636 21364 11656
rect 21364 11636 21416 11656
rect 21416 11636 21418 11656
rect 21362 11600 21418 11636
rect 21362 11192 21418 11248
rect 21362 10240 21418 10296
rect 22006 9696 22062 9752
rect 21362 8916 21364 8936
rect 21364 8916 21416 8936
rect 21416 8916 21418 8936
rect 21362 8880 21418 8916
rect 21362 7520 21418 7576
rect 21362 6976 21418 7032
rect 20534 6568 20590 6624
rect 20718 6024 20774 6080
rect 21362 5616 21418 5672
rect 20718 5208 20774 5264
rect 21362 4700 21364 4720
rect 21364 4700 21416 4720
rect 21416 4700 21418 4720
rect 21362 4664 21418 4700
rect 20626 4256 20682 4312
rect 21270 3848 21326 3904
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 20166 1944 20222 2000
rect 21270 3304 21326 3360
rect 21270 2916 21326 2952
rect 21270 2896 21272 2916
rect 21272 2896 21324 2916
rect 21324 2896 21326 2916
rect 20626 1536 20682 1592
rect 19430 992 19486 1048
rect 21270 2352 21326 2408
rect 20718 584 20774 640
rect 22006 176 22062 232
<< metal3 >>
rect 19701 22674 19767 22677
rect 22200 22674 23000 22704
rect 19701 22672 23000 22674
rect 19701 22616 19706 22672
rect 19762 22616 23000 22672
rect 19701 22614 23000 22616
rect 19701 22611 19767 22614
rect 22200 22584 23000 22614
rect 17953 22266 18019 22269
rect 22200 22266 23000 22296
rect 17953 22264 23000 22266
rect 17953 22208 17958 22264
rect 18014 22208 23000 22264
rect 17953 22206 23000 22208
rect 17953 22203 18019 22206
rect 22200 22176 23000 22206
rect 18597 21722 18663 21725
rect 22200 21722 23000 21752
rect 18597 21720 23000 21722
rect 18597 21664 18602 21720
rect 18658 21664 23000 21720
rect 18597 21662 23000 21664
rect 18597 21659 18663 21662
rect 22200 21632 23000 21662
rect 18965 21314 19031 21317
rect 22200 21314 23000 21344
rect 18965 21312 23000 21314
rect 18965 21256 18970 21312
rect 19026 21256 23000 21312
rect 18965 21254 23000 21256
rect 18965 21251 19031 21254
rect 22200 21224 23000 21254
rect 19517 20906 19583 20909
rect 22200 20906 23000 20936
rect 19517 20904 23000 20906
rect 19517 20848 19522 20904
rect 19578 20848 23000 20904
rect 19517 20846 23000 20848
rect 19517 20843 19583 20846
rect 22200 20816 23000 20846
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 6729 20498 6795 20501
rect 6913 20498 6979 20501
rect 6729 20496 6979 20498
rect 6729 20440 6734 20496
rect 6790 20440 6918 20496
rect 6974 20440 6979 20496
rect 6729 20438 6979 20440
rect 6729 20435 6795 20438
rect 6913 20435 6979 20438
rect 20805 20362 20871 20365
rect 22200 20362 23000 20392
rect 20805 20360 23000 20362
rect 20805 20304 20810 20360
rect 20866 20304 23000 20360
rect 20805 20302 23000 20304
rect 20805 20299 20871 20302
rect 22200 20272 23000 20302
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 21357 19954 21423 19957
rect 22200 19954 23000 19984
rect 21357 19952 23000 19954
rect 21357 19896 21362 19952
rect 21418 19896 23000 19952
rect 21357 19894 23000 19896
rect 21357 19891 21423 19894
rect 22200 19864 23000 19894
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 21357 19410 21423 19413
rect 22200 19410 23000 19440
rect 21357 19408 23000 19410
rect 21357 19352 21362 19408
rect 21418 19352 23000 19408
rect 21357 19350 23000 19352
rect 21357 19347 21423 19350
rect 22200 19320 23000 19350
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 21357 19002 21423 19005
rect 22200 19002 23000 19032
rect 21357 19000 23000 19002
rect 21357 18944 21362 19000
rect 21418 18944 23000 19000
rect 21357 18942 23000 18944
rect 21357 18939 21423 18942
rect 22200 18912 23000 18942
rect 21357 18594 21423 18597
rect 22200 18594 23000 18624
rect 21357 18592 23000 18594
rect 21357 18536 21362 18592
rect 21418 18536 23000 18592
rect 21357 18534 23000 18536
rect 21357 18531 21423 18534
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 22200 18504 23000 18534
rect 18270 18463 18590 18464
rect 21357 18050 21423 18053
rect 22200 18050 23000 18080
rect 21357 18048 23000 18050
rect 21357 17992 21362 18048
rect 21418 17992 23000 18048
rect 21357 17990 23000 17992
rect 21357 17987 21423 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 20805 17642 20871 17645
rect 22200 17642 23000 17672
rect 20805 17640 23000 17642
rect 20805 17584 20810 17640
rect 20866 17584 23000 17640
rect 20805 17582 23000 17584
rect 20805 17579 20871 17582
rect 22200 17552 23000 17582
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 0 17234 800 17264
rect 1669 17234 1735 17237
rect 0 17232 1735 17234
rect 0 17176 1674 17232
rect 1730 17176 1735 17232
rect 0 17174 1735 17176
rect 0 17144 800 17174
rect 1669 17171 1735 17174
rect 21357 17234 21423 17237
rect 22200 17234 23000 17264
rect 21357 17232 23000 17234
rect 21357 17176 21362 17232
rect 21418 17176 23000 17232
rect 21357 17174 23000 17176
rect 21357 17171 21423 17174
rect 22200 17144 23000 17174
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 21449 16690 21515 16693
rect 22200 16690 23000 16720
rect 21449 16688 23000 16690
rect 21449 16632 21454 16688
rect 21510 16632 23000 16688
rect 21449 16630 23000 16632
rect 21449 16627 21515 16630
rect 22200 16600 23000 16630
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 21357 16282 21423 16285
rect 22200 16282 23000 16312
rect 21357 16280 23000 16282
rect 21357 16224 21362 16280
rect 21418 16224 23000 16280
rect 21357 16222 23000 16224
rect 21357 16219 21423 16222
rect 22200 16192 23000 16222
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 21357 15738 21423 15741
rect 22200 15738 23000 15768
rect 21357 15736 23000 15738
rect 21357 15680 21362 15736
rect 21418 15680 23000 15736
rect 21357 15678 23000 15680
rect 21357 15675 21423 15678
rect 22200 15648 23000 15678
rect 21357 15330 21423 15333
rect 22200 15330 23000 15360
rect 21357 15328 23000 15330
rect 21357 15272 21362 15328
rect 21418 15272 23000 15328
rect 21357 15270 23000 15272
rect 21357 15267 21423 15270
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 22200 15240 23000 15270
rect 18270 15199 18590 15200
rect 21357 14922 21423 14925
rect 22200 14922 23000 14952
rect 21357 14920 23000 14922
rect 21357 14864 21362 14920
rect 21418 14864 23000 14920
rect 21357 14862 23000 14864
rect 21357 14859 21423 14862
rect 22200 14832 23000 14862
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 21265 14378 21331 14381
rect 22200 14378 23000 14408
rect 21265 14376 23000 14378
rect 21265 14320 21270 14376
rect 21326 14320 23000 14376
rect 21265 14318 23000 14320
rect 21265 14315 21331 14318
rect 22200 14288 23000 14318
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 21357 13970 21423 13973
rect 22200 13970 23000 14000
rect 21357 13968 23000 13970
rect 21357 13912 21362 13968
rect 21418 13912 23000 13968
rect 21357 13910 23000 13912
rect 21357 13907 21423 13910
rect 22200 13880 23000 13910
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 21357 13562 21423 13565
rect 22200 13562 23000 13592
rect 21357 13560 23000 13562
rect 21357 13504 21362 13560
rect 21418 13504 23000 13560
rect 21357 13502 23000 13504
rect 21357 13499 21423 13502
rect 22200 13472 23000 13502
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 20529 13018 20595 13021
rect 22200 13018 23000 13048
rect 20529 13016 23000 13018
rect 20529 12960 20534 13016
rect 20590 12960 23000 13016
rect 20529 12958 23000 12960
rect 20529 12955 20595 12958
rect 22200 12928 23000 12958
rect 19793 12610 19859 12613
rect 22200 12610 23000 12640
rect 19793 12608 23000 12610
rect 19793 12552 19798 12608
rect 19854 12552 23000 12608
rect 19793 12550 23000 12552
rect 19793 12547 19859 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 22200 12520 23000 12550
rect 14805 12479 15125 12480
rect 19241 12066 19307 12069
rect 22200 12066 23000 12096
rect 19241 12064 23000 12066
rect 19241 12008 19246 12064
rect 19302 12008 23000 12064
rect 19241 12006 23000 12008
rect 19241 12003 19307 12006
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 22200 11976 23000 12006
rect 18270 11935 18590 11936
rect 21357 11658 21423 11661
rect 22200 11658 23000 11688
rect 21357 11656 23000 11658
rect 21357 11600 21362 11656
rect 21418 11600 23000 11656
rect 21357 11598 23000 11600
rect 21357 11595 21423 11598
rect 22200 11568 23000 11598
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 21357 11250 21423 11253
rect 22200 11250 23000 11280
rect 21357 11248 23000 11250
rect 21357 11192 21362 11248
rect 21418 11192 23000 11248
rect 21357 11190 23000 11192
rect 21357 11187 21423 11190
rect 22200 11160 23000 11190
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 19885 10706 19951 10709
rect 22200 10706 23000 10736
rect 19885 10704 23000 10706
rect 19885 10648 19890 10704
rect 19946 10648 23000 10704
rect 19885 10646 23000 10648
rect 19885 10643 19951 10646
rect 22200 10616 23000 10646
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 21357 10298 21423 10301
rect 22200 10298 23000 10328
rect 21357 10296 23000 10298
rect 21357 10240 21362 10296
rect 21418 10240 23000 10296
rect 21357 10238 23000 10240
rect 21357 10235 21423 10238
rect 22200 10208 23000 10238
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 22001 9754 22067 9757
rect 22200 9754 23000 9784
rect 22001 9752 23000 9754
rect 22001 9696 22006 9752
rect 22062 9696 23000 9752
rect 22001 9694 23000 9696
rect 22001 9691 22067 9694
rect 22200 9664 23000 9694
rect 19885 9346 19951 9349
rect 22200 9346 23000 9376
rect 19885 9344 23000 9346
rect 19885 9288 19890 9344
rect 19946 9288 23000 9344
rect 19885 9286 23000 9288
rect 19885 9283 19951 9286
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 22200 9256 23000 9286
rect 14805 9215 15125 9216
rect 21357 8938 21423 8941
rect 22200 8938 23000 8968
rect 21357 8936 23000 8938
rect 21357 8880 21362 8936
rect 21418 8880 23000 8936
rect 21357 8878 23000 8880
rect 21357 8875 21423 8878
rect 22200 8848 23000 8878
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 19885 8394 19951 8397
rect 22200 8394 23000 8424
rect 19885 8392 23000 8394
rect 19885 8336 19890 8392
rect 19946 8336 23000 8392
rect 19885 8334 23000 8336
rect 19885 8331 19951 8334
rect 22200 8304 23000 8334
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 19885 7986 19951 7989
rect 22200 7986 23000 8016
rect 19885 7984 23000 7986
rect 19885 7928 19890 7984
rect 19946 7928 23000 7984
rect 19885 7926 23000 7928
rect 19885 7923 19951 7926
rect 22200 7896 23000 7926
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 21357 7578 21423 7581
rect 22200 7578 23000 7608
rect 21357 7576 23000 7578
rect 21357 7520 21362 7576
rect 21418 7520 23000 7576
rect 21357 7518 23000 7520
rect 21357 7515 21423 7518
rect 22200 7488 23000 7518
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 21357 7034 21423 7037
rect 22200 7034 23000 7064
rect 21357 7032 23000 7034
rect 21357 6976 21362 7032
rect 21418 6976 23000 7032
rect 21357 6974 23000 6976
rect 21357 6971 21423 6974
rect 22200 6944 23000 6974
rect 20529 6626 20595 6629
rect 22200 6626 23000 6656
rect 20529 6624 23000 6626
rect 20529 6568 20534 6624
rect 20590 6568 23000 6624
rect 20529 6566 23000 6568
rect 20529 6563 20595 6566
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 22200 6536 23000 6566
rect 18270 6495 18590 6496
rect 20713 6082 20779 6085
rect 22200 6082 23000 6112
rect 20713 6080 23000 6082
rect 20713 6024 20718 6080
rect 20774 6024 23000 6080
rect 20713 6022 23000 6024
rect 20713 6019 20779 6022
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 22200 5992 23000 6022
rect 14805 5951 15125 5952
rect 0 5810 800 5840
rect 1577 5810 1643 5813
rect 0 5808 1643 5810
rect 0 5752 1582 5808
rect 1638 5752 1643 5808
rect 0 5750 1643 5752
rect 0 5720 800 5750
rect 1577 5747 1643 5750
rect 21357 5674 21423 5677
rect 22200 5674 23000 5704
rect 21357 5672 23000 5674
rect 21357 5616 21362 5672
rect 21418 5616 23000 5672
rect 21357 5614 23000 5616
rect 21357 5611 21423 5614
rect 22200 5584 23000 5614
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 20713 5266 20779 5269
rect 22200 5266 23000 5296
rect 20713 5264 23000 5266
rect 20713 5208 20718 5264
rect 20774 5208 23000 5264
rect 20713 5206 23000 5208
rect 20713 5203 20779 5206
rect 22200 5176 23000 5206
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 21357 4722 21423 4725
rect 22200 4722 23000 4752
rect 21357 4720 23000 4722
rect 21357 4664 21362 4720
rect 21418 4664 23000 4720
rect 21357 4662 23000 4664
rect 21357 4659 21423 4662
rect 22200 4632 23000 4662
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 20621 4314 20687 4317
rect 22200 4314 23000 4344
rect 20621 4312 23000 4314
rect 20621 4256 20626 4312
rect 20682 4256 23000 4312
rect 20621 4254 23000 4256
rect 20621 4251 20687 4254
rect 22200 4224 23000 4254
rect 21265 3906 21331 3909
rect 22200 3906 23000 3936
rect 21265 3904 23000 3906
rect 21265 3848 21270 3904
rect 21326 3848 23000 3904
rect 21265 3846 23000 3848
rect 21265 3843 21331 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22200 3816 23000 3846
rect 14805 3775 15125 3776
rect 21265 3362 21331 3365
rect 22200 3362 23000 3392
rect 21265 3360 23000 3362
rect 21265 3304 21270 3360
rect 21326 3304 23000 3360
rect 21265 3302 23000 3304
rect 21265 3299 21331 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 22200 3272 23000 3302
rect 18270 3231 18590 3232
rect 21265 2954 21331 2957
rect 22200 2954 23000 2984
rect 21265 2952 23000 2954
rect 21265 2896 21270 2952
rect 21326 2896 23000 2952
rect 21265 2894 23000 2896
rect 21265 2891 21331 2894
rect 22200 2864 23000 2894
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 21265 2410 21331 2413
rect 22200 2410 23000 2440
rect 21265 2408 23000 2410
rect 21265 2352 21270 2408
rect 21326 2352 23000 2408
rect 21265 2350 23000 2352
rect 21265 2347 21331 2350
rect 22200 2320 23000 2350
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 20161 2002 20227 2005
rect 22200 2002 23000 2032
rect 20161 2000 23000 2002
rect 20161 1944 20166 2000
rect 20222 1944 23000 2000
rect 20161 1942 23000 1944
rect 20161 1939 20227 1942
rect 22200 1912 23000 1942
rect 20621 1594 20687 1597
rect 22200 1594 23000 1624
rect 20621 1592 23000 1594
rect 20621 1536 20626 1592
rect 20682 1536 23000 1592
rect 20621 1534 23000 1536
rect 20621 1531 20687 1534
rect 22200 1504 23000 1534
rect 19425 1050 19491 1053
rect 22200 1050 23000 1080
rect 19425 1048 23000 1050
rect 19425 992 19430 1048
rect 19486 992 23000 1048
rect 19425 990 23000 992
rect 19425 987 19491 990
rect 22200 960 23000 990
rect 20713 642 20779 645
rect 22200 642 23000 672
rect 20713 640 23000 642
rect 20713 584 20718 640
rect 20774 584 23000 640
rect 20713 582 23000 584
rect 20713 579 20779 582
rect 22200 552 23000 582
rect 22001 234 22067 237
rect 22200 234 23000 264
rect 22001 232 23000 234
rect 22001 176 22006 232
rect 22062 176 23000 232
rect 22001 174 23000 176
rect 22001 171 22067 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1624635492
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1624635492
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 3772 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1624635492
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1624635492
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_30
timestamp 1624635492
transform 1 0 3864 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1624635492
transform 1 0 4968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_42
timestamp 1624635492
transform 1 0 4968 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_54
timestamp 1624635492
transform 1 0 6072 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1624635492
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1624635492
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_66
timestamp 1624635492
transform 1 0 7176 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 8280 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 9016 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_88
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_100
timestamp 1624635492
transform 1 0 10304 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_87
timestamp 1624635492
transform 1 0 9108 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_99
timestamp 1624635492
transform 1 0 10212 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1624635492
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_111
timestamp 1624635492
transform 1 0 11316 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1624635492
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 14260 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_129
timestamp 1624635492
transform 1 0 12972 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1624635492
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_135
timestamp 1624635492
transform 1 0 13524 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_144
timestamp 1624635492
transform 1 0 14352 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_146
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_158
timestamp 1624635492
transform 1 0 15640 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_156
timestamp 1624635492
transform 1 0 15456 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1624635492
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_175
timestamp 1624635492
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_187 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_168
timestamp 1624635492
transform 1 0 16560 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_180
timestamp 1624635492
transform 1 0 17664 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 18952 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_194
timestamp 1624635492
transform 1 0 18952 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_195
timestamp 1624635492
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 19320 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 19044 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 19596 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_198
timestamp 1624635492
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_201
timestamp 1624635492
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform -1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 19504 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1624635492
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_204
timestamp 1624635492
transform 1 0 19872 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1624635492
transform -1 0 20332 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1624635492
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1624635492
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1624635492
transform -1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1624635492
transform -1 0 20884 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_215
timestamp 1624635492
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1624635492
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1624635492
transform -1 0 21436 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1624635492
transform -1 0 21436 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1624635492
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1624635492
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1624635492
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1624635492
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1624635492
transform 1 0 3588 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1624635492
transform 1 0 4692 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 6348 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_51
timestamp 1624635492
transform 1 0 5796 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_58
timestamp 1624635492
transform 1 0 6440 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_70
timestamp 1624635492
transform 1 0 7544 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_82
timestamp 1624635492
transform 1 0 8648 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_94
timestamp 1624635492
transform 1 0 9752 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 11592 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_106
timestamp 1624635492
transform 1 0 10856 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_115
timestamp 1624635492
transform 1 0 11684 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_127
timestamp 1624635492
transform 1 0 12788 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_139
timestamp 1624635492
transform 1 0 13892 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_151
timestamp 1624635492
transform 1 0 14996 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_163
timestamp 1624635492
transform 1 0 16100 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 16836 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_172
timestamp 1624635492
transform 1 0 16928 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1624635492
transform 1 0 18032 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 20332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 19412 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_196 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 19136 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_199
timestamp 1624635492
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1624635492
transform 1 0 19780 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1624635492
transform -1 0 21436 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1624635492
transform -1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1624635492
transform 1 0 20332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1624635492
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1624635492
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1624635492
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_27
timestamp 1624635492
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_30
timestamp 1624635492
transform 1 0 3864 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_42
timestamp 1624635492
transform 1 0 4968 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_54
timestamp 1624635492
transform 1 0 6072 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_66
timestamp 1624635492
transform 1 0 7176 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_78
timestamp 1624635492
transform 1 0 8280 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 9016 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_87
timestamp 1624635492
transform 1 0 9108 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_99
timestamp 1624635492
transform 1 0 10212 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_111
timestamp 1624635492
transform 1 0 11316 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1624635492
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 14260 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_135
timestamp 1624635492
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_144
timestamp 1624635492
transform 1 0 14352 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_156
timestamp 1624635492
transform 1 0 15456 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_168
timestamp 1624635492
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_180
timestamp 1624635492
transform 1 0 17664 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 19504 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 20424 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 20056 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_192
timestamp 1624635492
transform 1 0 18768 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_201
timestamp 1624635492
transform 1 0 19596 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_206
timestamp 1624635492
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 20884 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1624635492
transform -1 0 21436 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_210
timestamp 1624635492
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_215
timestamp 1624635492
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1624635492
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1624635492
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1624635492
transform 1 0 3588 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1624635492
transform 1 0 4692 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 6348 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_51
timestamp 1624635492
transform 1 0 5796 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_58
timestamp 1624635492
transform 1 0 6440 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_70
timestamp 1624635492
transform 1 0 7544 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_82
timestamp 1624635492
transform 1 0 8648 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_94
timestamp 1624635492
transform 1 0 9752 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 11592 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_106
timestamp 1624635492
transform 1 0 10856 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_115
timestamp 1624635492
transform 1 0 11684 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_127
timestamp 1624635492
transform 1 0 12788 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_139
timestamp 1624635492
transform 1 0 13892 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_151
timestamp 1624635492
transform 1 0 14996 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_163
timestamp 1624635492
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 16836 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_172
timestamp 1624635492
transform 1 0 16928 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1624635492
transform 1 0 18032 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1624635492
transform 1 0 19136 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_208
timestamp 1624635492
transform 1 0 20240 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _87_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 21068 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 21436 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_217
timestamp 1624635492
transform 1 0 21068 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1624635492
transform 1 0 21436 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1624635492
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 3772 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_27
timestamp 1624635492
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_30
timestamp 1624635492
transform 1 0 3864 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_42
timestamp 1624635492
transform 1 0 4968 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_54
timestamp 1624635492
transform 1 0 6072 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_66
timestamp 1624635492
transform 1 0 7176 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_78
timestamp 1624635492
transform 1 0 8280 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 9016 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_87
timestamp 1624635492
transform 1 0 9108 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_99
timestamp 1624635492
transform 1 0 10212 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_111
timestamp 1624635492
transform 1 0 11316 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1624635492
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 14260 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_135
timestamp 1624635492
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_144
timestamp 1624635492
transform 1 0 14352 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_156
timestamp 1624635492
transform 1 0 15456 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_168
timestamp 1624635492
transform 1 0 16560 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_180
timestamp 1624635492
transform 1 0 17664 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 19504 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_192
timestamp 1624635492
transform 1 0 18768 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_201
timestamp 1624635492
transform 1 0 19596 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1624635492
transform -1 0 21436 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1624635492
transform -1 0 20976 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 20516 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_211
timestamp 1624635492
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_216
timestamp 1624635492
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1624635492
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624635492
transform -1 0 1840 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_8
timestamp 1624635492
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_12
timestamp 1624635492
transform 1 0 2208 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1624635492
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 3772 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_24
timestamp 1624635492
transform 1 0 3312 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_36
timestamp 1624635492
transform 1 0 4416 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_27
timestamp 1624635492
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_30
timestamp 1624635492
transform 1 0 3864 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 6348 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_48
timestamp 1624635492
transform 1 0 5520 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_56
timestamp 1624635492
transform 1 0 6256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_58
timestamp 1624635492
transform 1 0 6440 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_42
timestamp 1624635492
transform 1 0 4968 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_54
timestamp 1624635492
transform 1 0 6072 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_70
timestamp 1624635492
transform 1 0 7544 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_82
timestamp 1624635492
transform 1 0 8648 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_66
timestamp 1624635492
transform 1 0 7176 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_78
timestamp 1624635492
transform 1 0 8280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 9016 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_94
timestamp 1624635492
transform 1 0 9752 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_87
timestamp 1624635492
transform 1 0 9108 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_99
timestamp 1624635492
transform 1 0 10212 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 11592 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_106
timestamp 1624635492
transform 1 0 10856 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_115
timestamp 1624635492
transform 1 0 11684 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_111
timestamp 1624635492
transform 1 0 11316 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1624635492
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 14260 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_127
timestamp 1624635492
transform 1 0 12788 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1624635492
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_135
timestamp 1624635492
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_144
timestamp 1624635492
transform 1 0 14352 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_151
timestamp 1624635492
transform 1 0 14996 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_163
timestamp 1624635492
transform 1 0 16100 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_156
timestamp 1624635492
transform 1 0 15456 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 16836 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_172
timestamp 1624635492
transform 1 0 16928 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1624635492
transform 1 0 18032 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_168
timestamp 1624635492
transform 1 0 16560 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_180
timestamp 1624635492
transform 1 0 17664 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 19504 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1624635492
transform 1 0 19136 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1624635492
transform 1 0 20240 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_192
timestamp 1624635492
transform 1 0 18768 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_201
timestamp 1624635492
transform 1 0 19596 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_211
timestamp 1624635492
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 20516 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1624635492
transform -1 0 20976 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_216
timestamp 1624635492
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_218
timestamp 1624635492
transform 1 0 21160 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1624635492
transform 1 0 21160 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _69_
timestamp 1624635492
transform -1 0 21160 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1624635492
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1624635492
transform 1 0 21528 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1624635492
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1624635492
transform 1 0 3588 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1624635492
transform 1 0 4692 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 6348 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_51
timestamp 1624635492
transform 1 0 5796 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_58
timestamp 1624635492
transform 1 0 6440 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 8188 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_8_70
timestamp 1624635492
transform 1 0 7544 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_76
timestamp 1624635492
transform 1 0 8096 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1624635492
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 11592 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_105
timestamp 1624635492
transform 1 0 10764 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_109
timestamp 1624635492
transform 1 0 11132 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_112
timestamp 1624635492
transform 1 0 11408 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_115
timestamp 1624635492
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15272 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 14260 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_126
timestamp 1624635492
transform 1 0 12696 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_138
timestamp 1624635492
transform 1 0 13800 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_143
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1624635492
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_166
timestamp 1624635492
transform 1 0 16376 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1624635492
transform 1 0 17664 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 16836 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_170
timestamp 1624635492
transform 1 0 16744 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_172
timestamp 1624635492
transform 1 0 16928 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_178
timestamp 1624635492
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 20148 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_189
timestamp 1624635492
transform 1 0 18492 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_201
timestamp 1624635492
transform 1 0 19596 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_207
timestamp 1624635492
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _71_
timestamp 1624635492
transform -1 0 21068 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1624635492
transform 1 0 20332 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 21436 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1624635492
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_217
timestamp 1624635492
transform 1 0 21068 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1624635492
transform 1 0 21436 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1624635492
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1624635492
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_30
timestamp 1624635492
transform 1 0 3864 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_42
timestamp 1624635492
transform 1 0 4968 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_54
timestamp 1624635492
transform 1 0 6072 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_66
timestamp 1624635492
transform 1 0 7176 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_78
timestamp 1624635492
transform 1 0 8280 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9660 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 9016 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_87
timestamp 1624635492
transform 1 0 9108 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 11684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11868 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1624635492
transform 1 0 11132 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_115
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 14260 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_133
timestamp 1624635492
transform 1 0 13340 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_141
timestamp 1624635492
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_144
timestamp 1624635492
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1624635492
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15364 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_9_149
timestamp 1624635492
transform 1 0 14812 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17020 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_171
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 19504 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 20148 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_189
timestamp 1624635492
transform 1 0 18492 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_197
timestamp 1624635492
transform 1 0 19228 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_201
timestamp 1624635492
transform 1 0 19596 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_207
timestamp 1624635492
transform 1 0 20148 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _73_
timestamp 1624635492
transform -1 0 21068 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1624635492
transform -1 0 20608 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1624635492
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_217
timestamp 1624635492
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1624635492
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1624635492
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1624635492
transform 1 0 3588 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1624635492
transform 1 0 4692 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_51
timestamp 1624635492
transform 1 0 5796 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_58
timestamp 1624635492
transform 1 0 6440 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_70
timestamp 1624635492
transform 1 0 7544 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_82
timestamp 1624635492
transform 1 0 8648 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_94
timestamp 1624635492
transform 1 0 9752 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11868 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 11592 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_106
timestamp 1624635492
transform 1 0 10856 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_115
timestamp 1624635492
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 13616 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_126
timestamp 1624635492
transform 1 0 12696 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_134
timestamp 1624635492
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_152
timestamp 1624635492
transform 1 0 15088 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_164
timestamp 1624635492
transform 1 0 16192 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 18216 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 17112 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 16836 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1624635492
transform 1 0 16744 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_172
timestamp 1624635492
transform 1 0 16928 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_183
timestamp 1624635492
transform 1 0 17940 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1624635492
transform -1 0 20148 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_202
timestamp 1624635492
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_207
timestamp 1624635492
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _74_
timestamp 1624635492
transform -1 0 21068 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1624635492
transform -1 0 20608 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1624635492
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_217
timestamp 1624635492
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1624635492
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1624635492
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 3772 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_27
timestamp 1624635492
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_30
timestamp 1624635492
transform 1 0 3864 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_42
timestamp 1624635492
transform 1 0 4968 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_54
timestamp 1624635492
transform 1 0 6072 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_66
timestamp 1624635492
transform 1 0 7176 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_78
timestamp 1624635492
transform 1 0 8280 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 9016 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_87
timestamp 1624635492
transform 1 0 9108 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_99
timestamp 1624635492
transform 1 0 10212 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11500 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_107
timestamp 1624635492
transform 1 0 10948 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1624635492
transform 1 0 11500 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_125
timestamp 1624635492
transform 1 0 12604 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _70_
timestamp 1624635492
transform -1 0 13524 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 13708 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 14260 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp 1624635492
transform 1 0 13156 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_135
timestamp 1624635492
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_140
timestamp 1624635492
transform 1 0 13984 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_144
timestamp 1624635492
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14536 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 16192 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_155
timestamp 1624635492
transform 1 0 15364 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_163
timestamp 1624635492
transform 1 0 16100 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1624635492
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_167
timestamp 1624635492
transform 1 0 16468 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_175
timestamp 1624635492
transform 1 0 17204 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1624635492
transform 1 0 17756 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 19504 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1624635492
transform -1 0 20148 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 19320 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_193
timestamp 1624635492
transform 1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_198
timestamp 1624635492
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_201
timestamp 1624635492
transform 1 0 19596 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_207
timestamp 1624635492
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _75_
timestamp 1624635492
transform -1 0 21068 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1624635492
transform -1 0 20608 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1624635492
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1624635492
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1624635492
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1624635492
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1624635492
transform 1 0 3588 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1624635492
transform 1 0 4692 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 6348 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_51
timestamp 1624635492
transform 1 0 5796 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_58
timestamp 1624635492
transform 1 0 6440 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_70
timestamp 1624635492
transform 1 0 7544 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_82
timestamp 1624635492
transform 1 0 8648 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_94
timestamp 1624635492
transform 1 0 9752 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _68_
timestamp 1624635492
transform 1 0 11868 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 11592 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_106
timestamp 1624635492
transform 1 0 10856 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_115
timestamp 1624635492
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_120
timestamp 1624635492
transform 1 0 12144 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_132
timestamp 1624635492
transform 1 0 13248 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _72_
timestamp 1624635492
transform -1 0 16008 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_156
timestamp 1624635492
transform 1 0 15456 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_162
timestamp 1624635492
transform 1 0 16008 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 16836 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_170
timestamp 1624635492
transform 1 0 16744 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_172
timestamp 1624635492
transform 1 0 16928 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_184
timestamp 1624635492
transform 1 0 18032 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1624635492
transform -1 0 20148 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 19688 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_196
timestamp 1624635492
transform 1 0 19136 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_202
timestamp 1624635492
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_207
timestamp 1624635492
transform 1 0 20148 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _76_
timestamp 1624635492
transform -1 0 21068 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1624635492
transform -1 0 20608 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1624635492
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_217
timestamp 1624635492
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1624635492
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1624635492
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1624635492
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 3772 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1624635492
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_30
timestamp 1624635492
transform 1 0 3864 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1624635492
transform 1 0 3588 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_39
timestamp 1624635492
transform 1 0 4692 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 6348 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_42
timestamp 1624635492
transform 1 0 4968 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_54
timestamp 1624635492
transform 1 0 6072 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_51
timestamp 1624635492
transform 1 0 5796 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_58
timestamp 1624635492
transform 1 0 6440 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 8004 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_13_66
timestamp 1624635492
transform 1 0 7176 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_78
timestamp 1624635492
transform 1 0 8280 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_70
timestamp 1624635492
transform 1 0 7544 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_74
timestamp 1624635492
transform 1 0 7912 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 11408 0 -1 10336
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 9016 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 9108 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_89
timestamp 1624635492
transform 1 0 9292 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_101
timestamp 1624635492
transform 1 0 10396 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_91
timestamp 1624635492
transform 1 0 9476 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 13248 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 11592 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp 1624635492
transform 1 0 11500 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_112
timestamp 1624635492
transform 1 0 11408 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_115
timestamp 1624635492
transform 1 0 11684 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14076 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13064 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 14260 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 13432 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1624635492
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_141
timestamp 1624635492
transform 1 0 14076 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_127
timestamp 1624635492
transform 1 0 12788 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_139
timestamp 1624635492
transform 1 0 13892 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1624635492
transform 1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1624635492
transform 1 0 14812 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_146
timestamp 1624635492
transform 1 0 14536 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 1624635492
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1624635492
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_157
timestamp 1624635492
transform 1 0 15548 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 18676 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 16836 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_167
timestamp 1624635492
transform 1 0 16468 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_173
timestamp 1624635492
transform 1 0 17020 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_169
timestamp 1624635492
transform 1 0 16652 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_172
timestamp 1624635492
transform 1 0 16928 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_184
timestamp 1624635492
transform 1 0 18032 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 18768 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1624635492
transform 1 0 19780 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 19504 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 1624635492
transform 1 0 18676 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_195
timestamp 1624635492
transform 1 0 19044 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_198
timestamp 1624635492
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_201
timestamp 1624635492
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_208
timestamp 1624635492
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_213
timestamp 1624635492
transform 1 0 20700 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1624635492
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _78_
timestamp 1624635492
transform -1 0 21160 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _77_
timestamp 1624635492
transform -1 0 21068 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1624635492
transform 1 0 20424 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_222
timestamp 1624635492
transform 1 0 21528 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_218
timestamp 1624635492
transform 1 0 21160 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1624635492
transform 1 0 21068 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1624635492
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 3772 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_27
timestamp 1624635492
transform 1 0 3588 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_30
timestamp 1624635492
transform 1 0 3864 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_42
timestamp 1624635492
transform 1 0 4968 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_54
timestamp 1624635492
transform 1 0 6072 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1624635492
transform -1 0 8832 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_66
timestamp 1624635492
transform 1 0 7176 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_74
timestamp 1624635492
transform 1 0 7912 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1624635492
transform -1 0 10856 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 9016 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1
timestamp 1624635492
transform -1 0 9936 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1624635492
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_87
timestamp 1624635492
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1624635492
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_100
timestamp 1624635492
transform 1 0 10304 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1624635492
transform 1 0 11040 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 12052 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1624635492
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_117
timestamp 1624635492
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_121
timestamp 1624635492
transform 1 0 12236 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1624635492
transform 1 0 12604 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13800 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 14260 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_138
timestamp 1624635492
transform 1 0 13800 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_142
timestamp 1624635492
transform 1 0 14168 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 17572 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_146
timestamp 1624635492
transform 1 0 14536 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_158
timestamp 1624635492
transform 1 0 15640 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_162
timestamp 1624635492
transform 1 0 16008 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp 1624635492
transform -1 0 18400 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1624635492
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1624635492
transform 1 0 19780 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 19504 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1624635492
transform 1 0 18400 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_192
timestamp 1624635492
transform 1 0 18768 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_195
timestamp 1624635492
transform 1 0 19044 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp 1624635492
transform 1 0 19412 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_201
timestamp 1624635492
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _79_
timestamp 1624635492
transform -1 0 21068 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1624635492
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1624635492
transform 1 0 21068 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1624635492
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1624635492
transform 1 0 3588 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_39
timestamp 1624635492
transform 1 0 4692 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_51
timestamp 1624635492
transform 1 0 5796 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_58
timestamp 1624635492
transform 1 0 6440 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1624635492
transform -1 0 8832 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_70
timestamp 1624635492
transform 1 0 7544 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_74
timestamp 1624635492
transform 1 0 7912 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1624635492
transform -1 0 9844 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11224 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1624635492
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_95
timestamp 1624635492
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_99
timestamp 1624635492
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 11592 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_110
timestamp 1624635492
transform 1 0 11224 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_115
timestamp 1624635492
transform 1 0 11684 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1624635492
transform -1 0 13984 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_16_127
timestamp 1624635492
transform 1 0 12788 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_140
timestamp 1624635492
transform 1 0 13984 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_right_track_0.prog_clk
timestamp 1624635492
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_149
timestamp 1624635492
transform 1 0 14812 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_161
timestamp 1624635492
transform 1 0 15916 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 18032 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 16836 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_169
timestamp 1624635492
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_172
timestamp 1624635492
transform 1 0 16928 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_182
timestamp 1624635492
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 19044 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1624635492
transform -1 0 20148 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 19688 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_193
timestamp 1624635492
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_198
timestamp 1624635492
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_202
timestamp 1624635492
transform 1 0 19688 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_207
timestamp 1624635492
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _81_
timestamp 1624635492
transform -1 0 21068 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1624635492
transform 1 0 20332 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform 1 0 21252 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1624635492
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 1624635492
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1624635492
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1624635492
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624635492
transform 1 0 3772 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1624635492
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_30
timestamp 1624635492
transform 1 0 3864 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_42
timestamp 1624635492
transform 1 0 4968 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_54
timestamp 1624635492
transform 1 0 6072 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_66
timestamp 1624635492
transform 1 0 7176 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_78
timestamp 1624635492
transform 1 0 8280 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 9292 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624635492
transform 1 0 9016 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1624635492
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1624635492
transform -1 0 11776 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_105
timestamp 1624635492
transform 1 0 10764 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_116
timestamp 1624635492
transform 1 0 11776 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_124
timestamp 1624635492
transform 1 0 12512 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1624635492
transform 1 0 13156 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624635492
transform 1 0 14260 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_129
timestamp 1624635492
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_140
timestamp 1624635492
transform 1 0 13984 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 16284 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_146
timestamp 1624635492
transform 1 0 14536 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_165
timestamp 1624635492
transform 1 0 16284 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 17388 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_186
timestamp 1624635492
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1624635492
transform 1 0 18400 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _80_
timestamp 1624635492
transform -1 0 19320 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624635492
transform 1 0 19504 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1624635492
transform -1 0 20148 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_191
timestamp 1624635492
transform 1 0 18676 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_198
timestamp 1624635492
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_201
timestamp 1624635492
transform 1 0 19596 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_207
timestamp 1624635492
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _82_
timestamp 1624635492
transform -1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1624635492
transform -1 0 20608 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1624635492
transform 1 0 20608 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1624635492
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1624635492
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1624635492
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_27
timestamp 1624635492
transform 1 0 3588 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_39
timestamp 1624635492
transform 1 0 4692 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624635492
transform 1 0 6348 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_51
timestamp 1624635492
transform 1 0 5796 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_58
timestamp 1624635492
transform 1 0 6440 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_right_track_0.prog_clk
timestamp 1624635492
transform 1 0 8464 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_70
timestamp 1624635492
transform 1 0 7544 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_78
timestamp 1624635492
transform 1 0 8280 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_83
timestamp 1624635492
transform 1 0 8740 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_95
timestamp 1624635492
transform 1 0 9844 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1624635492
transform 1 0 11040 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12144 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624635492
transform 1 0 11592 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_105
timestamp 1624635492
transform 1 0 10764 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_111
timestamp 1624635492
transform 1 0 11316 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_115
timestamp 1624635492
transform 1 0 11684 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_120
timestamp 1624635492
transform 1 0 12144 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 14536 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_128
timestamp 1624635492
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16652 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_18_146
timestamp 1624635492
transform 1 0 14536 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_158
timestamp 1624635492
transform 1 0 15640 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17112 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624635492
transform 1 0 16836 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 18124 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_169
timestamp 1624635492
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_172
timestamp 1624635492
transform 1 0 16928 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_183
timestamp 1624635492
transform 1 0 17940 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1624635492
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20056 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1624635492
transform -1 0 19596 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 19136 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_191
timestamp 1624635492
transform 1 0 18676 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_196
timestamp 1624635492
transform 1 0 19136 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp 1624635492
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_206
timestamp 1624635492
transform 1 0 20056 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _83_
timestamp 1624635492
transform -1 0 21068 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _84_
timestamp 1624635492
transform -1 0 20608 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1624635492
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_217
timestamp 1624635492
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1624635492
transform 1 0 21436 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1624635492
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1624635492
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624635492
transform 1 0 3772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_27
timestamp 1624635492
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_30
timestamp 1624635492
transform 1 0 3864 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_27
timestamp 1624635492
transform 1 0 3588 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_39
timestamp 1624635492
transform 1 0 4692 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 8096 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624635492
transform 1 0 6348 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_42
timestamp 1624635492
transform 1 0 4968 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_54
timestamp 1624635492
transform 1 0 6072 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_51
timestamp 1624635492
transform 1 0 5796 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_58
timestamp 1624635492
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1624635492
transform -1 0 9384 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_19_66
timestamp 1624635492
transform 1 0 7176 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_78
timestamp 1624635492
transform 1 0 8280 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_76
timestamp 1624635492
transform 1 0 8096 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_80
timestamp 1624635492
transform 1 0 8464 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 11040 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1624635492
transform 1 0 9752 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624635492
transform 1 0 9016 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_87
timestamp 1624635492
transform 1 0 9108 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_93
timestamp 1624635492
transform 1 0 9660 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_103
timestamp 1624635492
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1624635492
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10764 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1624635492
transform -1 0 13064 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624635492
transform 1 0 11592 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_121
timestamp 1624635492
transform 1 0 12236 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_108
timestamp 1624635492
transform 1 0 11040 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_115
timestamp 1624635492
transform 1 0 11684 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_135
timestamp 1624635492
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_130
timestamp 1624635492
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_133
timestamp 1624635492
transform 1 0 13340 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_right_track_0.prog_clk
timestamp 1624635492
transform -1 0 13524 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_139
timestamp 1624635492
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_139
timestamp 1624635492
transform 1 0 13892 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 14076 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624635492
transform 1 0 14260 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 13892 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_143
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_144
timestamp 1624635492
transform 1 0 14352 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 15916 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1624635492
transform 1 0 15456 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_160
timestamp 1624635492
transform 1 0 15824 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_155
timestamp 1624635492
transform 1 0 15364 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_161
timestamp 1624635492
transform 1 0 15916 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1624635492
transform -1 0 17756 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624635492
transform 1 0 16836 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1624635492
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1624635492
transform 1 0 17756 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_169
timestamp 1624635492
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_174
timestamp 1624635492
transform 1 0 17112 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1624635492
transform 1 0 18216 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_193
timestamp 1624635492
transform 1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 19320 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1624635492
transform -1 0 19412 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_204
timestamp 1624635492
transform 1 0 19872 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1624635492
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_206
timestamp 1624635492
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_201
timestamp 1624635492
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_198
timestamp 1624635492
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1624635492
transform -1 0 20056 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624635492
transform 1 0 19504 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp 1624635492
transform -1 0 20424 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1624635492
transform 1 0 19596 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1624635492
transform -1 0 20516 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1624635492
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1624635492
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp 1624635492
transform 1 0 20608 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1624635492
transform -1 0 20976 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1624635492
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_216
timestamp 1624635492
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output53
timestamp 1624635492
transform 1 0 21068 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1624635492
transform 1 0 21160 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1624635492
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1624635492
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1624635492
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 5612 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624635492
transform 1 0 3772 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_27
timestamp 1624635492
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_30
timestamp 1624635492
transform 1 0 3864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_49
timestamp 1624635492
transform 1 0 5612 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_61
timestamp 1624635492
transform 1 0 6716 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8740 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_83
timestamp 1624635492
transform 1 0 8740 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624635492
transform 1 0 9016 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_track_0.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 12420 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_21_87
timestamp 1624635492
transform 1 0 9108 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_99
timestamp 1624635492
transform 1 0 10212 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12604 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1624635492
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624635492
transform 1 0 14260 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_141
timestamp 1624635492
transform 1 0 14076 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_144
timestamp 1624635492
transform 1 0 14352 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1624635492
transform 1 0 15916 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1624635492
transform -1 0 15732 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 16652 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_159
timestamp 1624635492
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_164
timestamp 1624635492
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17296 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1624635492
transform 1 0 16652 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_175
timestamp 1624635492
transform 1 0 17204 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624635492
transform 1 0 19504 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 20424 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 19780 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 18952 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_192
timestamp 1624635492
transform 1 0 18768 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_196
timestamp 1624635492
transform 1 0 19136 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1624635492
transform 1 0 19780 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_207
timestamp 1624635492
transform 1 0 20148 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1624635492
transform 1 0 20608 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform 1 0 21068 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_210
timestamp 1624635492
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1624635492
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1624635492
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 3956 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1624635492
transform 1 0 4232 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_22_31
timestamp 1624635492
transform 1 0 3956 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624635492
transform 1 0 6348 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_43
timestamp 1624635492
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_47
timestamp 1624635492
transform 1 0 5428 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1624635492
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_58
timestamp 1624635492
transform 1 0 6440 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9108 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_70
timestamp 1624635492
transform 1 0 7544 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9476 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_94
timestamp 1624635492
transform 1 0 9752 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_98
timestamp 1624635492
transform 1 0 10120 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12696 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624635492
transform 1 0 11592 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_110
timestamp 1624635492
transform 1 0 11224 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_115
timestamp 1624635492
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 15088 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_126
timestamp 1624635492
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_130
timestamp 1624635492
transform 1 0 13064 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1624635492
transform -1 0 16100 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_152
timestamp 1624635492
transform 1 0 15088 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_163
timestamp 1624635492
transform 1 0 16100 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18492 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624635492
transform 1 0 16836 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_172
timestamp 1624635492
transform 1 0 16928 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1624635492
transform -1 0 19504 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20240 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_189
timestamp 1624635492
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_200
timestamp 1624635492
transform 1 0 19504 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_204
timestamp 1624635492
transform 1 0 19872 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_208
timestamp 1624635492
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1624635492
transform -1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 21068 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1624635492
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1624635492
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1624635492
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1624635492
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1624635492
transform -1 0 4876 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624635492
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_27
timestamp 1624635492
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_30
timestamp 1624635492
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_41
timestamp 1624635492
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1624635492
transform 1 0 5060 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 7544 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_46
timestamp 1624635492
transform 1 0 5336 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1624635492
transform 1 0 7728 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_70
timestamp 1624635492
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_81
timestamp 1624635492
transform 1 0 8556 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624635492
transform 1 0 9016 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_right_track_0.prog_clk
timestamp 1624635492
transform 1 0 9292 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_85
timestamp 1624635492
transform 1 0 8924 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_87
timestamp 1624635492
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_92
timestamp 1624635492
transform 1 0 9568 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_104
timestamp 1624635492
transform 1 0 10672 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13156 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_23_116
timestamp 1624635492
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624635492
transform 1 0 14260 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_131
timestamp 1624635492
transform 1 0 13156 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1624635492
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_right_track_0.prog_clk
timestamp 1624635492
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1624635492
transform 1 0 14812 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_161
timestamp 1624635492
transform 1 0 15916 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17756 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_173
timestamp 1624635492
transform 1 0 17020 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1624635492
transform -1 0 20424 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624635492
transform 1 0 19504 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_197
timestamp 1624635492
transform 1 0 19228 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_201
timestamp 1624635492
transform 1 0 19596 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1624635492
transform -1 0 20884 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1624635492
transform 1 0 21068 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_210
timestamp 1624635492
transform 1 0 20424 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_215
timestamp 1624635492
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1624635492
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 1840 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1624635492
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1624635492
transform 1 0 1748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_24
timestamp 1624635492
transform 1 0 3312 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_36
timestamp 1624635492
transform 1 0 4416 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624635492
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_48
timestamp 1624635492
transform 1 0 5520 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_56
timestamp 1624635492
transform 1 0 6256 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_58
timestamp 1624635492
transform 1 0 6440 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1624635492
transform 1 0 8096 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1624635492
transform -1 0 7912 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_right_track_0.prog_clk
timestamp 1624635492
transform 1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_64
timestamp 1624635492
transform 1 0 6992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_74
timestamp 1624635492
transform 1 0 7912 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_79
timestamp 1624635492
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1624635492
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_88
timestamp 1624635492
transform 1 0 9200 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_100
timestamp 1624635492
transform 1 0 10304 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624635492
transform 1 0 11592 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_112
timestamp 1624635492
transform 1 0 11408 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_115
timestamp 1624635492
transform 1 0 11684 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_127
timestamp 1624635492
transform 1 0 12788 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_139
timestamp 1624635492
transform 1 0 13892 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 14904 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_147
timestamp 1624635492
transform 1 0 14628 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_152
timestamp 1624635492
transform 1 0 15088 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_164
timestamp 1624635492
transform 1 0 16192 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17112 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624635492
transform 1 0 16836 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_170
timestamp 1624635492
transform 1 0 16744 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_172
timestamp 1624635492
transform 1 0 16928 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20240 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1624635492
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_202
timestamp 1624635492
transform 1 0 19688 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_208
timestamp 1624635492
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1624635492
transform -1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform 1 0 21068 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1624635492
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1624635492
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1624635492
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1624635492
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 6348 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624635492
transform 1 0 3772 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_27
timestamp 1624635492
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_30
timestamp 1624635492
transform 1 0 3864 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_38
timestamp 1624635492
transform 1 0 4600 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1624635492
transform 1 0 7452 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_81
timestamp 1624635492
transform 1 0 8556 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9292 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624635492
transform 1 0 9016 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_85
timestamp 1624635492
transform 1 0 8924 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_87
timestamp 1624635492
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 10948 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 1624635492
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1624635492
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624635492
transform 1 0 14260 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1624635492
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_144
timestamp 1624635492
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14536 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1624635492
transform -1 0 17112 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_162
timestamp 1624635492
transform 1 0 16008 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1624635492
transform -1 0 18584 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_174
timestamp 1624635492
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_178
timestamp 1624635492
transform 1 0 17480 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1624635492
transform 1 0 18768 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20148 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624635492
transform 1 0 19504 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_190
timestamp 1624635492
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_195
timestamp 1624635492
transform 1 0 19044 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_199
timestamp 1624635492
transform 1 0 19412 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_201
timestamp 1624635492
transform 1 0 19596 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1624635492
transform 1 0 20148 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1624635492
transform -1 0 20884 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform 1 0 21068 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_211
timestamp 1624635492
transform 1 0 20516 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1624635492
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1624635492
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 3220 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3588 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1624635492
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_15
timestamp 1624635492
transform 1 0 2484 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1624635492
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_30
timestamp 1624635492
transform 1 0 3864 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_23
timestamp 1624635492
transform 1 0 3220 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1624635492
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624635492
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_36
timestamp 1624635492
transform 1 0 4416 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_36
timestamp 1624635492
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1624635492
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 4508 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_40
timestamp 1624635492
transform 1 0 4784 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4508 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624635492
transform 1 0 6348 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_53
timestamp 1624635492
transform 1 0 5980 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_58
timestamp 1624635492
transform 1 0 6440 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_52
timestamp 1624635492
transform 1 0 5888 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7268 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1624635492
transform -1 0 8188 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_66
timestamp 1624635492
transform 1 0 7176 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_83
timestamp 1624635492
transform 1 0 8740 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_64
timestamp 1624635492
transform 1 0 6992 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_77
timestamp 1624635492
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_81
timestamp 1624635492
transform 1 0 8556 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_85
timestamp 1624635492
transform 1 0 8924 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624635492
transform 1 0 9016 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1624635492
transform -1 0 9752 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_99
timestamp 1624635492
transform 1 0 10212 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_104
timestamp 1624635492
transform 1 0 10672 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_99
timestamp 1624635492
transform 1 0 10212 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_94
timestamp 1624635492
transform 1 0 9752 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 10396 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1624635492
transform 1 0 9936 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_87
timestamp 1624635492
transform 1 0 9108 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_107
timestamp 1624635492
transform 1 0 10948 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_112
timestamp 1624635492
transform 1 0 11408 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624635492
transform 1 0 11592 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12052 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_119
timestamp 1624635492
transform 1 0 12052 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_121
timestamp 1624635492
transform 1 0 12236 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_115
timestamp 1624635492
transform 1 0 11684 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13064 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1624635492
transform -1 0 12236 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12420 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14904 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624635492
transform 1 0 14260 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_139
timestamp 1624635492
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_130
timestamp 1624635492
transform 1 0 13064 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_142
timestamp 1624635492
transform 1 0 14168 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_144
timestamp 1624635492
transform 1 0 14352 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1624635492
transform 1 0 15732 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15180 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1624635492
transform -1 0 15548 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1624635492
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_157
timestamp 1624635492
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_162
timestamp 1624635492
transform 1 0 16008 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624635492
transform 1 0 16836 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_169
timestamp 1624635492
transform 1 0 16652 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_172
timestamp 1624635492
transform 1 0 16928 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_184
timestamp 1624635492
transform 1 0 18032 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_174
timestamp 1624635492
transform 1 0 17112 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_186
timestamp 1624635492
transform 1 0 18216 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_194
timestamp 1624635492
transform 1 0 18952 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_194
timestamp 1624635492
transform 1 0 18952 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_190
timestamp 1624635492
transform 1 0 18584 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19320 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18952 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_201
timestamp 1624635492
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_198
timestamp 1624635492
transform 1 0 19320 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_205
timestamp 1624635492
transform 1 0 19964 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624635492
transform 1 0 19504 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 20056 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19964 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_206
timestamp 1624635492
transform 1 0 20056 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1624635492
transform -1 0 20424 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1624635492
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1624635492
transform 1 0 20608 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1624635492
transform -1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1624635492
transform 1 0 20884 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1624635492
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform 1 0 21068 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform 1 0 21068 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1624635492
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1624635492
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output52
timestamp 1624635492
transform -1 0 1932 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1624635492
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_9
timestamp 1624635492
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1624635492
transform 1 0 3128 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 4140 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_21
timestamp 1624635492
transform 1 0 3036 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_31
timestamp 1624635492
transform 1 0 3956 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_35
timestamp 1624635492
transform 1 0 4324 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1624635492
transform -1 0 7636 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624635492
transform 1 0 6348 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 5888 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_47
timestamp 1624635492
transform 1 0 5428 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_52
timestamp 1624635492
transform 1 0 5888 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_56
timestamp 1624635492
transform 1 0 6256 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1624635492
transform 1 0 6440 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_71
timestamp 1624635492
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_75
timestamp 1624635492
transform 1 0 8004 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10396 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_87
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1624635492
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1624635492
transform 1 0 10396 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624635492
transform 1 0 11592 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 12052 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_105
timestamp 1624635492
transform 1 0 10764 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_113
timestamp 1624635492
transform 1 0 11500 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_115
timestamp 1624635492
transform 1 0 11684 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1624635492
transform 1 0 12236 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_133
timestamp 1624635492
transform 1 0 13340 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_145
timestamp 1624635492
transform 1 0 14444 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_157
timestamp 1624635492
transform 1 0 15548 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17112 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624635492
transform 1 0 16836 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_169
timestamp 1624635492
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_172
timestamp 1624635492
transform 1 0 16928 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1624635492
transform -1 0 20332 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19872 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1624635492
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1624635492
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_199
timestamp 1624635492
transform 1 0 19412 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_204
timestamp 1624635492
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform 1 0 21068 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform 1 0 20516 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_209
timestamp 1624635492
transform 1 0 20332 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1624635492
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1624635492
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1624635492
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1624635492
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624635492
transform 1 0 3772 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_27
timestamp 1624635492
transform 1 0 3588 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_30
timestamp 1624635492
transform 1 0 3864 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 5244 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_42
timestamp 1624635492
transform 1 0 4968 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_61
timestamp 1624635492
transform 1 0 6716 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1624635492
transform 1 0 6900 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_72
timestamp 1624635492
transform 1 0 7728 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9292 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624635492
transform 1 0 9016 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_84
timestamp 1624635492
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_87
timestamp 1624635492
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1624635492
transform 1 0 11960 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11776 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_105
timestamp 1624635492
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_116
timestamp 1624635492
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_121
timestamp 1624635492
transform 1 0 12236 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_125
timestamp 1624635492
transform 1 0 12604 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1624635492
transform -1 0 13892 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624635492
transform 1 0 14260 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_128
timestamp 1624635492
transform 1 0 12880 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_139
timestamp 1624635492
transform 1 0 13892 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_144
timestamp 1624635492
transform 1 0 14352 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15548 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_29_156
timestamp 1624635492
transform 1 0 15456 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1624635492
transform -1 0 19044 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_173
timestamp 1624635492
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1624635492
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1624635492
transform -1 0 20424 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624635492
transform 1 0 19504 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform -1 0 19780 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_195
timestamp 1624635492
transform 1 0 19044 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_199
timestamp 1624635492
transform 1 0 19412 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_203
timestamp 1624635492
transform 1 0 19780 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1624635492
transform -1 0 20884 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output54
timestamp 1624635492
transform 1 0 21068 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1624635492
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1624635492
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1624635492
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 2300 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1624635492
transform 1 0 1380 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1624635492
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4232 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_29
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_33
timestamp 1624635492
transform 1 0 4140 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1624635492
transform 1 0 5244 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1624635492
transform -1 0 6992 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624635492
transform 1 0 6348 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 5888 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_43
timestamp 1624635492
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_48
timestamp 1624635492
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_52
timestamp 1624635492
transform 1 0 5888 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_56
timestamp 1624635492
transform 1 0 6256 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_58
timestamp 1624635492
transform 1 0 6440 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 7176 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 8188 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_64
timestamp 1624635492
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_69
timestamp 1624635492
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_73
timestamp 1624635492
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1624635492
transform 1 0 8188 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1624635492
transform 1 0 8740 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9936 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_86
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_94
timestamp 1624635492
transform 1 0 9752 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12696 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624635492
transform 1 0 11592 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_112
timestamp 1624635492
transform 1 0 11408 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1624635492
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1624635492
transform -1 0 13156 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 13340 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_126
timestamp 1624635492
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_131
timestamp 1624635492
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 16652 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 15088 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_149
timestamp 1624635492
transform 1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1624635492
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17572 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 18308 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624635492
transform 1 0 16836 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_169
timestamp 1624635492
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1624635492
transform 1 0 16928 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 1624635492
transform 1 0 17572 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_183
timestamp 1624635492
transform 1 0 17940 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_187
timestamp 1624635492
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1624635492
transform 1 0 18492 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1624635492
transform 1 0 19504 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1624635492
transform 1 0 19044 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform 1 0 19964 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_192
timestamp 1624635492
transform 1 0 18768 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_198
timestamp 1624635492
transform 1 0 19320 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_203
timestamp 1624635492
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output55
timestamp 1624635492
transform 1 0 21068 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform 1 0 20516 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_209
timestamp 1624635492
transform 1 0 20332 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1624635492
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1624635492
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1624635492
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_15
timestamp 1624635492
transform 1 0 2484 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 4048 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624635492
transform 1 0 3772 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 3588 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 1624635492
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_27
timestamp 1624635492
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_30
timestamp 1624635492
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 5888 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_31_48
timestamp 1624635492
transform 1 0 5520 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1624635492
transform -1 0 8832 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 7728 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_68
timestamp 1624635492
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_72
timestamp 1624635492
transform 1 0 7728 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1624635492
transform -1 0 10120 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624635492
transform 1 0 9016 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_84
timestamp 1624635492
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_87
timestamp 1624635492
transform 1 0 9108 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_98
timestamp 1624635492
transform 1 0 10120 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_104
timestamp 1624635492
transform 1 0 10672 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10764 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_121
timestamp 1624635492
transform 1 0 12236 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624635492
transform 1 0 14260 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_139
timestamp 1624635492
transform 1 0 13892 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1624635492
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14536 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1624635492
transform -1 0 17020 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_162
timestamp 1624635492
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1624635492
transform -1 0 18400 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform -1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_173
timestamp 1624635492
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_179
timestamp 1624635492
transform 1 0 17572 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1624635492
transform -1 0 19320 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1624635492
transform 1 0 18584 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624635492
transform 1 0 19504 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform 1 0 19872 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_188
timestamp 1624635492
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_193
timestamp 1624635492
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_198
timestamp 1624635492
transform 1 0 19320 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_201
timestamp 1624635492
transform 1 0 19596 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_208
timestamp 1624635492
transform 1 0 20240 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output56
timestamp 1624635492
transform 1 0 21068 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform -1 0 20792 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_214
timestamp 1624635492
transform 1 0 20792 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1624635492
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 2576 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 3036 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 1564 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_5
timestamp 1624635492
transform 1 0 1564 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1624635492
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_16
timestamp 1624635492
transform 1 0 2576 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1624635492
transform -1 0 4968 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 3956 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_21
timestamp 1624635492
transform 1 0 3036 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1624635492
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_31
timestamp 1624635492
transform 1 0 3956 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_42
timestamp 1624635492
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 5336 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_46
timestamp 1624635492
transform 1 0 5336 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 5704 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_50
timestamp 1624635492
transform 1 0 5704 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1624635492
transform -1 0 6164 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_55
timestamp 1624635492
transform 1 0 6164 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624635492
transform 1 0 6348 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_58
timestamp 1624635492
transform 1 0 6440 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1624635492
transform 1 0 6624 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7544 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 7268 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_63
timestamp 1624635492
transform 1 0 6900 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_67
timestamp 1624635492
transform 1 0 7268 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1624635492
transform -1 0 9476 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 10212 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 10580 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_86
timestamp 1624635492
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1624635492
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_95
timestamp 1624635492
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_99
timestamp 1624635492
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_103
timestamp 1624635492
transform 1 0 10580 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_107
timestamp 1624635492
transform 1 0 10948 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 10948 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_111
timestamp 1624635492
transform 1 0 11316 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_115
timestamp 1624635492
transform 1 0 11684 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624635492
transform 1 0 11592 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1624635492
transform 1 0 11868 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_120
timestamp 1624635492
transform 1 0 12144 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 12512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_124
timestamp 1624635492
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15088 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output84_A
timestamp 1624635492
transform 1 0 13064 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_128
timestamp 1624635492
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1624635492
transform 1 0 13248 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_140
timestamp 1624635492
transform 1 0 13984 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1624635492
transform -1 0 16652 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform -1 0 15640 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform -1 0 16192 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_152
timestamp 1624635492
transform 1 0 15088 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_158
timestamp 1624635492
transform 1 0 15640 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_164
timestamp 1624635492
transform 1 0 16192 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624635492
transform 1 0 16836 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform -1 0 17480 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform -1 0 18032 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_169
timestamp 1624635492
transform 1 0 16652 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_172
timestamp 1624635492
transform 1 0 16928 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_178
timestamp 1624635492
transform 1 0 17480 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1624635492
transform 1 0 18032 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 19596 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform -1 0 20148 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_188
timestamp 1624635492
transform 1 0 18400 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_201
timestamp 1624635492
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_207
timestamp 1624635492
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output57
timestamp 1624635492
transform 1 0 21068 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform -1 0 20700 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_213
timestamp 1624635492
transform 1 0 20700 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1624635492
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1624635492
transform 1 0 2116 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1624635492
transform 1 0 2576 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1624635492
transform 1 0 1564 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1624635492
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_9
timestamp 1624635492
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_14
timestamp 1624635492
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_19
timestamp 1624635492
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624635492
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1624635492
transform 1 0 3036 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1624635492
transform 1 0 4048 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1624635492
transform -1 0 4784 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_24
timestamp 1624635492
transform 1 0 3312 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_28
timestamp 1624635492
transform 1 0 3680 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_30
timestamp 1624635492
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_35
timestamp 1624635492
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_40
timestamp 1624635492
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624635492
transform 1 0 6440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1624635492
transform 1 0 6716 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1624635492
transform 1 0 4968 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1624635492
transform 1 0 5428 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1624635492
transform -1 0 6164 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_45
timestamp 1624635492
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_50
timestamp 1624635492
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_55
timestamp 1624635492
transform 1 0 6164 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1624635492
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1624635492
transform 1 0 7176 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1624635492
transform -1 0 7912 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1624635492
transform 1 0 8096 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1624635492
transform 1 0 8648 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_64
timestamp 1624635492
transform 1 0 6992 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1624635492
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_74
timestamp 1624635492
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_79
timestamp 1624635492
transform 1 0 8372 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624635492
transform 1 0 9108 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1624635492
transform -1 0 9660 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1624635492
transform -1 0 10120 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1624635492
transform -1 0 10580 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_85
timestamp 1624635492
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_88
timestamp 1624635492
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_93
timestamp 1624635492
transform 1 0 9660 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_98
timestamp 1624635492
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_103
timestamp 1624635492
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624635492
transform 1 0 11776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1624635492
transform -1 0 11040 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform -1 0 12420 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform -1 0 12972 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform 1 0 11224 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_108
timestamp 1624635492
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1624635492
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1624635492
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_123
timestamp 1624635492
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624635492
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform -1 0 13524 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform -1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_129
timestamp 1624635492
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1624635492
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_141
timestamp 1624635492
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform 1 0 16008 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform 1 0 15456 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform 1 0 14904 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1624635492
transform -1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_148
timestamp 1624635492
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_154
timestamp 1624635492
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_160
timestamp 1624635492
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1624635492
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624635492
transform 1 0 17112 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1624635492
transform 1 0 18124 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform 1 0 16560 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_172
timestamp 1624635492
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_175
timestamp 1624635492
transform 1 0 17204 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_183
timestamp 1624635492
transform 1 0 17940 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1624635492
transform 1 0 20056 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624635492
transform 1 0 19780 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output60
timestamp 1624635492
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1624635492
transform 1 0 18676 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_189
timestamp 1624635492
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_195
timestamp 1624635492
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1624635492
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1624635492
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output58
timestamp 1624635492
transform 1 0 21068 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output59
timestamp 1624635492
transform 1 0 20516 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1624635492
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1624635492
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1624635492
transform 1 0 21436 0 1 20128
box -38 -48 222 592
<< labels >>
rlabel metal3 s 0 5720 800 5840 6 ccff_head
port 0 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 ccff_tail
port 1 nsew signal tristate
rlabel metal3 s 22200 4224 23000 4344 6 chanx_right_in[0]
port 2 nsew signal input
rlabel metal3 s 22200 8848 23000 8968 6 chanx_right_in[10]
port 3 nsew signal input
rlabel metal3 s 22200 9256 23000 9376 6 chanx_right_in[11]
port 4 nsew signal input
rlabel metal3 s 22200 9664 23000 9784 6 chanx_right_in[12]
port 5 nsew signal input
rlabel metal3 s 22200 10208 23000 10328 6 chanx_right_in[13]
port 6 nsew signal input
rlabel metal3 s 22200 10616 23000 10736 6 chanx_right_in[14]
port 7 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[15]
port 8 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[16]
port 9 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_in[17]
port 10 nsew signal input
rlabel metal3 s 22200 12520 23000 12640 6 chanx_right_in[18]
port 11 nsew signal input
rlabel metal3 s 22200 12928 23000 13048 6 chanx_right_in[19]
port 12 nsew signal input
rlabel metal3 s 22200 4632 23000 4752 6 chanx_right_in[1]
port 13 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[2]
port 14 nsew signal input
rlabel metal3 s 22200 5584 23000 5704 6 chanx_right_in[3]
port 15 nsew signal input
rlabel metal3 s 22200 5992 23000 6112 6 chanx_right_in[4]
port 16 nsew signal input
rlabel metal3 s 22200 6536 23000 6656 6 chanx_right_in[5]
port 17 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[6]
port 18 nsew signal input
rlabel metal3 s 22200 7488 23000 7608 6 chanx_right_in[7]
port 19 nsew signal input
rlabel metal3 s 22200 7896 23000 8016 6 chanx_right_in[8]
port 20 nsew signal input
rlabel metal3 s 22200 8304 23000 8424 6 chanx_right_in[9]
port 21 nsew signal input
rlabel metal3 s 22200 13472 23000 13592 6 chanx_right_out[0]
port 22 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[10]
port 23 nsew signal tristate
rlabel metal3 s 22200 18504 23000 18624 6 chanx_right_out[11]
port 24 nsew signal tristate
rlabel metal3 s 22200 18912 23000 19032 6 chanx_right_out[12]
port 25 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[13]
port 26 nsew signal tristate
rlabel metal3 s 22200 19864 23000 19984 6 chanx_right_out[14]
port 27 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[15]
port 28 nsew signal tristate
rlabel metal3 s 22200 20816 23000 20936 6 chanx_right_out[16]
port 29 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[17]
port 30 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[18]
port 31 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[19]
port 32 nsew signal tristate
rlabel metal3 s 22200 13880 23000 14000 6 chanx_right_out[1]
port 33 nsew signal tristate
rlabel metal3 s 22200 14288 23000 14408 6 chanx_right_out[2]
port 34 nsew signal tristate
rlabel metal3 s 22200 14832 23000 14952 6 chanx_right_out[3]
port 35 nsew signal tristate
rlabel metal3 s 22200 15240 23000 15360 6 chanx_right_out[4]
port 36 nsew signal tristate
rlabel metal3 s 22200 15648 23000 15768 6 chanx_right_out[5]
port 37 nsew signal tristate
rlabel metal3 s 22200 16192 23000 16312 6 chanx_right_out[6]
port 38 nsew signal tristate
rlabel metal3 s 22200 16600 23000 16720 6 chanx_right_out[7]
port 39 nsew signal tristate
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[8]
port 40 nsew signal tristate
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[9]
port 41 nsew signal tristate
rlabel metal2 s 846 22200 902 23000 6 chany_top_in[0]
port 42 nsew signal input
rlabel metal2 s 6458 22200 6514 23000 6 chany_top_in[10]
port 43 nsew signal input
rlabel metal2 s 7010 22200 7066 23000 6 chany_top_in[11]
port 44 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[12]
port 45 nsew signal input
rlabel metal2 s 8114 22200 8170 23000 6 chany_top_in[13]
port 46 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[14]
port 47 nsew signal input
rlabel metal2 s 9218 22200 9274 23000 6 chany_top_in[15]
port 48 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[16]
port 49 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[17]
port 50 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_in[18]
port 51 nsew signal input
rlabel metal2 s 11426 22200 11482 23000 6 chany_top_in[19]
port 52 nsew signal input
rlabel metal2 s 1398 22200 1454 23000 6 chany_top_in[1]
port 53 nsew signal input
rlabel metal2 s 1950 22200 2006 23000 6 chany_top_in[2]
port 54 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 chany_top_in[3]
port 55 nsew signal input
rlabel metal2 s 3054 22200 3110 23000 6 chany_top_in[4]
port 56 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 chany_top_in[5]
port 57 nsew signal input
rlabel metal2 s 4158 22200 4214 23000 6 chany_top_in[6]
port 58 nsew signal input
rlabel metal2 s 4710 22200 4766 23000 6 chany_top_in[7]
port 59 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[8]
port 60 nsew signal input
rlabel metal2 s 5814 22200 5870 23000 6 chany_top_in[9]
port 61 nsew signal input
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_out[0]
port 62 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 63 nsew signal tristate
rlabel metal2 s 18234 22200 18290 23000 6 chany_top_out[11]
port 64 nsew signal tristate
rlabel metal2 s 18786 22200 18842 23000 6 chany_top_out[12]
port 65 nsew signal tristate
rlabel metal2 s 19338 22200 19394 23000 6 chany_top_out[13]
port 66 nsew signal tristate
rlabel metal2 s 19890 22200 19946 23000 6 chany_top_out[14]
port 67 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[15]
port 68 nsew signal tristate
rlabel metal2 s 20994 22200 21050 23000 6 chany_top_out[16]
port 69 nsew signal tristate
rlabel metal2 s 21546 22200 21602 23000 6 chany_top_out[17]
port 70 nsew signal tristate
rlabel metal2 s 22098 22200 22154 23000 6 chany_top_out[18]
port 71 nsew signal tristate
rlabel metal2 s 22650 22200 22706 23000 6 chany_top_out[19]
port 72 nsew signal tristate
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_out[1]
port 73 nsew signal tristate
rlabel metal2 s 13174 22200 13230 23000 6 chany_top_out[2]
port 74 nsew signal tristate
rlabel metal2 s 13726 22200 13782 23000 6 chany_top_out[3]
port 75 nsew signal tristate
rlabel metal2 s 14278 22200 14334 23000 6 chany_top_out[4]
port 76 nsew signal tristate
rlabel metal2 s 14830 22200 14886 23000 6 chany_top_out[5]
port 77 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[6]
port 78 nsew signal tristate
rlabel metal2 s 15934 22200 15990 23000 6 chany_top_out[7]
port 79 nsew signal tristate
rlabel metal2 s 16486 22200 16542 23000 6 chany_top_out[8]
port 80 nsew signal tristate
rlabel metal2 s 17038 22200 17094 23000 6 chany_top_out[9]
port 81 nsew signal tristate
rlabel metal3 s 22200 22584 23000 22704 6 prog_clk_0_E_in
port 82 nsew signal input
rlabel metal3 s 22200 2320 23000 2440 6 right_bottom_grid_pin_11_
port 83 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_13_
port 84 nsew signal input
rlabel metal3 s 22200 3272 23000 3392 6 right_bottom_grid_pin_15_
port 85 nsew signal input
rlabel metal3 s 22200 3816 23000 3936 6 right_bottom_grid_pin_17_
port 86 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_1_
port 87 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_3_
port 88 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_5_
port 89 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_7_
port 90 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_9_
port 91 nsew signal input
rlabel metal2 s 294 22200 350 23000 6 top_left_grid_pin_1_
port 92 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 93 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 94 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 95 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 96 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 97 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
