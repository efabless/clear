magic
tech sky130A
magscale 1 2
timestamp 1656405897
<< viali >>
rect 2053 20553 2087 20587
rect 5917 20553 5951 20587
rect 9873 20553 9907 20587
rect 11069 20553 11103 20587
rect 16313 20553 16347 20587
rect 17509 20553 17543 20587
rect 11805 20485 11839 20519
rect 1685 20417 1719 20451
rect 2237 20417 2271 20451
rect 2697 20417 2731 20451
rect 2973 20417 3007 20451
rect 4905 20417 4939 20451
rect 6377 20417 6411 20451
rect 6653 20417 6687 20451
rect 7941 20417 7975 20451
rect 9321 20417 9355 20451
rect 9965 20417 9999 20451
rect 12541 20417 12575 20451
rect 16129 20417 16163 20451
rect 16681 20417 16715 20451
rect 17325 20417 17359 20451
rect 19717 20417 19751 20451
rect 19993 20417 20027 20451
rect 20545 20417 20579 20451
rect 21097 20417 21131 20451
rect 4537 20349 4571 20383
rect 7665 20349 7699 20383
rect 7849 20349 7883 20383
rect 9781 20349 9815 20383
rect 13461 20349 13495 20383
rect 15485 20349 15519 20383
rect 18245 20349 18279 20383
rect 18889 20349 18923 20383
rect 12909 20281 12943 20315
rect 16865 20281 16899 20315
rect 1501 20213 1535 20247
rect 2513 20213 2547 20247
rect 3157 20213 3191 20247
rect 3893 20213 3927 20247
rect 4169 20213 4203 20247
rect 5273 20213 5307 20247
rect 8309 20213 8343 20247
rect 10333 20213 10367 20247
rect 10793 20213 10827 20247
rect 14381 20213 14415 20247
rect 14841 20213 14875 20247
rect 17877 20213 17911 20247
rect 19533 20213 19567 20247
rect 20177 20213 20211 20247
rect 20729 20213 20763 20247
rect 21281 20213 21315 20247
rect 2513 20009 2547 20043
rect 2973 20009 3007 20043
rect 6009 20009 6043 20043
rect 19993 20009 20027 20043
rect 20729 20009 20763 20043
rect 2053 19941 2087 19975
rect 14749 19941 14783 19975
rect 3985 19873 4019 19907
rect 8033 19873 8067 19907
rect 10057 19873 10091 19907
rect 10149 19873 10183 19907
rect 11069 19873 11103 19907
rect 13093 19873 13127 19907
rect 13277 19873 13311 19907
rect 15209 19873 15243 19907
rect 16589 19873 16623 19907
rect 17601 19873 17635 19907
rect 19441 19873 19475 19907
rect 1685 19805 1719 19839
rect 2237 19805 2271 19839
rect 2697 19805 2731 19839
rect 3157 19805 3191 19839
rect 4077 19805 4111 19839
rect 8125 19805 8159 19839
rect 9505 19805 9539 19839
rect 10241 19805 10275 19839
rect 12081 19805 12115 19839
rect 12449 19805 12483 19839
rect 14565 19805 14599 19839
rect 15393 19805 15427 19839
rect 18705 19805 18739 19839
rect 20545 19805 20579 19839
rect 21097 19805 21131 19839
rect 4169 19737 4203 19771
rect 4813 19737 4847 19771
rect 6837 19737 6871 19771
rect 8217 19737 8251 19771
rect 8953 19737 8987 19771
rect 13369 19737 13403 19771
rect 14105 19737 14139 19771
rect 15301 19737 15335 19771
rect 16497 19737 16531 19771
rect 17417 19737 17451 19771
rect 18061 19737 18095 19771
rect 1501 19669 1535 19703
rect 4537 19669 4571 19703
rect 5457 19669 5491 19703
rect 6285 19669 6319 19703
rect 7113 19669 7147 19703
rect 7573 19669 7607 19703
rect 8585 19669 8619 19703
rect 10609 19669 10643 19703
rect 11161 19669 11195 19703
rect 11253 19669 11287 19703
rect 11621 19669 11655 19703
rect 13737 19669 13771 19703
rect 15761 19669 15795 19703
rect 16037 19669 16071 19703
rect 16405 19669 16439 19703
rect 17049 19669 17083 19703
rect 17509 19669 17543 19703
rect 18521 19669 18555 19703
rect 19533 19669 19567 19703
rect 19625 19669 19659 19703
rect 21281 19669 21315 19703
rect 3985 19465 4019 19499
rect 5365 19465 5399 19499
rect 7757 19465 7791 19499
rect 10609 19465 10643 19499
rect 13093 19465 13127 19499
rect 13461 19465 13495 19499
rect 15209 19465 15243 19499
rect 16037 19465 16071 19499
rect 17417 19465 17451 19499
rect 18245 19465 18279 19499
rect 18337 19465 18371 19499
rect 19625 19465 19659 19499
rect 19993 19465 20027 19499
rect 20729 19465 20763 19499
rect 5457 19397 5491 19431
rect 9965 19397 9999 19431
rect 10517 19397 10551 19431
rect 16957 19397 16991 19431
rect 1685 19329 1719 19363
rect 2237 19329 2271 19363
rect 2513 19329 2547 19363
rect 3525 19329 3559 19363
rect 3617 19329 3651 19363
rect 7389 19329 7423 19363
rect 11805 19329 11839 19363
rect 11897 19329 11931 19363
rect 12541 19329 12575 19363
rect 17049 19329 17083 19363
rect 20545 19329 20579 19363
rect 21097 19329 21131 19363
rect 3341 19261 3375 19295
rect 5641 19261 5675 19295
rect 7205 19261 7239 19295
rect 7297 19261 7331 19295
rect 8401 19261 8435 19295
rect 10425 19261 10459 19295
rect 11713 19261 11747 19295
rect 13553 19261 13587 19295
rect 13645 19261 13679 19295
rect 14197 19261 14231 19295
rect 15025 19261 15059 19295
rect 15117 19261 15151 19295
rect 16865 19261 16899 19295
rect 18429 19261 18463 19295
rect 19441 19261 19475 19295
rect 19533 19261 19567 19295
rect 2053 19193 2087 19227
rect 4353 19193 4387 19227
rect 4721 19193 4755 19227
rect 8953 19193 8987 19227
rect 12265 19193 12299 19227
rect 14565 19193 14599 19227
rect 15577 19193 15611 19227
rect 1501 19125 1535 19159
rect 2697 19125 2731 19159
rect 4997 19125 5031 19159
rect 6745 19125 6779 19159
rect 8033 19125 8067 19159
rect 9229 19125 9263 19159
rect 10977 19125 11011 19159
rect 12725 19125 12759 19159
rect 17877 19125 17911 19159
rect 18889 19125 18923 19159
rect 21281 19125 21315 19159
rect 2421 18921 2455 18955
rect 4537 18921 4571 18955
rect 11713 18921 11747 18955
rect 12449 18921 12483 18955
rect 15485 18921 15519 18955
rect 18889 18921 18923 18955
rect 2881 18853 2915 18887
rect 3893 18853 3927 18887
rect 5641 18853 5675 18887
rect 9689 18853 9723 18887
rect 17049 18853 17083 18887
rect 17509 18853 17543 18887
rect 19717 18853 19751 18887
rect 5181 18785 5215 18819
rect 8033 18785 8067 18819
rect 10609 18785 10643 18819
rect 14933 18785 14967 18819
rect 16313 18785 16347 18819
rect 1685 18717 1719 18751
rect 2145 18717 2179 18751
rect 2605 18717 2639 18751
rect 3065 18717 3099 18751
rect 4905 18717 4939 18751
rect 6009 18717 6043 18751
rect 8217 18717 8251 18751
rect 13093 18717 13127 18751
rect 16865 18717 16899 18751
rect 17325 18717 17359 18751
rect 17785 18717 17819 18751
rect 18429 18717 18463 18751
rect 18705 18717 18739 18751
rect 19533 18717 19567 18751
rect 20177 18717 20211 18751
rect 20637 18717 20671 18751
rect 21097 18717 21131 18751
rect 6285 18649 6319 18683
rect 8125 18649 8159 18683
rect 9321 18649 9355 18683
rect 15117 18649 15151 18683
rect 15945 18649 15979 18683
rect 1501 18581 1535 18615
rect 1961 18581 1995 18615
rect 3341 18581 3375 18615
rect 4261 18581 4295 18615
rect 4997 18581 5031 18615
rect 6653 18581 6687 18615
rect 7021 18581 7055 18615
rect 7481 18581 7515 18615
rect 8585 18581 8619 18615
rect 8953 18581 8987 18615
rect 11345 18581 11379 18615
rect 12725 18581 12759 18615
rect 13645 18581 13679 18615
rect 14381 18581 14415 18615
rect 15025 18581 15059 18615
rect 17969 18581 18003 18615
rect 18245 18581 18279 18615
rect 19993 18581 20027 18615
rect 20453 18581 20487 18615
rect 21281 18581 21315 18615
rect 2145 18377 2179 18411
rect 2421 18377 2455 18411
rect 2881 18377 2915 18411
rect 4721 18377 4755 18411
rect 6929 18377 6963 18411
rect 7665 18377 7699 18411
rect 9965 18377 9999 18411
rect 10609 18377 10643 18411
rect 11989 18377 12023 18411
rect 12817 18377 12851 18411
rect 13461 18377 13495 18411
rect 15117 18377 15151 18411
rect 15485 18377 15519 18411
rect 16313 18377 16347 18411
rect 18613 18377 18647 18411
rect 19901 18377 19935 18411
rect 4629 18309 4663 18343
rect 8033 18309 8067 18343
rect 9045 18309 9079 18343
rect 14381 18309 14415 18343
rect 15577 18309 15611 18343
rect 1685 18241 1719 18275
rect 1961 18241 1995 18275
rect 2605 18241 2639 18275
rect 3065 18241 3099 18275
rect 6837 18241 6871 18275
rect 12449 18241 12483 18275
rect 14473 18241 14507 18275
rect 16129 18241 16163 18275
rect 17325 18241 17359 18275
rect 18245 18241 18279 18275
rect 18889 18241 18923 18275
rect 19257 18241 19291 18275
rect 19717 18241 19751 18275
rect 20177 18241 20211 18275
rect 20821 18241 20855 18275
rect 21097 18241 21131 18275
rect 4537 18173 4571 18207
rect 7113 18173 7147 18207
rect 8125 18173 8159 18207
rect 8309 18173 8343 18207
rect 9689 18173 9723 18207
rect 9873 18173 9907 18207
rect 13185 18173 13219 18207
rect 13369 18173 13403 18207
rect 14197 18173 14231 18207
rect 15669 18173 15703 18207
rect 17049 18173 17083 18207
rect 18061 18173 18095 18207
rect 18153 18173 18187 18207
rect 5089 18105 5123 18139
rect 10333 18105 10367 18139
rect 14841 18105 14875 18139
rect 19441 18105 19475 18139
rect 20361 18105 20395 18139
rect 1501 18037 1535 18071
rect 3341 18037 3375 18071
rect 3801 18037 3835 18071
rect 5365 18037 5399 18071
rect 5733 18037 5767 18071
rect 6469 18037 6503 18071
rect 8677 18037 8711 18071
rect 13829 18037 13863 18071
rect 20637 18037 20671 18071
rect 21281 18037 21315 18071
rect 2973 17833 3007 17867
rect 6837 17833 6871 17867
rect 7481 17833 7515 17867
rect 7849 17833 7883 17867
rect 18429 17833 18463 17867
rect 19349 17833 19383 17867
rect 16589 17765 16623 17799
rect 4629 17697 4663 17731
rect 8493 17697 8527 17731
rect 10333 17697 10367 17731
rect 11069 17697 11103 17731
rect 11897 17697 11931 17731
rect 12725 17697 12759 17731
rect 15669 17697 15703 17731
rect 17141 17697 17175 17731
rect 19901 17697 19935 17731
rect 1685 17629 1719 17663
rect 2237 17629 2271 17663
rect 2697 17629 2731 17663
rect 3157 17629 3191 17663
rect 5273 17629 5307 17663
rect 5733 17629 5767 17663
rect 8217 17629 8251 17663
rect 9413 17629 9447 17663
rect 10057 17629 10091 17663
rect 11345 17629 11379 17663
rect 15025 17629 15059 17663
rect 17325 17629 17359 17663
rect 18245 17629 18279 17663
rect 18705 17629 18739 17663
rect 20545 17629 20579 17663
rect 21097 17629 21131 17663
rect 4353 17561 4387 17595
rect 9045 17561 9079 17595
rect 12633 17561 12667 17595
rect 15853 17561 15887 17595
rect 19717 17561 19751 17595
rect 1501 17493 1535 17527
rect 2053 17493 2087 17527
rect 2513 17493 2547 17527
rect 3985 17493 4019 17527
rect 4445 17493 4479 17527
rect 6101 17493 6135 17527
rect 7113 17493 7147 17527
rect 8309 17493 8343 17527
rect 9689 17493 9723 17527
rect 10149 17493 10183 17527
rect 12173 17493 12207 17527
rect 12541 17493 12575 17527
rect 13185 17493 13219 17527
rect 13645 17493 13679 17527
rect 14381 17493 14415 17527
rect 14749 17493 14783 17527
rect 15209 17493 15243 17527
rect 15761 17493 15795 17527
rect 16221 17493 16255 17527
rect 17233 17493 17267 17527
rect 17693 17493 17727 17527
rect 18889 17493 18923 17527
rect 19809 17493 19843 17527
rect 20729 17493 20763 17527
rect 21281 17493 21315 17527
rect 2329 17289 2363 17323
rect 2789 17289 2823 17323
rect 3341 17289 3375 17323
rect 5641 17289 5675 17323
rect 5733 17289 5767 17323
rect 6745 17289 6779 17323
rect 7573 17289 7607 17323
rect 7941 17289 7975 17323
rect 9229 17289 9263 17323
rect 10333 17289 10367 17323
rect 10425 17289 10459 17323
rect 13185 17289 13219 17323
rect 13829 17289 13863 17323
rect 14473 17289 14507 17323
rect 15577 17289 15611 17323
rect 17693 17289 17727 17323
rect 19257 17289 19291 17323
rect 8585 17221 8619 17255
rect 9321 17221 9355 17255
rect 13737 17221 13771 17255
rect 1685 17153 1719 17187
rect 2697 17153 2731 17187
rect 3709 17153 3743 17187
rect 6837 17153 6871 17187
rect 12265 17153 12299 17187
rect 12633 17153 12667 17187
rect 14841 17153 14875 17187
rect 15945 17153 15979 17187
rect 16037 17153 16071 17187
rect 18889 17153 18923 17187
rect 19901 17153 19935 17187
rect 20545 17153 20579 17187
rect 21097 17153 21131 17187
rect 2973 17085 3007 17119
rect 3801 17085 3835 17119
rect 3985 17085 4019 17119
rect 4997 17085 5031 17119
rect 5917 17085 5951 17119
rect 6929 17085 6963 17119
rect 8033 17085 8067 17119
rect 8217 17085 8251 17119
rect 9045 17085 9079 17119
rect 10149 17085 10183 17119
rect 11529 17085 11563 17119
rect 13645 17085 13679 17119
rect 14933 17085 14967 17119
rect 15025 17085 15059 17119
rect 16221 17085 16255 17119
rect 17509 17085 17543 17119
rect 17601 17085 17635 17119
rect 18705 17085 18739 17119
rect 18797 17085 18831 17119
rect 19993 17085 20027 17119
rect 20085 17085 20119 17119
rect 6377 17017 6411 17051
rect 9689 17017 9723 17051
rect 11161 17017 11195 17051
rect 16681 17017 16715 17051
rect 19533 17017 19567 17051
rect 1501 16949 1535 16983
rect 2053 16949 2087 16983
rect 4445 16949 4479 16983
rect 5273 16949 5307 16983
rect 10793 16949 10827 16983
rect 14197 16949 14231 16983
rect 18061 16949 18095 16983
rect 20729 16949 20763 16983
rect 21281 16949 21315 16983
rect 4537 16745 4571 16779
rect 6193 16745 6227 16779
rect 16405 16745 16439 16779
rect 17233 16745 17267 16779
rect 18245 16745 18279 16779
rect 19625 16745 19659 16779
rect 6929 16677 6963 16711
rect 9965 16677 9999 16711
rect 4169 16609 4203 16643
rect 4905 16609 4939 16643
rect 7849 16609 7883 16643
rect 9505 16609 9539 16643
rect 10333 16609 10367 16643
rect 10793 16609 10827 16643
rect 11069 16609 11103 16643
rect 12633 16609 12667 16643
rect 13093 16609 13127 16643
rect 13645 16609 13679 16643
rect 14565 16609 14599 16643
rect 15117 16609 15151 16643
rect 16037 16609 16071 16643
rect 16865 16609 16899 16643
rect 17601 16609 17635 16643
rect 17785 16609 17819 16643
rect 20177 16609 20211 16643
rect 21189 16609 21223 16643
rect 1685 16541 1719 16575
rect 2329 16541 2363 16575
rect 2973 16541 3007 16575
rect 3433 16541 3467 16575
rect 5181 16541 5215 16575
rect 7665 16541 7699 16575
rect 9321 16541 9355 16575
rect 11897 16541 11931 16575
rect 12265 16541 12299 16575
rect 18521 16541 18555 16575
rect 21097 16541 21131 16575
rect 6561 16473 6595 16507
rect 7573 16473 7607 16507
rect 15301 16473 15335 16507
rect 17877 16473 17911 16507
rect 1501 16405 1535 16439
rect 2145 16405 2179 16439
rect 2789 16405 2823 16439
rect 3249 16405 3283 16439
rect 5089 16405 5123 16439
rect 5549 16405 5583 16439
rect 7205 16405 7239 16439
rect 8217 16405 8251 16439
rect 8953 16405 8987 16439
rect 9413 16405 9447 16439
rect 15209 16405 15243 16439
rect 15669 16405 15703 16439
rect 18705 16405 18739 16439
rect 19257 16405 19291 16439
rect 19993 16405 20027 16439
rect 20085 16405 20119 16439
rect 20637 16405 20671 16439
rect 21005 16405 21039 16439
rect 2513 16201 2547 16235
rect 3341 16201 3375 16235
rect 5825 16201 5859 16235
rect 7665 16201 7699 16235
rect 8217 16201 8251 16235
rect 8677 16201 8711 16235
rect 11529 16201 11563 16235
rect 11897 16201 11931 16235
rect 12633 16201 12667 16235
rect 15485 16201 15519 16235
rect 17233 16201 17267 16235
rect 18981 16201 19015 16235
rect 20729 16201 20763 16235
rect 3709 16133 3743 16167
rect 5457 16133 5491 16167
rect 7205 16133 7239 16167
rect 13001 16133 13035 16167
rect 15853 16133 15887 16167
rect 16221 16133 16255 16167
rect 17509 16133 17543 16167
rect 19441 16133 19475 16167
rect 1685 16065 1719 16099
rect 2237 16065 2271 16099
rect 2697 16065 2731 16099
rect 3801 16065 3835 16099
rect 7297 16065 7331 16099
rect 8309 16065 8343 16099
rect 14933 16065 14967 16099
rect 16681 16065 16715 16099
rect 18797 16065 18831 16099
rect 19717 16065 19751 16099
rect 20637 16065 20671 16099
rect 3893 15997 3927 16031
rect 6653 15997 6687 16031
rect 7113 15997 7147 16031
rect 8125 15997 8159 16031
rect 14289 15997 14323 16031
rect 20821 15997 20855 16031
rect 2053 15929 2087 15963
rect 4997 15929 5031 15963
rect 9781 15929 9815 15963
rect 10517 15929 10551 15963
rect 13921 15929 13955 15963
rect 18153 15929 18187 15963
rect 18429 15929 18463 15963
rect 20269 15929 20303 15963
rect 1501 15861 1535 15895
rect 2973 15861 3007 15895
rect 4721 15861 4755 15895
rect 8953 15861 8987 15895
rect 9413 15861 9447 15895
rect 10057 15861 10091 15895
rect 10885 15861 10919 15895
rect 12357 15861 12391 15895
rect 13369 15861 13403 15895
rect 14657 15861 14691 15895
rect 19901 15861 19935 15895
rect 21281 15861 21315 15895
rect 2237 15657 2271 15691
rect 2697 15657 2731 15691
rect 6101 15657 6135 15691
rect 9321 15657 9355 15691
rect 11345 15657 11379 15691
rect 11713 15657 11747 15691
rect 17693 15657 17727 15691
rect 3893 15521 3927 15555
rect 5549 15521 5583 15555
rect 6745 15521 6779 15555
rect 7573 15521 7607 15555
rect 7757 15521 7791 15555
rect 8401 15521 8435 15555
rect 13277 15521 13311 15555
rect 18245 15521 18279 15555
rect 1685 15453 1719 15487
rect 2421 15453 2455 15487
rect 2881 15453 2915 15487
rect 4169 15453 4203 15487
rect 6469 15453 6503 15487
rect 7481 15453 7515 15487
rect 10701 15453 10735 15487
rect 10977 15453 11011 15487
rect 16598 15453 16632 15487
rect 16865 15453 16899 15487
rect 18153 15453 18187 15487
rect 18705 15453 18739 15487
rect 19441 15453 19475 15487
rect 19993 15453 20027 15487
rect 20545 15453 20579 15487
rect 21097 15453 21131 15487
rect 5457 15385 5491 15419
rect 8953 15385 8987 15419
rect 10434 15385 10468 15419
rect 13645 15385 13679 15419
rect 14105 15385 14139 15419
rect 14841 15385 14875 15419
rect 1501 15317 1535 15351
rect 3249 15317 3283 15351
rect 4077 15317 4111 15351
rect 4537 15317 4571 15351
rect 4997 15317 5031 15351
rect 5365 15317 5399 15351
rect 6561 15317 6595 15351
rect 7113 15317 7147 15351
rect 12081 15317 12115 15351
rect 12449 15317 12483 15351
rect 12817 15317 12851 15351
rect 14473 15317 14507 15351
rect 15485 15317 15519 15351
rect 17233 15317 17267 15351
rect 18061 15317 18095 15351
rect 19625 15317 19659 15351
rect 20177 15317 20211 15351
rect 20729 15317 20763 15351
rect 21281 15317 21315 15351
rect 1961 15113 1995 15147
rect 2789 15113 2823 15147
rect 3801 15113 3835 15147
rect 4629 15113 4663 15147
rect 11069 15113 11103 15147
rect 11529 15113 11563 15147
rect 12541 15113 12575 15147
rect 12909 15113 12943 15147
rect 19625 15113 19659 15147
rect 9934 15045 9968 15079
rect 1685 14977 1719 15011
rect 2145 14977 2179 15011
rect 5641 14977 5675 15011
rect 7389 14977 7423 15011
rect 8401 14977 8435 15011
rect 9689 14977 9723 15011
rect 14022 14977 14056 15011
rect 14289 14977 14323 15011
rect 15770 14977 15804 15011
rect 16037 14977 16071 15011
rect 16681 14977 16715 15011
rect 18898 14977 18932 15011
rect 19165 14977 19199 15011
rect 20738 14977 20772 15011
rect 21005 14977 21039 15011
rect 21281 14977 21315 15011
rect 2605 14909 2639 14943
rect 2697 14909 2731 14943
rect 4721 14909 4755 14943
rect 4905 14909 4939 14943
rect 5733 14909 5767 14943
rect 5917 14909 5951 14943
rect 7481 14909 7515 14943
rect 7573 14909 7607 14943
rect 3525 14841 3559 14875
rect 5273 14841 5307 14875
rect 6745 14841 6779 14875
rect 8769 14841 8803 14875
rect 1501 14773 1535 14807
rect 3157 14773 3191 14807
rect 4261 14773 4295 14807
rect 7021 14773 7055 14807
rect 8033 14773 8067 14807
rect 9137 14773 9171 14807
rect 11989 14773 12023 14807
rect 14657 14773 14691 14807
rect 17325 14773 17359 14807
rect 17785 14773 17819 14807
rect 10425 14569 10459 14603
rect 10701 14569 10735 14603
rect 14105 14569 14139 14603
rect 15853 14569 15887 14603
rect 19441 14569 19475 14603
rect 3065 14501 3099 14535
rect 7849 14501 7883 14535
rect 4261 14433 4295 14467
rect 4445 14433 4479 14467
rect 6101 14433 6135 14467
rect 6929 14433 6963 14467
rect 7113 14433 7147 14467
rect 12081 14433 12115 14467
rect 12357 14433 12391 14467
rect 1685 14365 1719 14399
rect 2237 14365 2271 14399
rect 2689 14365 2723 14399
rect 3433 14365 3467 14399
rect 4169 14365 4203 14399
rect 4905 14365 4939 14399
rect 6469 14365 6503 14399
rect 9045 14365 9079 14399
rect 12624 14365 12658 14399
rect 15218 14365 15252 14399
rect 15485 14365 15519 14399
rect 16966 14365 17000 14399
rect 17233 14365 17267 14399
rect 17509 14365 17543 14399
rect 17765 14365 17799 14399
rect 20821 14365 20855 14399
rect 21097 14365 21131 14399
rect 9312 14297 9346 14331
rect 11836 14297 11870 14331
rect 20554 14297 20588 14331
rect 1501 14229 1535 14263
rect 2053 14229 2087 14263
rect 2513 14229 2547 14263
rect 3801 14229 3835 14263
rect 5273 14229 5307 14263
rect 5825 14229 5859 14263
rect 7205 14229 7239 14263
rect 7573 14229 7607 14263
rect 8309 14229 8343 14263
rect 13737 14229 13771 14263
rect 18889 14229 18923 14263
rect 21281 14229 21315 14263
rect 1961 14025 1995 14059
rect 2421 14025 2455 14059
rect 3985 14025 4019 14059
rect 4445 14025 4479 14059
rect 5089 14025 5123 14059
rect 5549 14025 5583 14059
rect 7113 14025 7147 14059
rect 9505 14025 9539 14059
rect 11161 14025 11195 14059
rect 14197 14025 14231 14059
rect 17417 14025 17451 14059
rect 17693 14025 17727 14059
rect 18797 14025 18831 14059
rect 19533 14025 19567 14059
rect 21189 14025 21223 14059
rect 7389 13957 7423 13991
rect 8392 13957 8426 13991
rect 10048 13957 10082 13991
rect 11621 13957 11655 13991
rect 12173 13957 12207 13991
rect 20646 13957 20680 13991
rect 1685 13889 1719 13923
rect 2145 13889 2179 13923
rect 2605 13889 2639 13923
rect 3065 13889 3099 13923
rect 4353 13889 4387 13923
rect 5457 13889 5491 13923
rect 13654 13889 13688 13923
rect 13921 13889 13955 13923
rect 15310 13889 15344 13923
rect 17049 13889 17083 13923
rect 20913 13889 20947 13923
rect 21373 13889 21407 13923
rect 4537 13821 4571 13855
rect 5641 13821 5675 13855
rect 6377 13821 6411 13855
rect 7849 13821 7883 13855
rect 8125 13821 8159 13855
rect 9781 13821 9815 13855
rect 15577 13821 15611 13855
rect 15853 13821 15887 13855
rect 16221 13821 16255 13855
rect 18061 13821 18095 13855
rect 2881 13753 2915 13787
rect 12541 13753 12575 13787
rect 18429 13753 18463 13787
rect 19165 13753 19199 13787
rect 1501 13685 1535 13719
rect 3433 13685 3467 13719
rect 3157 13481 3191 13515
rect 4813 13481 4847 13515
rect 10333 13481 10367 13515
rect 14105 13481 14139 13515
rect 15117 13481 15151 13515
rect 15853 13481 15887 13515
rect 18889 13481 18923 13515
rect 19349 13481 19383 13515
rect 2237 13413 2271 13447
rect 7205 13413 7239 13447
rect 14473 13413 14507 13447
rect 20361 13413 20395 13447
rect 5457 13345 5491 13379
rect 6469 13345 6503 13379
rect 6929 13345 6963 13379
rect 7849 13345 7883 13379
rect 8953 13345 8987 13379
rect 20913 13345 20947 13379
rect 1685 13277 1719 13311
rect 2697 13277 2731 13311
rect 3341 13277 3375 13311
rect 5181 13277 5215 13311
rect 6285 13277 6319 13311
rect 7573 13277 7607 13311
rect 10609 13277 10643 13311
rect 10977 13277 11011 13311
rect 17233 13277 17267 13311
rect 17509 13277 17543 13311
rect 20085 13277 20119 13311
rect 2053 13209 2087 13243
rect 4353 13209 4387 13243
rect 6193 13209 6227 13243
rect 8217 13209 8251 13243
rect 9220 13209 9254 13243
rect 12817 13209 12851 13243
rect 13737 13209 13771 13243
rect 16966 13209 17000 13243
rect 17776 13209 17810 13243
rect 1501 13141 1535 13175
rect 2881 13141 2915 13175
rect 3985 13141 4019 13175
rect 5273 13141 5307 13175
rect 5825 13141 5859 13175
rect 7665 13141 7699 13175
rect 11345 13141 11379 13175
rect 11805 13141 11839 13175
rect 12173 13141 12207 13175
rect 12541 13141 12575 13175
rect 13277 13141 13311 13175
rect 15577 13141 15611 13175
rect 19901 13141 19935 13175
rect 20729 13141 20763 13175
rect 20821 13141 20855 13175
rect 2329 12937 2363 12971
rect 2881 12937 2915 12971
rect 3617 12937 3651 12971
rect 4537 12937 4571 12971
rect 5273 12937 5307 12971
rect 5733 12937 5767 12971
rect 10793 12937 10827 12971
rect 13093 12937 13127 12971
rect 14933 12937 14967 12971
rect 19165 12937 19199 12971
rect 19441 12937 19475 12971
rect 20269 12937 20303 12971
rect 7481 12869 7515 12903
rect 10250 12869 10284 12903
rect 13369 12869 13403 12903
rect 13829 12869 13863 12903
rect 18052 12869 18086 12903
rect 1961 12801 1995 12835
rect 2973 12801 3007 12835
rect 3801 12801 3835 12835
rect 4077 12801 4111 12835
rect 4997 12801 5031 12835
rect 5641 12801 5675 12835
rect 7573 12801 7607 12835
rect 8125 12801 8159 12835
rect 10517 12801 10551 12835
rect 11713 12801 11747 12835
rect 11969 12801 12003 12835
rect 16046 12801 16080 12835
rect 20085 12801 20119 12835
rect 20821 12801 20855 12835
rect 1685 12733 1719 12767
rect 1869 12733 1903 12767
rect 2789 12733 2823 12767
rect 5825 12733 5859 12767
rect 7757 12733 7791 12767
rect 14657 12733 14691 12767
rect 16313 12733 16347 12767
rect 17785 12733 17819 12767
rect 20545 12733 20579 12767
rect 8585 12665 8619 12699
rect 14197 12665 14231 12699
rect 3341 12597 3375 12631
rect 4261 12597 4295 12631
rect 6653 12597 6687 12631
rect 7113 12597 7147 12631
rect 9137 12597 9171 12631
rect 16773 12597 16807 12631
rect 17325 12597 17359 12631
rect 8033 12393 8067 12427
rect 11161 12393 11195 12427
rect 13737 12393 13771 12427
rect 16589 12393 16623 12427
rect 18797 12393 18831 12427
rect 19717 12393 19751 12427
rect 20821 12393 20855 12427
rect 21189 12393 21223 12427
rect 7665 12325 7699 12359
rect 8401 12325 8435 12359
rect 10517 12325 10551 12359
rect 16221 12325 16255 12359
rect 19441 12325 19475 12359
rect 1961 12257 1995 12291
rect 2605 12257 2639 12291
rect 2789 12257 2823 12291
rect 4353 12257 4387 12291
rect 5273 12257 5307 12291
rect 6837 12257 6871 12291
rect 6929 12257 6963 12291
rect 13001 12257 13035 12291
rect 14197 12257 14231 12291
rect 14565 12257 14599 12291
rect 14841 12257 14875 12291
rect 20361 12257 20395 12291
rect 2237 12189 2271 12223
rect 4169 12189 4203 12223
rect 9137 12189 9171 12223
rect 15108 12189 15142 12223
rect 17417 12189 17451 12223
rect 19257 12189 19291 12223
rect 21281 12189 21315 12223
rect 2881 12121 2915 12155
rect 5457 12121 5491 12155
rect 6101 12121 6135 12155
rect 7021 12121 7055 12155
rect 9404 12121 9438 12155
rect 10793 12121 10827 12155
rect 12633 12121 12667 12155
rect 17662 12121 17696 12155
rect 20085 12121 20119 12155
rect 3249 12053 3283 12087
rect 3801 12053 3835 12087
rect 4261 12053 4295 12087
rect 5365 12053 5399 12087
rect 5825 12053 5859 12087
rect 7389 12053 7423 12087
rect 11529 12053 11563 12087
rect 11989 12053 12023 12087
rect 13369 12053 13403 12087
rect 17049 12053 17083 12087
rect 20177 12053 20211 12087
rect 2513 11849 2547 11883
rect 2973 11849 3007 11883
rect 3801 11849 3835 11883
rect 4261 11849 4295 11883
rect 6929 11849 6963 11883
rect 9505 11849 9539 11883
rect 12081 11849 12115 11883
rect 12541 11849 12575 11883
rect 18061 11849 18095 11883
rect 19165 11849 19199 11883
rect 19809 11849 19843 11883
rect 20177 11849 20211 11883
rect 20453 11849 20487 11883
rect 2881 11781 2915 11815
rect 4997 11781 5031 11815
rect 10618 11781 10652 11815
rect 11621 11781 11655 11815
rect 14390 11781 14424 11815
rect 15200 11781 15234 11815
rect 19717 11781 19751 11815
rect 4169 11713 4203 11747
rect 7297 11713 7331 11747
rect 16681 11713 16715 11747
rect 16937 11713 16971 11747
rect 18981 11713 19015 11747
rect 20821 11713 20855 11747
rect 1961 11645 1995 11679
rect 2237 11645 2271 11679
rect 3065 11645 3099 11679
rect 4445 11645 4479 11679
rect 5365 11645 5399 11679
rect 5733 11645 5767 11679
rect 7389 11645 7423 11679
rect 7573 11645 7607 11679
rect 10878 11645 10912 11679
rect 12909 11645 12943 11679
rect 14657 11645 14691 11679
rect 14933 11645 14967 11679
rect 19625 11645 19659 11679
rect 20913 11645 20947 11679
rect 21005 11645 21039 11679
rect 7941 11577 7975 11611
rect 8769 11577 8803 11611
rect 13277 11577 13311 11611
rect 6469 11509 6503 11543
rect 8309 11509 8343 11543
rect 9137 11509 9171 11543
rect 16313 11509 16347 11543
rect 18429 11509 18463 11543
rect 1593 11305 1627 11339
rect 3341 11305 3375 11339
rect 3985 11305 4019 11339
rect 4537 11305 4571 11339
rect 10885 11305 10919 11339
rect 11253 11305 11287 11339
rect 17601 11305 17635 11339
rect 19349 11305 19383 11339
rect 21189 11305 21223 11339
rect 7113 11237 7147 11271
rect 10517 11237 10551 11271
rect 13093 11237 13127 11271
rect 16129 11237 16163 11271
rect 17969 11237 18003 11271
rect 18337 11237 18371 11271
rect 18889 11237 18923 11271
rect 2237 11169 2271 11203
rect 2789 11169 2823 11203
rect 5181 11169 5215 11203
rect 6193 11169 6227 11203
rect 7665 11169 7699 11203
rect 9137 11169 9171 11203
rect 11713 11169 11747 11203
rect 14473 11169 14507 11203
rect 20729 11169 20763 11203
rect 6101 11101 6135 11135
rect 7573 11101 7607 11135
rect 9393 11101 9427 11135
rect 13369 11101 13403 11135
rect 16957 11101 16991 11135
rect 18705 11101 18739 11135
rect 2053 11033 2087 11067
rect 2881 11033 2915 11067
rect 3893 11033 3927 11067
rect 4905 11033 4939 11067
rect 4997 11033 5031 11067
rect 6009 11033 6043 11067
rect 6653 11033 6687 11067
rect 8125 11033 8159 11067
rect 11958 11033 11992 11067
rect 15301 11033 15335 11067
rect 20484 11033 20518 11067
rect 21281 11033 21315 11067
rect 1961 10965 1995 10999
rect 2973 10965 3007 10999
rect 5641 10965 5675 10999
rect 7481 10965 7515 10999
rect 8493 10965 8527 10999
rect 14841 10965 14875 10999
rect 15761 10965 15795 10999
rect 16497 10965 16531 10999
rect 17233 10965 17267 10999
rect 2881 10761 2915 10795
rect 4629 10761 4663 10795
rect 7757 10761 7791 10795
rect 10885 10761 10919 10795
rect 11989 10761 12023 10795
rect 17417 10761 17451 10795
rect 20545 10761 20579 10795
rect 3525 10693 3559 10727
rect 6377 10693 6411 10727
rect 7389 10693 7423 10727
rect 8125 10693 8159 10727
rect 10272 10693 10306 10727
rect 14298 10693 14332 10727
rect 18530 10693 18564 10727
rect 19432 10693 19466 10727
rect 21097 10693 21131 10727
rect 1961 10625 1995 10659
rect 5825 10625 5859 10659
rect 8769 10625 8803 10659
rect 10517 10625 10551 10659
rect 12817 10625 12851 10659
rect 18797 10625 18831 10659
rect 19165 10625 19199 10659
rect 21281 10625 21315 10659
rect 2237 10557 2271 10591
rect 2973 10557 3007 10591
rect 3065 10557 3099 10591
rect 4445 10557 4479 10591
rect 4537 10557 4571 10591
rect 5457 10557 5491 10591
rect 11621 10557 11655 10591
rect 14565 10557 14599 10591
rect 17049 10557 17083 10591
rect 13185 10489 13219 10523
rect 2513 10421 2547 10455
rect 4997 10421 5031 10455
rect 7021 10421 7055 10455
rect 9137 10421 9171 10455
rect 12449 10421 12483 10455
rect 14933 10421 14967 10455
rect 15485 10421 15519 10455
rect 15853 10421 15887 10455
rect 16221 10421 16255 10455
rect 16681 10421 16715 10455
rect 1685 10217 1719 10251
rect 3433 10217 3467 10251
rect 4905 10217 4939 10251
rect 6285 10217 6319 10251
rect 8953 10217 8987 10251
rect 10701 10217 10735 10251
rect 11529 10217 11563 10251
rect 14841 10217 14875 10251
rect 16865 10217 16899 10251
rect 2973 10149 3007 10183
rect 8585 10149 8619 10183
rect 11989 10149 12023 10183
rect 16589 10149 16623 10183
rect 2145 10081 2179 10115
rect 2329 10081 2363 10115
rect 4353 10081 4387 10115
rect 5733 10081 5767 10115
rect 5917 10081 5951 10115
rect 6837 10081 6871 10115
rect 8033 10081 8067 10115
rect 8125 10081 8159 10115
rect 10333 10081 10367 10115
rect 18245 10081 18279 10115
rect 19993 10081 20027 10115
rect 20545 10081 20579 10115
rect 20821 10081 20855 10115
rect 2053 10013 2087 10047
rect 3249 10013 3283 10047
rect 4445 10013 4479 10047
rect 5641 10013 5675 10047
rect 11805 10013 11839 10047
rect 13645 10013 13679 10047
rect 15209 10013 15243 10047
rect 19717 10013 19751 10047
rect 2789 9945 2823 9979
rect 6653 9945 6687 9979
rect 7481 9945 7515 9979
rect 8217 9945 8251 9979
rect 10066 9945 10100 9979
rect 11161 9945 11195 9979
rect 13378 9945 13412 9979
rect 14565 9945 14599 9979
rect 15476 9945 15510 9979
rect 17978 9945 18012 9979
rect 20177 9945 20211 9979
rect 3893 9877 3927 9911
rect 4537 9877 4571 9911
rect 5273 9877 5307 9911
rect 6745 9877 6779 9911
rect 12265 9877 12299 9911
rect 14105 9877 14139 9911
rect 18797 9877 18831 9911
rect 19533 9877 19567 9911
rect 10885 9673 10919 9707
rect 1501 9605 1535 9639
rect 3249 9605 3283 9639
rect 16681 9605 16715 9639
rect 2145 9537 2179 9571
rect 3157 9537 3191 9571
rect 3893 9537 3927 9571
rect 4537 9537 4571 9571
rect 5181 9537 5215 9571
rect 7021 9537 7055 9571
rect 7757 9537 7791 9571
rect 8401 9537 8435 9571
rect 9485 9537 9519 9571
rect 12918 9537 12952 9571
rect 14177 9537 14211 9571
rect 16313 9537 16347 9571
rect 17417 9537 17451 9571
rect 19450 9537 19484 9571
rect 20269 9537 20303 9571
rect 20545 9537 20579 9571
rect 1961 9469 1995 9503
rect 2053 9469 2087 9503
rect 3341 9469 3375 9503
rect 4905 9469 4939 9503
rect 5089 9469 5123 9503
rect 6745 9469 6779 9503
rect 7849 9469 7883 9503
rect 8033 9469 8067 9503
rect 9229 9469 9263 9503
rect 13185 9469 13219 9503
rect 13921 9469 13955 9503
rect 17509 9469 17543 9503
rect 17601 9469 17635 9503
rect 19717 9469 19751 9503
rect 20821 9469 20855 9503
rect 4353 9401 4387 9435
rect 13553 9401 13587 9435
rect 17049 9401 17083 9435
rect 18337 9401 18371 9435
rect 20085 9401 20119 9435
rect 2513 9333 2547 9367
rect 2789 9333 2823 9367
rect 3985 9333 4019 9367
rect 5549 9333 5583 9367
rect 5917 9333 5951 9367
rect 7389 9333 7423 9367
rect 8861 9333 8895 9367
rect 10609 9333 10643 9367
rect 11805 9333 11839 9367
rect 15301 9333 15335 9367
rect 15577 9333 15611 9367
rect 7941 9129 7975 9163
rect 8585 9129 8619 9163
rect 9321 9129 9355 9163
rect 10977 9129 11011 9163
rect 19809 9129 19843 9163
rect 6285 9061 6319 9095
rect 7665 9061 7699 9095
rect 11529 9061 11563 9095
rect 14197 9061 14231 9095
rect 19349 9061 19383 9095
rect 1961 8993 1995 9027
rect 3157 8993 3191 9027
rect 3985 8993 4019 9027
rect 5457 8993 5491 9027
rect 7113 8993 7147 9027
rect 10701 8993 10735 9027
rect 11897 8993 11931 9027
rect 15577 8993 15611 9027
rect 18061 8993 18095 9027
rect 20361 8993 20395 9027
rect 2237 8925 2271 8959
rect 5273 8925 5307 8959
rect 7297 8925 7331 8959
rect 12153 8925 12187 8959
rect 13553 8925 13587 8959
rect 17509 8925 17543 8959
rect 18337 8925 18371 8959
rect 19533 8925 19567 8959
rect 21281 8925 21315 8959
rect 2513 8857 2547 8891
rect 2697 8857 2731 8891
rect 4169 8857 4203 8891
rect 5365 8857 5399 8891
rect 10456 8857 10490 8891
rect 15310 8857 15344 8891
rect 17242 8857 17276 8891
rect 17877 8857 17911 8891
rect 21097 8857 21131 8891
rect 4077 8789 4111 8823
rect 4537 8789 4571 8823
rect 4905 8789 4939 8823
rect 5917 8789 5951 8823
rect 7205 8789 7239 8823
rect 9045 8789 9079 8823
rect 13277 8789 13311 8823
rect 16129 8789 16163 8823
rect 18705 8789 18739 8823
rect 20177 8789 20211 8823
rect 20269 8789 20303 8823
rect 3525 8585 3559 8619
rect 5825 8585 5859 8619
rect 6469 8585 6503 8619
rect 8769 8585 8803 8619
rect 9137 8585 9171 8619
rect 10793 8585 10827 8619
rect 11713 8585 11747 8619
rect 16681 8585 16715 8619
rect 20085 8585 20119 8619
rect 20453 8585 20487 8619
rect 2973 8517 3007 8551
rect 7573 8517 7607 8551
rect 8217 8517 8251 8551
rect 16037 8517 16071 8551
rect 17794 8517 17828 8551
rect 18337 8517 18371 8551
rect 18705 8517 18739 8551
rect 20545 8517 20579 8551
rect 21281 8517 21315 8551
rect 1961 8449 1995 8483
rect 2881 8449 2915 8483
rect 5089 8449 5123 8483
rect 5457 8449 5491 8483
rect 7481 8449 7515 8483
rect 9413 8449 9447 8483
rect 9669 8449 9703 8483
rect 13113 8449 13147 8483
rect 14657 8449 14691 8483
rect 15025 8449 15059 8483
rect 19441 8449 19475 8483
rect 2237 8381 2271 8415
rect 3157 8381 3191 8415
rect 4077 8381 4111 8415
rect 4445 8381 4479 8415
rect 7757 8381 7791 8415
rect 13369 8381 13403 8415
rect 18061 8381 18095 8415
rect 19257 8381 19291 8415
rect 19349 8381 19383 8415
rect 20637 8381 20671 8415
rect 2513 8313 2547 8347
rect 7113 8313 7147 8347
rect 11989 8313 12023 8347
rect 15393 8313 15427 8347
rect 21097 8313 21131 8347
rect 6837 8245 6871 8279
rect 11161 8245 11195 8279
rect 13737 8245 13771 8279
rect 14105 8245 14139 8279
rect 15761 8245 15795 8279
rect 19809 8245 19843 8279
rect 3801 8041 3835 8075
rect 4261 8041 4295 8075
rect 5917 8041 5951 8075
rect 8953 8041 8987 8075
rect 9413 8041 9447 8075
rect 12173 8041 12207 8075
rect 18889 8041 18923 8075
rect 21189 8041 21223 8075
rect 2881 7973 2915 8007
rect 3341 7973 3375 8007
rect 8585 7973 8619 8007
rect 13185 7973 13219 8007
rect 2053 7905 2087 7939
rect 2237 7905 2271 7939
rect 4997 7905 5031 7939
rect 5181 7905 5215 7939
rect 6929 7905 6963 7939
rect 7113 7905 7147 7939
rect 7573 7905 7607 7939
rect 7757 7905 7791 7939
rect 12541 7905 12575 7939
rect 12725 7905 12759 7939
rect 2697 7837 2731 7871
rect 3157 7837 3191 7871
rect 3985 7837 4019 7871
rect 5273 7837 5307 7871
rect 7849 7837 7883 7871
rect 10793 7837 10827 7871
rect 12817 7837 12851 7871
rect 14657 7837 14691 7871
rect 16865 7837 16899 7871
rect 17132 7837 17166 7871
rect 18705 7837 18739 7871
rect 20729 7837 20763 7871
rect 10526 7769 10560 7803
rect 14381 7769 14415 7803
rect 16129 7769 16163 7803
rect 16497 7769 16531 7803
rect 20484 7769 20518 7803
rect 21281 7769 21315 7803
rect 1593 7701 1627 7735
rect 1961 7701 1995 7735
rect 5641 7701 5675 7735
rect 6469 7701 6503 7735
rect 6837 7701 6871 7735
rect 8217 7701 8251 7735
rect 11161 7701 11195 7735
rect 11805 7701 11839 7735
rect 13737 7701 13771 7735
rect 15025 7701 15059 7735
rect 15761 7701 15795 7735
rect 18245 7701 18279 7735
rect 19349 7701 19383 7735
rect 1869 7497 1903 7531
rect 2329 7497 2363 7531
rect 3985 7497 4019 7531
rect 4353 7497 4387 7531
rect 4997 7497 5031 7531
rect 5089 7497 5123 7531
rect 6745 7497 6779 7531
rect 9321 7497 9355 7531
rect 14381 7497 14415 7531
rect 17509 7497 17543 7531
rect 20637 7497 20671 7531
rect 21097 7497 21131 7531
rect 2881 7429 2915 7463
rect 8677 7429 8711 7463
rect 14902 7429 14936 7463
rect 20094 7429 20128 7463
rect 21005 7429 21039 7463
rect 1961 7361 1995 7395
rect 2697 7361 2731 7395
rect 3341 7361 3375 7395
rect 6837 7361 6871 7395
rect 7389 7361 7423 7395
rect 10445 7361 10479 7395
rect 12817 7361 12851 7395
rect 13645 7361 13679 7395
rect 14657 7361 14691 7395
rect 16773 7361 16807 7395
rect 17325 7361 17359 7395
rect 18153 7361 18187 7395
rect 18245 7361 18279 7395
rect 1685 7293 1719 7327
rect 3709 7293 3743 7327
rect 3893 7293 3927 7327
rect 5273 7293 5307 7327
rect 6929 7293 6963 7327
rect 8309 7293 8343 7327
rect 10701 7293 10735 7327
rect 12357 7293 12391 7327
rect 18429 7293 18463 7327
rect 20361 7293 20395 7327
rect 21281 7293 21315 7327
rect 4629 7225 4663 7259
rect 6009 7225 6043 7259
rect 7573 7225 7607 7259
rect 11069 7225 11103 7259
rect 12633 7225 12667 7259
rect 17785 7225 17819 7259
rect 3157 7157 3191 7191
rect 6377 7157 6411 7191
rect 7941 7157 7975 7191
rect 9045 7157 9079 7191
rect 11529 7157 11563 7191
rect 11989 7157 12023 7191
rect 13185 7157 13219 7191
rect 14013 7157 14047 7191
rect 16037 7157 16071 7191
rect 18981 7157 19015 7191
rect 1685 6953 1719 6987
rect 7389 6953 7423 6987
rect 9137 6953 9171 6987
rect 15393 6953 15427 6987
rect 2329 6817 2363 6851
rect 3341 6817 3375 6851
rect 4445 6817 4479 6851
rect 5641 6817 5675 6851
rect 6837 6817 6871 6851
rect 6929 6817 6963 6851
rect 8033 6817 8067 6851
rect 10517 6817 10551 6851
rect 12449 6817 12483 6851
rect 14381 6817 14415 6851
rect 15945 6817 15979 6851
rect 16129 6817 16163 6851
rect 17417 6817 17451 6851
rect 18337 6817 18371 6851
rect 21097 6817 21131 6851
rect 3065 6749 3099 6783
rect 5457 6749 5491 6783
rect 10261 6749 10295 6783
rect 14657 6749 14691 6783
rect 17049 6749 17083 6783
rect 17693 6749 17727 6783
rect 18889 6749 18923 6783
rect 20370 6749 20404 6783
rect 20637 6749 20671 6783
rect 2053 6681 2087 6715
rect 6745 6681 6779 6715
rect 8585 6681 8619 6715
rect 12182 6681 12216 6715
rect 21281 6681 21315 6715
rect 2145 6613 2179 6647
rect 2697 6613 2731 6647
rect 3157 6613 3191 6647
rect 3801 6613 3835 6647
rect 4169 6613 4203 6647
rect 4261 6613 4295 6647
rect 5089 6613 5123 6647
rect 5549 6613 5583 6647
rect 6377 6613 6411 6647
rect 7757 6613 7791 6647
rect 7849 6613 7883 6647
rect 11069 6613 11103 6647
rect 12817 6613 12851 6647
rect 13093 6613 13127 6647
rect 13645 6613 13679 6647
rect 14565 6613 14599 6647
rect 15025 6613 15059 6647
rect 16221 6613 16255 6647
rect 16589 6613 16623 6647
rect 16865 6613 16899 6647
rect 17601 6613 17635 6647
rect 18061 6613 18095 6647
rect 18705 6613 18739 6647
rect 19257 6613 19291 6647
rect 2697 6409 2731 6443
rect 3065 6409 3099 6443
rect 3985 6409 4019 6443
rect 4353 6409 4387 6443
rect 6561 6409 6595 6443
rect 7113 6409 7147 6443
rect 8953 6409 8987 6443
rect 12633 6409 12667 6443
rect 13001 6409 13035 6443
rect 16773 6409 16807 6443
rect 19809 6409 19843 6443
rect 1501 6341 1535 6375
rect 2605 6341 2639 6375
rect 8125 6341 8159 6375
rect 14114 6341 14148 6375
rect 4445 6273 4479 6307
rect 4997 6273 5031 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 7481 6273 7515 6307
rect 10353 6273 10387 6307
rect 10609 6273 10643 6307
rect 10977 6273 11011 6307
rect 11621 6273 11655 6307
rect 14381 6273 14415 6307
rect 16046 6273 16080 6307
rect 16313 6273 16347 6307
rect 17886 6273 17920 6307
rect 18153 6273 18187 6307
rect 18521 6273 18555 6307
rect 19165 6273 19199 6307
rect 19901 6273 19935 6307
rect 20821 6273 20855 6307
rect 2513 6205 2547 6239
rect 3341 6205 3375 6239
rect 4629 6205 4663 6239
rect 5549 6205 5583 6239
rect 7573 6205 7607 6239
rect 7665 6205 7699 6239
rect 19625 6205 19659 6239
rect 20545 6205 20579 6239
rect 5181 6137 5215 6171
rect 6009 6137 6043 6171
rect 1593 6069 1627 6103
rect 2053 6069 2087 6103
rect 8585 6069 8619 6103
rect 9229 6069 9263 6103
rect 12265 6069 12299 6103
rect 14933 6069 14967 6103
rect 18705 6069 18739 6103
rect 19073 6069 19107 6103
rect 20269 6069 20303 6103
rect 2421 5865 2455 5899
rect 3433 5865 3467 5899
rect 12357 5865 12391 5899
rect 14197 5865 14231 5899
rect 16313 5865 16347 5899
rect 20545 5865 20579 5899
rect 5733 5797 5767 5831
rect 6193 5797 6227 5831
rect 7113 5797 7147 5831
rect 20269 5797 20303 5831
rect 1869 5729 1903 5763
rect 1961 5729 1995 5763
rect 2789 5729 2823 5763
rect 2973 5729 3007 5763
rect 4813 5729 4847 5763
rect 10425 5729 10459 5763
rect 10977 5729 11011 5763
rect 12817 5729 12851 5763
rect 13277 5729 13311 5763
rect 14473 5729 14507 5763
rect 17049 5729 17083 5763
rect 19717 5729 19751 5763
rect 21189 5729 21223 5763
rect 2053 5661 2087 5695
rect 3065 5661 3099 5695
rect 3801 5661 3835 5695
rect 4445 5661 4479 5695
rect 5917 5661 5951 5695
rect 6377 5661 6411 5695
rect 6837 5661 6871 5695
rect 7297 5661 7331 5695
rect 7941 5661 7975 5695
rect 8309 5661 8343 5695
rect 14740 5661 14774 5695
rect 16129 5661 16163 5695
rect 16589 5661 16623 5695
rect 17305 5661 17339 5695
rect 18889 5661 18923 5695
rect 19901 5661 19935 5695
rect 21005 5661 21039 5695
rect 5089 5593 5123 5627
rect 10180 5593 10214 5627
rect 11244 5593 11278 5627
rect 20913 5593 20947 5627
rect 3985 5525 4019 5559
rect 4261 5525 4295 5559
rect 4997 5525 5031 5559
rect 5457 5525 5491 5559
rect 6653 5525 6687 5559
rect 9045 5525 9079 5559
rect 13737 5525 13771 5559
rect 15853 5525 15887 5559
rect 16773 5525 16807 5559
rect 18429 5525 18463 5559
rect 18705 5525 18739 5559
rect 19809 5525 19843 5559
rect 2513 5321 2547 5355
rect 3157 5321 3191 5355
rect 4261 5321 4295 5355
rect 5641 5321 5675 5355
rect 6469 5321 6503 5355
rect 6837 5321 6871 5355
rect 7481 5321 7515 5355
rect 7849 5321 7883 5355
rect 9137 5321 9171 5355
rect 13921 5321 13955 5355
rect 15853 5321 15887 5355
rect 17601 5321 17635 5355
rect 19349 5321 19383 5355
rect 1501 5253 1535 5287
rect 1685 5253 1719 5287
rect 2605 5253 2639 5287
rect 21281 5253 21315 5287
rect 3341 5185 3375 5219
rect 4077 5185 4111 5219
rect 4537 5185 4571 5219
rect 5549 5185 5583 5219
rect 8493 5185 8527 5219
rect 10250 5185 10284 5219
rect 10517 5185 10551 5219
rect 10793 5185 10827 5219
rect 13286 5185 13320 5219
rect 13553 5185 13587 5219
rect 14289 5185 14323 5219
rect 14933 5185 14967 5219
rect 15209 5185 15243 5219
rect 15669 5185 15703 5219
rect 16129 5185 16163 5219
rect 17141 5185 17175 5219
rect 17233 5185 17267 5219
rect 17877 5185 17911 5219
rect 18429 5185 18463 5219
rect 19073 5185 19107 5219
rect 20462 5185 20496 5219
rect 20729 5185 20763 5219
rect 2697 5117 2731 5151
rect 3617 5117 3651 5151
rect 5825 5117 5859 5151
rect 6929 5117 6963 5151
rect 7113 5117 7147 5151
rect 7941 5117 7975 5151
rect 8125 5117 8159 5151
rect 11805 5117 11839 5151
rect 17049 5117 17083 5151
rect 12173 5049 12207 5083
rect 14473 5049 14507 5083
rect 18889 5049 18923 5083
rect 21097 5049 21131 5083
rect 2145 4981 2179 5015
rect 4721 4981 4755 5015
rect 5181 4981 5215 5015
rect 8677 4981 8711 5015
rect 14749 4981 14783 5015
rect 15393 4981 15427 5015
rect 16313 4981 16347 5015
rect 18061 4981 18095 5015
rect 18613 4981 18647 5015
rect 4905 4777 4939 4811
rect 5917 4777 5951 4811
rect 7941 4777 7975 4811
rect 10517 4777 10551 4811
rect 10793 4777 10827 4811
rect 11253 4777 11287 4811
rect 12909 4777 12943 4811
rect 20269 4777 20303 4811
rect 9689 4709 9723 4743
rect 16129 4709 16163 4743
rect 16589 4709 16623 4743
rect 19349 4709 19383 4743
rect 21281 4709 21315 4743
rect 1961 4641 1995 4675
rect 2605 4641 2639 4675
rect 4261 4641 4295 4675
rect 5273 4641 5307 4675
rect 5457 4641 5491 4675
rect 6561 4641 6595 4675
rect 9137 4641 9171 4675
rect 12633 4641 12667 4675
rect 14105 4641 14139 4675
rect 18889 4641 18923 4675
rect 20821 4641 20855 4675
rect 2237 4573 2271 4607
rect 4445 4573 4479 4607
rect 6285 4573 6319 4607
rect 7297 4573 7331 4607
rect 7757 4573 7791 4607
rect 8401 4573 8435 4607
rect 9321 4573 9355 4607
rect 9965 4573 9999 4607
rect 10977 4573 11011 4607
rect 13553 4573 13587 4607
rect 15945 4573 15979 4607
rect 16405 4573 16439 4607
rect 16957 4573 16991 4607
rect 18633 4573 18667 4607
rect 19625 4573 19659 4607
rect 20729 4573 20763 4607
rect 2789 4505 2823 4539
rect 3893 4505 3927 4539
rect 12366 4505 12400 4539
rect 14350 4505 14384 4539
rect 2881 4437 2915 4471
rect 3249 4437 3283 4471
rect 4537 4437 4571 4471
rect 5549 4437 5583 4471
rect 7481 4437 7515 4471
rect 8217 4437 8251 4471
rect 9229 4437 9263 4471
rect 10149 4437 10183 4471
rect 13737 4437 13771 4471
rect 15485 4437 15519 4471
rect 17141 4437 17175 4471
rect 17509 4437 17543 4471
rect 19809 4437 19843 4471
rect 20637 4437 20671 4471
rect 1777 4233 1811 4267
rect 1869 4233 1903 4267
rect 4629 4233 4663 4267
rect 6009 4233 6043 4267
rect 8125 4233 8159 4267
rect 10701 4233 10735 4267
rect 11713 4233 11747 4267
rect 16129 4233 16163 4267
rect 13614 4165 13648 4199
rect 20821 4165 20855 4199
rect 2881 4097 2915 4131
rect 3893 4097 3927 4131
rect 4445 4097 4479 4131
rect 4905 4097 4939 4131
rect 5365 4097 5399 4131
rect 5825 4097 5859 4131
rect 7021 4097 7055 4131
rect 7481 4097 7515 4131
rect 7941 4097 7975 4131
rect 8585 4097 8619 4131
rect 8861 4097 8895 4131
rect 9321 4097 9355 4131
rect 9588 4097 9622 4131
rect 12837 4097 12871 4131
rect 13093 4097 13127 4131
rect 13369 4097 13403 4131
rect 15025 4097 15059 4131
rect 15485 4097 15519 4131
rect 15945 4097 15979 4131
rect 17049 4097 17083 4131
rect 18061 4097 18095 4131
rect 19450 4097 19484 4131
rect 20177 4097 20211 4131
rect 20913 4097 20947 4131
rect 1685 4029 1719 4063
rect 2605 4029 2639 4063
rect 2789 4029 2823 4063
rect 6561 4029 6595 4063
rect 17141 4029 17175 4063
rect 17325 4029 17359 4063
rect 19717 4029 19751 4063
rect 21005 4029 21039 4063
rect 3249 3961 3283 3995
rect 3617 3961 3651 3995
rect 5549 3961 5583 3995
rect 7205 3961 7239 3995
rect 8401 3961 8435 3995
rect 14749 3961 14783 3995
rect 16681 3961 16715 3995
rect 20453 3961 20487 3995
rect 2237 3893 2271 3927
rect 4077 3893 4111 3927
rect 5089 3893 5123 3927
rect 7665 3893 7699 3927
rect 9045 3893 9079 3927
rect 11161 3893 11195 3927
rect 15209 3893 15243 3927
rect 15669 3893 15703 3927
rect 17877 3893 17911 3927
rect 18337 3893 18371 3927
rect 19993 3893 20027 3927
rect 2697 3689 2731 3723
rect 4905 3689 4939 3723
rect 6193 3689 6227 3723
rect 7205 3689 7239 3723
rect 12817 3689 12851 3723
rect 16129 3689 16163 3723
rect 16589 3689 16623 3723
rect 17509 3689 17543 3723
rect 20637 3689 20671 3723
rect 2421 3621 2455 3655
rect 9045 3621 9079 3655
rect 12081 3621 12115 3655
rect 13553 3621 13587 3655
rect 19993 3621 20027 3655
rect 1869 3553 1903 3587
rect 1961 3553 1995 3587
rect 3157 3553 3191 3587
rect 3341 3553 3375 3587
rect 4353 3553 4387 3587
rect 5457 3553 5491 3587
rect 6837 3553 6871 3587
rect 7665 3553 7699 3587
rect 7849 3553 7883 3587
rect 10425 3553 10459 3587
rect 10701 3553 10735 3587
rect 14749 3553 14783 3587
rect 18153 3553 18187 3587
rect 21189 3553 21223 3587
rect 4261 3485 4295 3519
rect 5273 3485 5307 3519
rect 6561 3485 6595 3519
rect 7573 3485 7607 3519
rect 8401 3485 8435 3519
rect 10158 3485 10192 3519
rect 12541 3485 12575 3519
rect 13001 3485 13035 3519
rect 13369 3485 13403 3519
rect 14289 3485 14323 3519
rect 16405 3485 16439 3519
rect 16865 3485 16899 3519
rect 17877 3485 17911 3519
rect 18797 3485 18831 3519
rect 19257 3485 19291 3519
rect 19809 3485 19843 3519
rect 21097 3485 21131 3519
rect 2053 3417 2087 3451
rect 3065 3417 3099 3451
rect 6653 3417 6687 3451
rect 10946 3417 10980 3451
rect 14994 3417 15028 3451
rect 21005 3417 21039 3451
rect 3801 3349 3835 3383
rect 4169 3349 4203 3383
rect 5365 3349 5399 3383
rect 8585 3349 8619 3383
rect 12357 3349 12391 3383
rect 14105 3349 14139 3383
rect 17049 3349 17083 3383
rect 17969 3349 18003 3383
rect 18613 3349 18647 3383
rect 19441 3349 19475 3383
rect 6009 3145 6043 3179
rect 7021 3145 7055 3179
rect 7665 3145 7699 3179
rect 8861 3145 8895 3179
rect 15853 3145 15887 3179
rect 17877 3145 17911 3179
rect 18245 3145 18279 3179
rect 18889 3145 18923 3179
rect 19349 3145 19383 3179
rect 7573 3077 7607 3111
rect 13553 3077 13587 3111
rect 1961 3009 1995 3043
rect 2237 3009 2271 3043
rect 2697 3009 2731 3043
rect 3157 3009 3191 3043
rect 3617 3009 3651 3043
rect 4077 3009 4111 3043
rect 5365 3009 5399 3043
rect 5825 3009 5859 3043
rect 6377 3009 6411 3043
rect 6837 3009 6871 3043
rect 8953 3009 8987 3043
rect 9873 3009 9907 3043
rect 10885 3009 10919 3043
rect 11069 3009 11103 3043
rect 11989 3009 12023 3043
rect 12081 3009 12115 3043
rect 12725 3009 12759 3043
rect 14197 3009 14231 3043
rect 14841 3009 14875 3043
rect 15945 3009 15979 3043
rect 16681 3009 16715 3043
rect 17233 3009 17267 3043
rect 18337 3009 18371 3043
rect 19257 3009 19291 3043
rect 19993 3009 20027 3043
rect 21373 3009 21407 3043
rect 5089 2941 5123 2975
rect 7481 2941 7515 2975
rect 9045 2941 9079 2975
rect 9597 2941 9631 2975
rect 9781 2941 9815 2975
rect 12173 2941 12207 2975
rect 13369 2941 13403 2975
rect 13461 2941 13495 2975
rect 15669 2941 15703 2975
rect 18429 2941 18463 2975
rect 19441 2941 19475 2975
rect 20269 2941 20303 2975
rect 2881 2873 2915 2907
rect 3801 2873 3835 2907
rect 6561 2873 6595 2907
rect 16865 2873 16899 2907
rect 3341 2805 3375 2839
rect 4261 2805 4295 2839
rect 8033 2805 8067 2839
rect 8493 2805 8527 2839
rect 10241 2805 10275 2839
rect 11621 2805 11655 2839
rect 12909 2805 12943 2839
rect 13921 2805 13955 2839
rect 14381 2805 14415 2839
rect 15025 2805 15059 2839
rect 16313 2805 16347 2839
rect 17417 2805 17451 2839
rect 21189 2805 21223 2839
rect 1869 2601 1903 2635
rect 2881 2601 2915 2635
rect 6837 2601 6871 2635
rect 12265 2601 12299 2635
rect 20637 2601 20671 2635
rect 2421 2533 2455 2567
rect 14841 2533 14875 2567
rect 15945 2533 15979 2567
rect 17969 2533 18003 2567
rect 19901 2533 19935 2567
rect 4629 2465 4663 2499
rect 5457 2465 5491 2499
rect 7665 2465 7699 2499
rect 9505 2465 9539 2499
rect 10609 2465 10643 2499
rect 11713 2465 11747 2499
rect 21189 2465 21223 2499
rect 1685 2397 1719 2431
rect 2789 2397 2823 2431
rect 3249 2397 3283 2431
rect 4353 2397 4387 2431
rect 5733 2397 5767 2431
rect 6653 2397 6687 2431
rect 7941 2397 7975 2431
rect 8585 2397 8619 2431
rect 9229 2397 9263 2431
rect 10333 2397 10367 2431
rect 11805 2397 11839 2431
rect 12633 2397 12667 2431
rect 13185 2397 13219 2431
rect 14105 2397 14139 2431
rect 14657 2397 14691 2431
rect 15209 2397 15243 2431
rect 15761 2397 15795 2431
rect 16681 2397 16715 2431
rect 17233 2397 17267 2431
rect 17785 2397 17819 2431
rect 18337 2397 18371 2431
rect 19257 2397 19291 2431
rect 20085 2397 20119 2431
rect 21005 2397 21039 2431
rect 2237 2329 2271 2363
rect 11897 2329 11931 2363
rect 21097 2329 21131 2363
rect 3433 2261 3467 2295
rect 8401 2261 8435 2295
rect 12817 2261 12851 2295
rect 13369 2261 13403 2295
rect 14289 2261 14323 2295
rect 15393 2261 15427 2295
rect 16865 2261 16899 2295
rect 17417 2261 17451 2295
rect 18521 2261 18555 2295
rect 19441 2261 19475 2295
<< metal1 >>
rect 16114 20748 16120 20800
rect 16172 20788 16178 20800
rect 17954 20788 17960 20800
rect 16172 20760 17960 20788
rect 16172 20748 16178 20760
rect 17954 20748 17960 20760
rect 18012 20748 18018 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 2038 20584 2044 20596
rect 1999 20556 2044 20584
rect 2038 20544 2044 20556
rect 2096 20544 2102 20596
rect 5718 20544 5724 20596
rect 5776 20584 5782 20596
rect 5905 20587 5963 20593
rect 5905 20584 5917 20587
rect 5776 20556 5917 20584
rect 5776 20544 5782 20556
rect 5905 20553 5917 20556
rect 5951 20553 5963 20587
rect 9861 20587 9919 20593
rect 9861 20584 9873 20587
rect 5905 20547 5963 20553
rect 6472 20556 9873 20584
rect 1670 20448 1676 20460
rect 1631 20420 1676 20448
rect 1670 20408 1676 20420
rect 1728 20408 1734 20460
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20448 2283 20451
rect 2590 20448 2596 20460
rect 2271 20420 2596 20448
rect 2271 20417 2283 20420
rect 2225 20411 2283 20417
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20417 2743 20451
rect 2958 20448 2964 20460
rect 2871 20420 2964 20448
rect 2685 20411 2743 20417
rect 2700 20380 2728 20411
rect 2958 20408 2964 20420
rect 3016 20448 3022 20460
rect 4893 20451 4951 20457
rect 4893 20448 4905 20451
rect 3016 20420 4905 20448
rect 3016 20408 3022 20420
rect 4893 20417 4905 20420
rect 4939 20417 4951 20451
rect 5920 20448 5948 20547
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 5920 20420 6377 20448
rect 4893 20411 4951 20417
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 4525 20383 4583 20389
rect 4525 20380 4537 20383
rect 2700 20352 4537 20380
rect 4525 20349 4537 20352
rect 4571 20380 4583 20383
rect 5166 20380 5172 20392
rect 4571 20352 5172 20380
rect 4571 20349 4583 20352
rect 4525 20343 4583 20349
rect 5166 20340 5172 20352
rect 5224 20340 5230 20392
rect 4706 20272 4712 20324
rect 4764 20312 4770 20324
rect 6472 20312 6500 20556
rect 9861 20553 9873 20556
rect 9907 20584 9919 20587
rect 11057 20587 11115 20593
rect 11057 20584 11069 20587
rect 9907 20556 11069 20584
rect 9907 20553 9919 20556
rect 9861 20547 9919 20553
rect 11057 20553 11069 20556
rect 11103 20553 11115 20587
rect 11057 20547 11115 20553
rect 16301 20587 16359 20593
rect 16301 20553 16313 20587
rect 16347 20553 16359 20587
rect 16301 20547 16359 20553
rect 11793 20519 11851 20525
rect 11793 20516 11805 20519
rect 6656 20488 11805 20516
rect 6656 20457 6684 20488
rect 11793 20485 11805 20488
rect 11839 20516 11851 20519
rect 12066 20516 12072 20528
rect 11839 20488 12072 20516
rect 11839 20485 11851 20488
rect 11793 20479 11851 20485
rect 12066 20476 12072 20488
rect 12124 20476 12130 20528
rect 16316 20516 16344 20547
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 17497 20587 17555 20593
rect 17497 20584 17509 20587
rect 17276 20556 17509 20584
rect 17276 20544 17282 20556
rect 17497 20553 17509 20556
rect 17543 20553 17555 20587
rect 21634 20584 21640 20596
rect 17497 20547 17555 20553
rect 19812 20556 21640 20584
rect 19812 20516 19840 20556
rect 21634 20544 21640 20556
rect 21692 20544 21698 20596
rect 16316 20488 19840 20516
rect 19886 20476 19892 20528
rect 19944 20516 19950 20528
rect 19944 20488 21128 20516
rect 19944 20476 19950 20488
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20417 6699 20451
rect 6641 20411 6699 20417
rect 7466 20408 7472 20460
rect 7524 20448 7530 20460
rect 7929 20451 7987 20457
rect 7929 20448 7941 20451
rect 7524 20420 7941 20448
rect 7524 20408 7530 20420
rect 7929 20417 7941 20420
rect 7975 20417 7987 20451
rect 7929 20411 7987 20417
rect 9309 20451 9367 20457
rect 9309 20417 9321 20451
rect 9355 20448 9367 20451
rect 9953 20451 10011 20457
rect 9953 20448 9965 20451
rect 9355 20420 9965 20448
rect 9355 20417 9367 20420
rect 9309 20411 9367 20417
rect 9953 20417 9965 20420
rect 9999 20417 10011 20451
rect 9953 20411 10011 20417
rect 12529 20451 12587 20457
rect 12529 20417 12541 20451
rect 12575 20448 12587 20451
rect 16114 20448 16120 20460
rect 12575 20420 15700 20448
rect 16075 20420 16120 20448
rect 12575 20417 12587 20420
rect 12529 20411 12587 20417
rect 7558 20340 7564 20392
rect 7616 20380 7622 20392
rect 7653 20383 7711 20389
rect 7653 20380 7665 20383
rect 7616 20352 7665 20380
rect 7616 20340 7622 20352
rect 7653 20349 7665 20352
rect 7699 20349 7711 20383
rect 7653 20343 7711 20349
rect 7837 20383 7895 20389
rect 7837 20349 7849 20383
rect 7883 20349 7895 20383
rect 9324 20380 9352 20411
rect 7837 20343 7895 20349
rect 7944 20352 9352 20380
rect 9769 20383 9827 20389
rect 4764 20284 6500 20312
rect 4764 20272 4770 20284
rect 7006 20272 7012 20324
rect 7064 20312 7070 20324
rect 7852 20312 7880 20343
rect 7064 20284 7880 20312
rect 7064 20272 7070 20284
rect 1486 20244 1492 20256
rect 1447 20216 1492 20244
rect 1486 20204 1492 20216
rect 1544 20204 1550 20256
rect 2222 20204 2228 20256
rect 2280 20244 2286 20256
rect 2501 20247 2559 20253
rect 2501 20244 2513 20247
rect 2280 20216 2513 20244
rect 2280 20204 2286 20216
rect 2501 20213 2513 20216
rect 2547 20213 2559 20247
rect 2501 20207 2559 20213
rect 3145 20247 3203 20253
rect 3145 20213 3157 20247
rect 3191 20244 3203 20247
rect 3418 20244 3424 20256
rect 3191 20216 3424 20244
rect 3191 20213 3203 20216
rect 3145 20207 3203 20213
rect 3418 20204 3424 20216
rect 3476 20204 3482 20256
rect 3878 20244 3884 20256
rect 3839 20216 3884 20244
rect 3878 20204 3884 20216
rect 3936 20204 3942 20256
rect 4154 20244 4160 20256
rect 4115 20216 4160 20244
rect 4154 20204 4160 20216
rect 4212 20204 4218 20256
rect 5258 20244 5264 20256
rect 5219 20216 5264 20244
rect 5258 20204 5264 20216
rect 5316 20204 5322 20256
rect 7650 20204 7656 20256
rect 7708 20244 7714 20256
rect 7944 20244 7972 20352
rect 9769 20349 9781 20383
rect 9815 20380 9827 20383
rect 13446 20380 13452 20392
rect 9815 20352 11284 20380
rect 13407 20352 13452 20380
rect 9815 20349 9827 20352
rect 9769 20343 9827 20349
rect 8294 20244 8300 20256
rect 7708 20216 7972 20244
rect 8255 20216 8300 20244
rect 7708 20204 7714 20216
rect 8294 20204 8300 20216
rect 8352 20204 8358 20256
rect 10318 20244 10324 20256
rect 10279 20216 10324 20244
rect 10318 20204 10324 20216
rect 10376 20204 10382 20256
rect 10778 20244 10784 20256
rect 10739 20216 10784 20244
rect 10778 20204 10784 20216
rect 10836 20204 10842 20256
rect 11256 20244 11284 20352
rect 13446 20340 13452 20352
rect 13504 20340 13510 20392
rect 15378 20340 15384 20392
rect 15436 20380 15442 20392
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 15436 20352 15485 20380
rect 15436 20340 15442 20352
rect 15473 20349 15485 20352
rect 15519 20349 15531 20383
rect 15672 20380 15700 20420
rect 16114 20408 16120 20420
rect 16172 20408 16178 20460
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20417 16727 20451
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 16669 20411 16727 20417
rect 16776 20420 17325 20448
rect 16298 20380 16304 20392
rect 15672 20352 16304 20380
rect 15473 20343 15531 20349
rect 16298 20340 16304 20352
rect 16356 20340 16362 20392
rect 12897 20315 12955 20321
rect 12897 20281 12909 20315
rect 12943 20312 12955 20315
rect 13814 20312 13820 20324
rect 12943 20284 13820 20312
rect 12943 20281 12955 20284
rect 12897 20275 12955 20281
rect 13814 20272 13820 20284
rect 13872 20272 13878 20324
rect 14642 20272 14648 20324
rect 14700 20312 14706 20324
rect 16684 20312 16712 20411
rect 14700 20284 16712 20312
rect 14700 20272 14706 20284
rect 12710 20244 12716 20256
rect 11256 20216 12716 20244
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 13538 20204 13544 20256
rect 13596 20244 13602 20256
rect 14369 20247 14427 20253
rect 14369 20244 14381 20247
rect 13596 20216 14381 20244
rect 13596 20204 13602 20216
rect 14369 20213 14381 20216
rect 14415 20244 14427 20247
rect 14829 20247 14887 20253
rect 14829 20244 14841 20247
rect 14415 20216 14841 20244
rect 14415 20213 14427 20216
rect 14369 20207 14427 20213
rect 14829 20213 14841 20216
rect 14875 20213 14887 20247
rect 14829 20207 14887 20213
rect 14918 20204 14924 20256
rect 14976 20244 14982 20256
rect 16776 20244 16804 20420
rect 17313 20417 17325 20420
rect 17359 20417 17371 20451
rect 19702 20448 19708 20460
rect 19663 20420 19708 20448
rect 17313 20411 17371 20417
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 19794 20408 19800 20460
rect 19852 20448 19858 20460
rect 21100 20457 21128 20488
rect 19981 20451 20039 20457
rect 19981 20448 19993 20451
rect 19852 20420 19993 20448
rect 19852 20408 19858 20420
rect 19981 20417 19993 20420
rect 20027 20417 20039 20451
rect 19981 20411 20039 20417
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20417 20591 20451
rect 20533 20411 20591 20417
rect 21085 20451 21143 20457
rect 21085 20417 21097 20451
rect 21131 20417 21143 20451
rect 21085 20411 21143 20417
rect 18230 20380 18236 20392
rect 18191 20352 18236 20380
rect 18230 20340 18236 20352
rect 18288 20340 18294 20392
rect 18874 20380 18880 20392
rect 18835 20352 18880 20380
rect 18874 20340 18880 20352
rect 18932 20340 18938 20392
rect 16853 20315 16911 20321
rect 16853 20281 16865 20315
rect 16899 20312 16911 20315
rect 20548 20312 20576 20411
rect 16899 20284 20576 20312
rect 16899 20281 16911 20284
rect 16853 20275 16911 20281
rect 14976 20216 16804 20244
rect 14976 20204 14982 20216
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 17865 20247 17923 20253
rect 17865 20244 17877 20247
rect 17276 20216 17877 20244
rect 17276 20204 17282 20216
rect 17865 20213 17877 20216
rect 17911 20213 17923 20247
rect 19518 20244 19524 20256
rect 19479 20216 19524 20244
rect 17865 20207 17923 20213
rect 19518 20204 19524 20216
rect 19576 20204 19582 20256
rect 20162 20244 20168 20256
rect 20123 20216 20168 20244
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 20714 20244 20720 20256
rect 20675 20216 20720 20244
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 21266 20244 21272 20256
rect 21227 20216 21272 20244
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 1670 20000 1676 20052
rect 1728 20040 1734 20052
rect 2501 20043 2559 20049
rect 2501 20040 2513 20043
rect 1728 20012 2513 20040
rect 1728 20000 1734 20012
rect 2501 20009 2513 20012
rect 2547 20009 2559 20043
rect 2501 20003 2559 20009
rect 2590 20000 2596 20052
rect 2648 20040 2654 20052
rect 2961 20043 3019 20049
rect 2961 20040 2973 20043
rect 2648 20012 2973 20040
rect 2648 20000 2654 20012
rect 2961 20009 2973 20012
rect 3007 20009 3019 20043
rect 2961 20003 3019 20009
rect 5997 20043 6055 20049
rect 5997 20009 6009 20043
rect 6043 20040 6055 20043
rect 10870 20040 10876 20052
rect 6043 20012 10876 20040
rect 6043 20009 6055 20012
rect 5997 20003 6055 20009
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 19702 20000 19708 20052
rect 19760 20040 19766 20052
rect 19981 20043 20039 20049
rect 19981 20040 19993 20043
rect 19760 20012 19993 20040
rect 19760 20000 19766 20012
rect 19981 20009 19993 20012
rect 20027 20009 20039 20043
rect 19981 20003 20039 20009
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20680 20012 20729 20040
rect 20680 20000 20686 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 1946 19932 1952 19984
rect 2004 19972 2010 19984
rect 2041 19975 2099 19981
rect 2041 19972 2053 19975
rect 2004 19944 2053 19972
rect 2004 19932 2010 19944
rect 2041 19941 2053 19944
rect 2087 19941 2099 19975
rect 13354 19972 13360 19984
rect 2041 19935 2099 19941
rect 10060 19944 13360 19972
rect 3973 19907 4031 19913
rect 3973 19873 3985 19907
rect 4019 19904 4031 19907
rect 4338 19904 4344 19916
rect 4019 19876 4344 19904
rect 4019 19873 4031 19876
rect 3973 19867 4031 19873
rect 4338 19864 4344 19876
rect 4396 19864 4402 19916
rect 10060 19913 10088 19944
rect 13354 19932 13360 19944
rect 13412 19932 13418 19984
rect 14737 19975 14795 19981
rect 14737 19941 14749 19975
rect 14783 19972 14795 19975
rect 19794 19972 19800 19984
rect 14783 19944 19800 19972
rect 14783 19941 14795 19944
rect 14737 19935 14795 19941
rect 19794 19932 19800 19944
rect 19852 19932 19858 19984
rect 8021 19907 8079 19913
rect 8021 19873 8033 19907
rect 8067 19904 8079 19907
rect 10045 19907 10103 19913
rect 8067 19876 8340 19904
rect 8067 19873 8079 19876
rect 8021 19867 8079 19873
rect 8312 19848 8340 19876
rect 10045 19873 10057 19907
rect 10091 19873 10103 19907
rect 10045 19867 10103 19873
rect 10137 19907 10195 19913
rect 10137 19873 10149 19907
rect 10183 19904 10195 19907
rect 10778 19904 10784 19916
rect 10183 19876 10784 19904
rect 10183 19873 10195 19876
rect 10137 19867 10195 19873
rect 10778 19864 10784 19876
rect 10836 19864 10842 19916
rect 11057 19907 11115 19913
rect 11057 19873 11069 19907
rect 11103 19904 11115 19907
rect 11698 19904 11704 19916
rect 11103 19876 11704 19904
rect 11103 19873 11115 19876
rect 11057 19867 11115 19873
rect 11698 19864 11704 19876
rect 11756 19864 11762 19916
rect 11882 19864 11888 19916
rect 11940 19904 11946 19916
rect 13081 19907 13139 19913
rect 13081 19904 13093 19907
rect 11940 19876 13093 19904
rect 11940 19864 11946 19876
rect 13081 19873 13093 19876
rect 13127 19873 13139 19907
rect 13081 19867 13139 19873
rect 13265 19907 13323 19913
rect 13265 19873 13277 19907
rect 13311 19904 13323 19907
rect 13814 19904 13820 19916
rect 13311 19876 13820 19904
rect 13311 19873 13323 19876
rect 13265 19867 13323 19873
rect 13814 19864 13820 19876
rect 13872 19904 13878 19916
rect 14642 19904 14648 19916
rect 13872 19876 14648 19904
rect 13872 19864 13878 19876
rect 14642 19864 14648 19876
rect 14700 19864 14706 19916
rect 15194 19904 15200 19916
rect 15155 19876 15200 19904
rect 15194 19864 15200 19876
rect 15252 19864 15258 19916
rect 16298 19864 16304 19916
rect 16356 19904 16362 19916
rect 16577 19907 16635 19913
rect 16577 19904 16589 19907
rect 16356 19876 16589 19904
rect 16356 19864 16362 19876
rect 16577 19873 16589 19876
rect 16623 19873 16635 19907
rect 17589 19907 17647 19913
rect 17589 19904 17601 19907
rect 16577 19867 16635 19873
rect 16684 19876 17601 19904
rect 1670 19836 1676 19848
rect 1631 19808 1676 19836
rect 1670 19796 1676 19808
rect 1728 19796 1734 19848
rect 2222 19836 2228 19848
rect 2183 19808 2228 19836
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 2682 19836 2688 19848
rect 2643 19808 2688 19836
rect 2682 19796 2688 19808
rect 2740 19796 2746 19848
rect 3145 19839 3203 19845
rect 3145 19805 3157 19839
rect 3191 19836 3203 19839
rect 3786 19836 3792 19848
rect 3191 19808 3792 19836
rect 3191 19805 3203 19808
rect 3145 19799 3203 19805
rect 3786 19796 3792 19808
rect 3844 19796 3850 19848
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19836 4123 19839
rect 4430 19836 4436 19848
rect 4111 19808 4436 19836
rect 4111 19805 4123 19808
rect 4065 19799 4123 19805
rect 4430 19796 4436 19808
rect 4488 19796 4494 19848
rect 6914 19796 6920 19848
rect 6972 19836 6978 19848
rect 8113 19839 8171 19845
rect 8113 19836 8125 19839
rect 6972 19808 8125 19836
rect 6972 19796 6978 19808
rect 8113 19805 8125 19808
rect 8159 19805 8171 19839
rect 8113 19799 8171 19805
rect 8294 19796 8300 19848
rect 8352 19796 8358 19848
rect 8478 19796 8484 19848
rect 8536 19836 8542 19848
rect 9493 19839 9551 19845
rect 9493 19836 9505 19839
rect 8536 19808 9505 19836
rect 8536 19796 8542 19808
rect 9493 19805 9505 19808
rect 9539 19836 9551 19839
rect 10229 19839 10287 19845
rect 10229 19836 10241 19839
rect 9539 19808 10241 19836
rect 9539 19805 9551 19808
rect 9493 19799 9551 19805
rect 10229 19805 10241 19808
rect 10275 19805 10287 19839
rect 12066 19836 12072 19848
rect 12027 19808 12072 19836
rect 10229 19799 10287 19805
rect 12066 19796 12072 19808
rect 12124 19836 12130 19848
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 12124 19808 12449 19836
rect 12124 19796 12130 19808
rect 12437 19805 12449 19808
rect 12483 19836 12495 19839
rect 12618 19836 12624 19848
rect 12483 19808 12624 19836
rect 12483 19805 12495 19808
rect 12437 19799 12495 19805
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 13538 19796 13544 19848
rect 13596 19836 13602 19848
rect 14553 19839 14611 19845
rect 14553 19836 14565 19839
rect 13596 19808 14565 19836
rect 13596 19796 13602 19808
rect 14553 19805 14565 19808
rect 14599 19805 14611 19839
rect 15378 19836 15384 19848
rect 15339 19808 15384 19836
rect 14553 19799 14611 19805
rect 4157 19771 4215 19777
rect 4157 19737 4169 19771
rect 4203 19768 4215 19771
rect 4801 19771 4859 19777
rect 4801 19768 4813 19771
rect 4203 19740 4813 19768
rect 4203 19737 4215 19740
rect 4157 19731 4215 19737
rect 4801 19737 4813 19740
rect 4847 19737 4859 19771
rect 4801 19731 4859 19737
rect 6825 19771 6883 19777
rect 6825 19737 6837 19771
rect 6871 19768 6883 19771
rect 7466 19768 7472 19780
rect 6871 19740 7472 19768
rect 6871 19737 6883 19740
rect 6825 19731 6883 19737
rect 7466 19728 7472 19740
rect 7524 19728 7530 19780
rect 8205 19771 8263 19777
rect 8205 19737 8217 19771
rect 8251 19768 8263 19771
rect 8941 19771 8999 19777
rect 8941 19768 8953 19771
rect 8251 19740 8953 19768
rect 8251 19737 8263 19740
rect 8205 19731 8263 19737
rect 8941 19737 8953 19740
rect 8987 19737 8999 19771
rect 8941 19731 8999 19737
rect 13357 19771 13415 19777
rect 13357 19737 13369 19771
rect 13403 19768 13415 19771
rect 14093 19771 14151 19777
rect 14093 19768 14105 19771
rect 13403 19740 14105 19768
rect 13403 19737 13415 19740
rect 13357 19731 13415 19737
rect 14093 19737 14105 19740
rect 14139 19737 14151 19771
rect 14568 19768 14596 19799
rect 15378 19796 15384 19808
rect 15436 19796 15442 19848
rect 16206 19796 16212 19848
rect 16264 19836 16270 19848
rect 16684 19836 16712 19876
rect 17589 19873 17601 19876
rect 17635 19873 17647 19907
rect 17589 19867 17647 19873
rect 19429 19907 19487 19913
rect 19429 19873 19441 19907
rect 19475 19904 19487 19907
rect 20438 19904 20444 19916
rect 19475 19876 20444 19904
rect 19475 19873 19487 19876
rect 19429 19867 19487 19873
rect 20438 19864 20444 19876
rect 20496 19864 20502 19916
rect 16264 19808 16712 19836
rect 16264 19796 16270 19808
rect 17494 19796 17500 19848
rect 17552 19836 17558 19848
rect 18693 19839 18751 19845
rect 18693 19836 18705 19839
rect 17552 19808 18705 19836
rect 17552 19796 17558 19808
rect 18693 19805 18705 19808
rect 18739 19805 18751 19839
rect 18693 19799 18751 19805
rect 18874 19796 18880 19848
rect 18932 19836 18938 19848
rect 19794 19836 19800 19848
rect 18932 19808 19800 19836
rect 18932 19796 18938 19808
rect 19794 19796 19800 19808
rect 19852 19796 19858 19848
rect 20530 19836 20536 19848
rect 20491 19808 20536 19836
rect 20530 19796 20536 19808
rect 20588 19796 20594 19848
rect 20806 19796 20812 19848
rect 20864 19836 20870 19848
rect 21085 19839 21143 19845
rect 21085 19836 21097 19839
rect 20864 19808 21097 19836
rect 20864 19796 20870 19808
rect 21085 19805 21097 19808
rect 21131 19805 21143 19839
rect 21085 19799 21143 19805
rect 15289 19771 15347 19777
rect 15289 19768 15301 19771
rect 14568 19740 15301 19768
rect 14093 19731 14151 19737
rect 15289 19737 15301 19740
rect 15335 19737 15347 19771
rect 15289 19731 15347 19737
rect 16485 19771 16543 19777
rect 16485 19737 16497 19771
rect 16531 19768 16543 19771
rect 17218 19768 17224 19780
rect 16531 19740 17224 19768
rect 16531 19737 16543 19740
rect 16485 19731 16543 19737
rect 17218 19728 17224 19740
rect 17276 19728 17282 19780
rect 17405 19771 17463 19777
rect 17405 19737 17417 19771
rect 17451 19768 17463 19771
rect 18049 19771 18107 19777
rect 18049 19768 18061 19771
rect 17451 19740 18061 19768
rect 17451 19737 17463 19740
rect 17405 19731 17463 19737
rect 18049 19737 18061 19740
rect 18095 19737 18107 19771
rect 18049 19731 18107 19737
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 4522 19700 4528 19712
rect 4483 19672 4528 19700
rect 4522 19660 4528 19672
rect 4580 19660 4586 19712
rect 5350 19660 5356 19712
rect 5408 19700 5414 19712
rect 5445 19703 5503 19709
rect 5445 19700 5457 19703
rect 5408 19672 5457 19700
rect 5408 19660 5414 19672
rect 5445 19669 5457 19672
rect 5491 19669 5503 19703
rect 5445 19663 5503 19669
rect 5994 19660 6000 19712
rect 6052 19700 6058 19712
rect 6273 19703 6331 19709
rect 6273 19700 6285 19703
rect 6052 19672 6285 19700
rect 6052 19660 6058 19672
rect 6273 19669 6285 19672
rect 6319 19669 6331 19703
rect 6273 19663 6331 19669
rect 7006 19660 7012 19712
rect 7064 19700 7070 19712
rect 7101 19703 7159 19709
rect 7101 19700 7113 19703
rect 7064 19672 7113 19700
rect 7064 19660 7070 19672
rect 7101 19669 7113 19672
rect 7147 19669 7159 19703
rect 7558 19700 7564 19712
rect 7519 19672 7564 19700
rect 7101 19663 7159 19669
rect 7558 19660 7564 19672
rect 7616 19660 7622 19712
rect 8573 19703 8631 19709
rect 8573 19669 8585 19703
rect 8619 19700 8631 19703
rect 9306 19700 9312 19712
rect 8619 19672 9312 19700
rect 8619 19669 8631 19672
rect 8573 19663 8631 19669
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 10597 19703 10655 19709
rect 10597 19669 10609 19703
rect 10643 19700 10655 19703
rect 11149 19703 11207 19709
rect 11149 19700 11161 19703
rect 10643 19672 11161 19700
rect 10643 19669 10655 19672
rect 10597 19663 10655 19669
rect 11149 19669 11161 19672
rect 11195 19669 11207 19703
rect 11149 19663 11207 19669
rect 11238 19660 11244 19712
rect 11296 19700 11302 19712
rect 11609 19703 11667 19709
rect 11296 19672 11341 19700
rect 11296 19660 11302 19672
rect 11609 19669 11621 19703
rect 11655 19700 11667 19703
rect 11974 19700 11980 19712
rect 11655 19672 11980 19700
rect 11655 19669 11667 19672
rect 11609 19663 11667 19669
rect 11974 19660 11980 19672
rect 12032 19660 12038 19712
rect 13725 19703 13783 19709
rect 13725 19669 13737 19703
rect 13771 19700 13783 19703
rect 13814 19700 13820 19712
rect 13771 19672 13820 19700
rect 13771 19669 13783 19672
rect 13725 19663 13783 19669
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 15746 19700 15752 19712
rect 15707 19672 15752 19700
rect 15746 19660 15752 19672
rect 15804 19660 15810 19712
rect 15838 19660 15844 19712
rect 15896 19700 15902 19712
rect 16025 19703 16083 19709
rect 16025 19700 16037 19703
rect 15896 19672 16037 19700
rect 15896 19660 15902 19672
rect 16025 19669 16037 19672
rect 16071 19669 16083 19703
rect 16390 19700 16396 19712
rect 16351 19672 16396 19700
rect 16025 19663 16083 19669
rect 16390 19660 16396 19672
rect 16448 19660 16454 19712
rect 17034 19700 17040 19712
rect 16995 19672 17040 19700
rect 17034 19660 17040 19672
rect 17092 19660 17098 19712
rect 17236 19700 17264 19728
rect 17497 19703 17555 19709
rect 17497 19700 17509 19703
rect 17236 19672 17509 19700
rect 17497 19669 17509 19672
rect 17543 19669 17555 19703
rect 17497 19663 17555 19669
rect 17586 19660 17592 19712
rect 17644 19700 17650 19712
rect 18509 19703 18567 19709
rect 18509 19700 18521 19703
rect 17644 19672 18521 19700
rect 17644 19660 17650 19672
rect 18509 19669 18521 19672
rect 18555 19669 18567 19703
rect 18509 19663 18567 19669
rect 18598 19660 18604 19712
rect 18656 19700 18662 19712
rect 19521 19703 19579 19709
rect 19521 19700 19533 19703
rect 18656 19672 19533 19700
rect 18656 19660 18662 19672
rect 19521 19669 19533 19672
rect 19567 19669 19579 19703
rect 19521 19663 19579 19669
rect 19613 19703 19671 19709
rect 19613 19669 19625 19703
rect 19659 19700 19671 19703
rect 19978 19700 19984 19712
rect 19659 19672 19984 19700
rect 19659 19669 19671 19672
rect 19613 19663 19671 19669
rect 19978 19660 19984 19672
rect 20036 19660 20042 19712
rect 21266 19700 21272 19712
rect 21227 19672 21272 19700
rect 21266 19660 21272 19672
rect 21324 19660 21330 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 3973 19499 4031 19505
rect 3973 19465 3985 19499
rect 4019 19496 4031 19499
rect 4614 19496 4620 19508
rect 4019 19468 4620 19496
rect 4019 19465 4031 19468
rect 3973 19459 4031 19465
rect 4614 19456 4620 19468
rect 4672 19456 4678 19508
rect 5350 19496 5356 19508
rect 5311 19468 5356 19496
rect 5350 19456 5356 19468
rect 5408 19456 5414 19508
rect 7745 19499 7803 19505
rect 7745 19465 7757 19499
rect 7791 19496 7803 19499
rect 10042 19496 10048 19508
rect 7791 19468 10048 19496
rect 7791 19465 7803 19468
rect 7745 19459 7803 19465
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 10594 19496 10600 19508
rect 10555 19468 10600 19496
rect 10594 19456 10600 19468
rect 10652 19456 10658 19508
rect 11238 19456 11244 19508
rect 11296 19496 11302 19508
rect 13081 19499 13139 19505
rect 13081 19496 13093 19499
rect 11296 19468 13093 19496
rect 11296 19456 11302 19468
rect 13081 19465 13093 19468
rect 13127 19465 13139 19499
rect 13446 19496 13452 19508
rect 13407 19468 13452 19496
rect 13081 19459 13139 19465
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 15197 19499 15255 19505
rect 15197 19465 15209 19499
rect 15243 19496 15255 19499
rect 15838 19496 15844 19508
rect 15243 19468 15844 19496
rect 15243 19465 15255 19468
rect 15197 19459 15255 19465
rect 15838 19456 15844 19468
rect 15896 19456 15902 19508
rect 16025 19499 16083 19505
rect 16025 19465 16037 19499
rect 16071 19496 16083 19499
rect 16390 19496 16396 19508
rect 16071 19468 16396 19496
rect 16071 19465 16083 19468
rect 16025 19459 16083 19465
rect 16390 19456 16396 19468
rect 16448 19456 16454 19508
rect 17405 19499 17463 19505
rect 16776 19468 17080 19496
rect 2682 19428 2688 19440
rect 1688 19400 2688 19428
rect 1688 19369 1716 19400
rect 2682 19388 2688 19400
rect 2740 19388 2746 19440
rect 3142 19388 3148 19440
rect 3200 19428 3206 19440
rect 5445 19431 5503 19437
rect 5445 19428 5457 19431
rect 3200 19400 5457 19428
rect 3200 19388 3206 19400
rect 5445 19397 5457 19400
rect 5491 19397 5503 19431
rect 9950 19428 9956 19440
rect 9863 19400 9956 19428
rect 5445 19391 5503 19397
rect 9950 19388 9956 19400
rect 10008 19428 10014 19440
rect 10505 19431 10563 19437
rect 10505 19428 10517 19431
rect 10008 19400 10517 19428
rect 10008 19388 10014 19400
rect 10505 19397 10517 19400
rect 10551 19428 10563 19431
rect 16776 19428 16804 19468
rect 16942 19428 16948 19440
rect 10551 19400 12434 19428
rect 10551 19397 10563 19400
rect 10505 19391 10563 19397
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19329 1731 19363
rect 2222 19360 2228 19372
rect 2183 19332 2228 19360
rect 1673 19323 1731 19329
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 2498 19360 2504 19372
rect 2459 19332 2504 19360
rect 2498 19320 2504 19332
rect 2556 19320 2562 19372
rect 3418 19320 3424 19372
rect 3476 19360 3482 19372
rect 3513 19363 3571 19369
rect 3513 19360 3525 19363
rect 3476 19332 3525 19360
rect 3476 19320 3482 19332
rect 3513 19329 3525 19332
rect 3559 19329 3571 19363
rect 3513 19323 3571 19329
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 4246 19360 4252 19372
rect 3651 19332 4252 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 4246 19320 4252 19332
rect 4304 19320 4310 19372
rect 6730 19320 6736 19372
rect 6788 19360 6794 19372
rect 7377 19363 7435 19369
rect 7377 19360 7389 19363
rect 6788 19332 7389 19360
rect 6788 19320 6794 19332
rect 7377 19329 7389 19332
rect 7423 19360 7435 19363
rect 11790 19360 11796 19372
rect 7423 19332 8524 19360
rect 7423 19329 7435 19332
rect 7377 19323 7435 19329
rect 3329 19295 3387 19301
rect 3329 19261 3341 19295
rect 3375 19261 3387 19295
rect 5626 19292 5632 19304
rect 5587 19264 5632 19292
rect 3329 19255 3387 19261
rect 2038 19224 2044 19236
rect 1999 19196 2044 19224
rect 2038 19184 2044 19196
rect 2096 19184 2102 19236
rect 3344 19224 3372 19255
rect 5626 19252 5632 19264
rect 5684 19252 5690 19304
rect 7193 19295 7251 19301
rect 7193 19261 7205 19295
rect 7239 19261 7251 19295
rect 7193 19255 7251 19261
rect 7285 19295 7343 19301
rect 7285 19261 7297 19295
rect 7331 19292 7343 19295
rect 7926 19292 7932 19304
rect 7331 19264 7932 19292
rect 7331 19261 7343 19264
rect 7285 19255 7343 19261
rect 4338 19224 4344 19236
rect 3344 19196 4344 19224
rect 4338 19184 4344 19196
rect 4396 19224 4402 19236
rect 4709 19227 4767 19233
rect 4709 19224 4721 19227
rect 4396 19196 4721 19224
rect 4396 19184 4402 19196
rect 4709 19193 4721 19196
rect 4755 19224 4767 19227
rect 7208 19224 7236 19255
rect 7926 19252 7932 19264
rect 7984 19252 7990 19304
rect 8386 19292 8392 19304
rect 8347 19264 8392 19292
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 8496 19292 8524 19332
rect 10244 19332 10548 19360
rect 11751 19332 11796 19360
rect 10244 19292 10272 19332
rect 10410 19292 10416 19304
rect 8496 19264 10272 19292
rect 10371 19264 10416 19292
rect 10410 19252 10416 19264
rect 10468 19252 10474 19304
rect 10520 19292 10548 19332
rect 11790 19320 11796 19332
rect 11848 19320 11854 19372
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19329 11943 19363
rect 12406 19360 12434 19400
rect 12728 19400 16804 19428
rect 16903 19400 16948 19428
rect 12526 19360 12532 19372
rect 12406 19332 12532 19360
rect 11885 19323 11943 19329
rect 11238 19292 11244 19304
rect 10520 19264 11244 19292
rect 11238 19252 11244 19264
rect 11296 19252 11302 19304
rect 11701 19295 11759 19301
rect 11701 19261 11713 19295
rect 11747 19261 11759 19295
rect 11900 19292 11928 19323
rect 12526 19320 12532 19332
rect 12584 19320 12590 19372
rect 11974 19292 11980 19304
rect 11900 19264 11980 19292
rect 11701 19255 11759 19261
rect 7558 19224 7564 19236
rect 4755 19196 7144 19224
rect 7208 19196 7564 19224
rect 4755 19193 4767 19196
rect 4709 19187 4767 19193
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 2685 19159 2743 19165
rect 2685 19125 2697 19159
rect 2731 19156 2743 19159
rect 3050 19156 3056 19168
rect 2731 19128 3056 19156
rect 2731 19125 2743 19128
rect 2685 19119 2743 19125
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 4982 19156 4988 19168
rect 4943 19128 4988 19156
rect 4982 19116 4988 19128
rect 5040 19116 5046 19168
rect 6730 19156 6736 19168
rect 6691 19128 6736 19156
rect 6730 19116 6736 19128
rect 6788 19116 6794 19168
rect 7116 19156 7144 19196
rect 7558 19184 7564 19196
rect 7616 19224 7622 19236
rect 8941 19227 8999 19233
rect 8941 19224 8953 19227
rect 7616 19196 8953 19224
rect 7616 19184 7622 19196
rect 8941 19193 8953 19196
rect 8987 19224 8999 19227
rect 11716 19224 11744 19255
rect 11974 19252 11980 19264
rect 12032 19252 12038 19304
rect 12728 19292 12756 19400
rect 16942 19388 16948 19400
rect 17000 19388 17006 19440
rect 17052 19428 17080 19468
rect 17405 19465 17417 19499
rect 17451 19496 17463 19499
rect 17494 19496 17500 19508
rect 17451 19468 17500 19496
rect 17451 19465 17463 19468
rect 17405 19459 17463 19465
rect 17494 19456 17500 19468
rect 17552 19456 17558 19508
rect 18230 19496 18236 19508
rect 18191 19468 18236 19496
rect 18230 19456 18236 19468
rect 18288 19456 18294 19508
rect 18325 19499 18383 19505
rect 18325 19465 18337 19499
rect 18371 19496 18383 19499
rect 19058 19496 19064 19508
rect 18371 19468 19064 19496
rect 18371 19465 18383 19468
rect 18325 19459 18383 19465
rect 19058 19456 19064 19468
rect 19116 19456 19122 19508
rect 19613 19499 19671 19505
rect 19613 19465 19625 19499
rect 19659 19496 19671 19499
rect 19794 19496 19800 19508
rect 19659 19468 19800 19496
rect 19659 19465 19671 19468
rect 19613 19459 19671 19465
rect 19794 19456 19800 19468
rect 19852 19456 19858 19508
rect 19978 19496 19984 19508
rect 19939 19468 19984 19496
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 20717 19499 20775 19505
rect 20717 19496 20729 19499
rect 20680 19468 20729 19496
rect 20680 19456 20686 19468
rect 20717 19465 20729 19468
rect 20763 19465 20775 19499
rect 20717 19459 20775 19465
rect 20806 19428 20812 19440
rect 17052 19400 20812 19428
rect 20806 19388 20812 19400
rect 20864 19388 20870 19440
rect 14274 19360 14280 19372
rect 12912 19332 14280 19360
rect 12912 19304 12940 19332
rect 14274 19320 14280 19332
rect 14332 19320 14338 19372
rect 15194 19360 15200 19372
rect 14936 19332 15200 19360
rect 12728 19264 12848 19292
rect 11882 19224 11888 19236
rect 8987 19196 11652 19224
rect 11716 19196 11888 19224
rect 8987 19193 8999 19196
rect 8941 19187 8999 19193
rect 7742 19156 7748 19168
rect 7116 19128 7748 19156
rect 7742 19116 7748 19128
rect 7800 19116 7806 19168
rect 7926 19116 7932 19168
rect 7984 19156 7990 19168
rect 8021 19159 8079 19165
rect 8021 19156 8033 19159
rect 7984 19128 8033 19156
rect 7984 19116 7990 19128
rect 8021 19125 8033 19128
rect 8067 19125 8079 19159
rect 9214 19156 9220 19168
rect 9175 19128 9220 19156
rect 8021 19119 8079 19125
rect 9214 19116 9220 19128
rect 9272 19116 9278 19168
rect 10962 19156 10968 19168
rect 10923 19128 10968 19156
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 11624 19156 11652 19196
rect 11882 19184 11888 19196
rect 11940 19184 11946 19236
rect 12250 19224 12256 19236
rect 12211 19196 12256 19224
rect 12250 19184 12256 19196
rect 12308 19184 12314 19236
rect 12434 19156 12440 19168
rect 11624 19128 12440 19156
rect 12434 19116 12440 19128
rect 12492 19116 12498 19168
rect 12713 19159 12771 19165
rect 12713 19125 12725 19159
rect 12759 19156 12771 19159
rect 12820 19156 12848 19264
rect 12894 19252 12900 19304
rect 12952 19252 12958 19304
rect 13538 19292 13544 19304
rect 13499 19264 13544 19292
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19261 13691 19295
rect 13633 19255 13691 19261
rect 14185 19295 14243 19301
rect 14185 19261 14197 19295
rect 14231 19292 14243 19295
rect 14936 19292 14964 19332
rect 15194 19320 15200 19332
rect 15252 19360 15258 19372
rect 15378 19360 15384 19372
rect 15252 19332 15384 19360
rect 15252 19320 15258 19332
rect 15378 19320 15384 19332
rect 15436 19320 15442 19372
rect 17037 19363 17095 19369
rect 17037 19360 17049 19363
rect 15580 19332 17049 19360
rect 14231 19264 14964 19292
rect 15013 19295 15071 19301
rect 14231 19261 14243 19264
rect 14185 19255 14243 19261
rect 15013 19261 15025 19295
rect 15059 19261 15071 19295
rect 15013 19255 15071 19261
rect 15105 19295 15163 19301
rect 15105 19261 15117 19295
rect 15151 19292 15163 19295
rect 15470 19292 15476 19304
rect 15151 19264 15476 19292
rect 15151 19261 15163 19264
rect 15105 19255 15163 19261
rect 13446 19184 13452 19236
rect 13504 19224 13510 19236
rect 13648 19224 13676 19255
rect 13504 19196 13676 19224
rect 14553 19227 14611 19233
rect 13504 19184 13510 19196
rect 14553 19193 14565 19227
rect 14599 19224 14611 19227
rect 15028 19224 15056 19255
rect 15470 19252 15476 19264
rect 15528 19252 15534 19304
rect 15580 19233 15608 19332
rect 17037 19329 17049 19332
rect 17083 19329 17095 19363
rect 17037 19323 17095 19329
rect 18874 19320 18880 19372
rect 18932 19360 18938 19372
rect 20533 19363 20591 19369
rect 20533 19360 20545 19363
rect 18932 19332 20545 19360
rect 18932 19320 18938 19332
rect 20533 19329 20545 19332
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 20714 19320 20720 19372
rect 20772 19360 20778 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20772 19332 21097 19360
rect 20772 19320 20778 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 16853 19295 16911 19301
rect 16853 19261 16865 19295
rect 16899 19292 16911 19295
rect 17126 19292 17132 19304
rect 16899 19264 17132 19292
rect 16899 19261 16911 19264
rect 16853 19255 16911 19261
rect 17126 19252 17132 19264
rect 17184 19252 17190 19304
rect 18417 19295 18475 19301
rect 18417 19261 18429 19295
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 19429 19295 19487 19301
rect 19429 19261 19441 19295
rect 19475 19261 19487 19295
rect 19429 19255 19487 19261
rect 19521 19295 19579 19301
rect 19521 19261 19533 19295
rect 19567 19292 19579 19295
rect 19610 19292 19616 19304
rect 19567 19264 19616 19292
rect 19567 19261 19579 19264
rect 19521 19255 19579 19261
rect 15565 19227 15623 19233
rect 14599 19196 15139 19224
rect 14599 19193 14611 19196
rect 14553 19187 14611 19193
rect 12759 19128 12848 19156
rect 15111 19156 15139 19196
rect 15565 19193 15577 19227
rect 15611 19193 15623 19227
rect 15565 19187 15623 19193
rect 18046 19184 18052 19236
rect 18104 19224 18110 19236
rect 18432 19224 18460 19255
rect 18104 19196 18460 19224
rect 19444 19224 19472 19255
rect 19610 19252 19616 19264
rect 19668 19252 19674 19304
rect 21542 19224 21548 19236
rect 19444 19196 21548 19224
rect 18104 19184 18110 19196
rect 21542 19184 21548 19196
rect 21600 19184 21606 19236
rect 16298 19156 16304 19168
rect 15111 19128 16304 19156
rect 12759 19125 12771 19128
rect 12713 19119 12771 19125
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 17862 19156 17868 19168
rect 17823 19128 17868 19156
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 18506 19116 18512 19168
rect 18564 19156 18570 19168
rect 18877 19159 18935 19165
rect 18877 19156 18889 19159
rect 18564 19128 18889 19156
rect 18564 19116 18570 19128
rect 18877 19125 18889 19128
rect 18923 19156 18935 19159
rect 19610 19156 19616 19168
rect 18923 19128 19616 19156
rect 18923 19125 18935 19128
rect 18877 19119 18935 19125
rect 19610 19116 19616 19128
rect 19668 19116 19674 19168
rect 21269 19159 21327 19165
rect 21269 19125 21281 19159
rect 21315 19156 21327 19159
rect 21358 19156 21364 19168
rect 21315 19128 21364 19156
rect 21315 19125 21327 19128
rect 21269 19119 21327 19125
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 2222 18912 2228 18964
rect 2280 18952 2286 18964
rect 2409 18955 2467 18961
rect 2409 18952 2421 18955
rect 2280 18924 2421 18952
rect 2280 18912 2286 18924
rect 2409 18921 2421 18924
rect 2455 18921 2467 18955
rect 2409 18915 2467 18921
rect 2498 18912 2504 18964
rect 2556 18952 2562 18964
rect 4525 18955 4583 18961
rect 4525 18952 4537 18955
rect 2556 18924 4537 18952
rect 2556 18912 2562 18924
rect 4525 18921 4537 18924
rect 4571 18921 4583 18955
rect 4525 18915 4583 18921
rect 5074 18912 5080 18964
rect 5132 18952 5138 18964
rect 9950 18952 9956 18964
rect 5132 18924 9956 18952
rect 5132 18912 5138 18924
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10410 18912 10416 18964
rect 10468 18952 10474 18964
rect 11701 18955 11759 18961
rect 11701 18952 11713 18955
rect 10468 18924 11713 18952
rect 10468 18912 10474 18924
rect 11701 18921 11713 18924
rect 11747 18921 11759 18955
rect 11701 18915 11759 18921
rect 12437 18955 12495 18961
rect 12437 18921 12449 18955
rect 12483 18952 12495 18955
rect 12526 18952 12532 18964
rect 12483 18924 12532 18952
rect 12483 18921 12495 18924
rect 12437 18915 12495 18921
rect 12526 18912 12532 18924
rect 12584 18912 12590 18964
rect 12618 18912 12624 18964
rect 12676 18952 12682 18964
rect 14734 18952 14740 18964
rect 12676 18924 14740 18952
rect 12676 18912 12682 18924
rect 14734 18912 14740 18924
rect 14792 18912 14798 18964
rect 15470 18952 15476 18964
rect 15431 18924 15476 18952
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 15562 18912 15568 18964
rect 15620 18952 15626 18964
rect 18506 18952 18512 18964
rect 15620 18924 18512 18952
rect 15620 18912 15626 18924
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 18874 18952 18880 18964
rect 18835 18924 18880 18952
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 20530 18952 20536 18964
rect 19392 18924 20536 18952
rect 19392 18912 19398 18924
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 1670 18844 1676 18896
rect 1728 18884 1734 18896
rect 2869 18887 2927 18893
rect 2869 18884 2881 18887
rect 1728 18856 2881 18884
rect 1728 18844 1734 18856
rect 2869 18853 2881 18856
rect 2915 18853 2927 18887
rect 2869 18847 2927 18853
rect 3881 18887 3939 18893
rect 3881 18853 3893 18887
rect 3927 18884 3939 18887
rect 4706 18884 4712 18896
rect 3927 18856 4712 18884
rect 3927 18853 3939 18856
rect 3881 18847 3939 18853
rect 3896 18816 3924 18847
rect 4706 18844 4712 18856
rect 4764 18844 4770 18896
rect 5629 18887 5687 18893
rect 5629 18884 5641 18887
rect 5184 18856 5641 18884
rect 5184 18825 5212 18856
rect 5629 18853 5641 18856
rect 5675 18884 5687 18887
rect 9674 18884 9680 18896
rect 5675 18856 9435 18884
rect 9635 18856 9680 18884
rect 5675 18853 5687 18856
rect 5629 18847 5687 18853
rect 2608 18788 3924 18816
rect 5169 18819 5227 18825
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18717 1731 18751
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 1673 18711 1731 18717
rect 1688 18680 1716 18711
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 2608 18757 2636 18788
rect 5169 18785 5181 18819
rect 5215 18785 5227 18819
rect 7834 18816 7840 18828
rect 5169 18779 5227 18785
rect 5460 18788 7840 18816
rect 2593 18751 2651 18757
rect 2593 18717 2605 18751
rect 2639 18717 2651 18751
rect 3050 18748 3056 18760
rect 3011 18720 3056 18748
rect 2593 18711 2651 18717
rect 3050 18708 3056 18720
rect 3108 18708 3114 18760
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18748 4951 18751
rect 4982 18748 4988 18760
rect 4939 18720 4988 18748
rect 4939 18717 4951 18720
rect 4893 18711 4951 18717
rect 4982 18708 4988 18720
rect 5040 18708 5046 18760
rect 2774 18680 2780 18692
rect 1688 18652 2780 18680
rect 2774 18640 2780 18652
rect 2832 18640 2838 18692
rect 5460 18680 5488 18788
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 8021 18819 8079 18825
rect 8021 18785 8033 18819
rect 8067 18816 8079 18819
rect 8662 18816 8668 18828
rect 8067 18788 8668 18816
rect 8067 18785 8079 18788
rect 8021 18779 8079 18785
rect 8662 18776 8668 18788
rect 8720 18776 8726 18828
rect 5626 18708 5632 18760
rect 5684 18748 5690 18760
rect 5997 18751 6055 18757
rect 5997 18748 6009 18751
rect 5684 18720 6009 18748
rect 5684 18708 5690 18720
rect 5997 18717 6009 18720
rect 6043 18748 6055 18751
rect 6546 18748 6552 18760
rect 6043 18720 6552 18748
rect 6043 18717 6055 18720
rect 5997 18711 6055 18717
rect 6546 18708 6552 18720
rect 6604 18708 6610 18760
rect 8205 18751 8263 18757
rect 8205 18717 8217 18751
rect 8251 18748 8263 18751
rect 8386 18748 8392 18760
rect 8251 18720 8392 18748
rect 8251 18717 8263 18720
rect 8205 18711 8263 18717
rect 8386 18708 8392 18720
rect 8444 18708 8450 18760
rect 3344 18652 5488 18680
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 1670 18572 1676 18624
rect 1728 18612 1734 18624
rect 1949 18615 2007 18621
rect 1949 18612 1961 18615
rect 1728 18584 1961 18612
rect 1728 18572 1734 18584
rect 1949 18581 1961 18584
rect 1995 18581 2007 18615
rect 1949 18575 2007 18581
rect 3050 18572 3056 18624
rect 3108 18612 3114 18624
rect 3344 18621 3372 18652
rect 5534 18640 5540 18692
rect 5592 18680 5598 18692
rect 6273 18683 6331 18689
rect 6273 18680 6285 18683
rect 5592 18652 6285 18680
rect 5592 18640 5598 18652
rect 6273 18649 6285 18652
rect 6319 18649 6331 18683
rect 6273 18643 6331 18649
rect 7282 18640 7288 18692
rect 7340 18680 7346 18692
rect 8113 18683 8171 18689
rect 8113 18680 8125 18683
rect 7340 18652 8125 18680
rect 7340 18640 7346 18652
rect 8113 18649 8125 18652
rect 8159 18649 8171 18683
rect 8113 18643 8171 18649
rect 8294 18640 8300 18692
rect 8352 18680 8358 18692
rect 9309 18683 9367 18689
rect 9309 18680 9321 18683
rect 8352 18652 9321 18680
rect 8352 18640 8358 18652
rect 9309 18649 9321 18652
rect 9355 18649 9367 18683
rect 9407 18680 9435 18856
rect 9674 18844 9680 18856
rect 9732 18844 9738 18896
rect 14182 18844 14188 18896
rect 14240 18884 14246 18896
rect 16942 18884 16948 18896
rect 14240 18856 16948 18884
rect 14240 18844 14246 18856
rect 16942 18844 16948 18856
rect 17000 18844 17006 18896
rect 17037 18887 17095 18893
rect 17037 18853 17049 18887
rect 17083 18853 17095 18887
rect 17037 18847 17095 18853
rect 17497 18887 17555 18893
rect 17497 18853 17509 18887
rect 17543 18884 17555 18887
rect 19705 18887 19763 18893
rect 17543 18856 19656 18884
rect 17543 18853 17555 18856
rect 17497 18847 17555 18853
rect 10594 18816 10600 18828
rect 10555 18788 10600 18816
rect 10594 18776 10600 18788
rect 10652 18776 10658 18828
rect 12802 18776 12808 18828
rect 12860 18816 12866 18828
rect 14826 18816 14832 18828
rect 12860 18788 14832 18816
rect 12860 18776 12866 18788
rect 14826 18776 14832 18788
rect 14884 18776 14890 18828
rect 14921 18819 14979 18825
rect 14921 18785 14933 18819
rect 14967 18785 14979 18819
rect 14921 18779 14979 18785
rect 9490 18708 9496 18760
rect 9548 18748 9554 18760
rect 13081 18751 13139 18757
rect 13081 18748 13093 18751
rect 9548 18720 13093 18748
rect 9548 18708 9554 18720
rect 13081 18717 13093 18720
rect 13127 18748 13139 18751
rect 13538 18748 13544 18760
rect 13127 18720 13544 18748
rect 13127 18717 13139 18720
rect 13081 18711 13139 18717
rect 13538 18708 13544 18720
rect 13596 18708 13602 18760
rect 14936 18748 14964 18779
rect 15102 18776 15108 18828
rect 15160 18816 15166 18828
rect 16301 18819 16359 18825
rect 16301 18816 16313 18819
rect 15160 18788 16313 18816
rect 15160 18776 15166 18788
rect 16301 18785 16313 18788
rect 16347 18785 16359 18819
rect 17052 18816 17080 18847
rect 19334 18816 19340 18828
rect 17052 18788 19340 18816
rect 16301 18779 16359 18785
rect 19334 18776 19340 18788
rect 19392 18776 19398 18828
rect 16390 18748 16396 18760
rect 14936 18720 16396 18748
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 17218 18748 17224 18760
rect 16899 18720 17224 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 17218 18708 17224 18720
rect 17276 18708 17282 18760
rect 17313 18751 17371 18757
rect 17313 18717 17325 18751
rect 17359 18748 17371 18751
rect 17586 18748 17592 18760
rect 17359 18720 17592 18748
rect 17359 18717 17371 18720
rect 17313 18711 17371 18717
rect 17586 18708 17592 18720
rect 17644 18708 17650 18760
rect 17773 18751 17831 18757
rect 17773 18717 17785 18751
rect 17819 18748 17831 18751
rect 18414 18748 18420 18760
rect 17819 18720 18276 18748
rect 18375 18720 18420 18748
rect 17819 18717 17831 18720
rect 17773 18711 17831 18717
rect 12802 18680 12808 18692
rect 9407 18652 12808 18680
rect 9309 18643 9367 18649
rect 12802 18640 12808 18652
rect 12860 18640 12866 18692
rect 15105 18683 15163 18689
rect 15105 18680 15117 18683
rect 13648 18652 15117 18680
rect 13648 18624 13676 18652
rect 15105 18649 15117 18652
rect 15151 18680 15163 18683
rect 15933 18683 15991 18689
rect 15933 18680 15945 18683
rect 15151 18652 15945 18680
rect 15151 18649 15163 18652
rect 15105 18643 15163 18649
rect 15933 18649 15945 18652
rect 15979 18680 15991 18683
rect 16114 18680 16120 18692
rect 15979 18652 16120 18680
rect 15979 18649 15991 18652
rect 15933 18643 15991 18649
rect 16114 18640 16120 18652
rect 16172 18640 16178 18692
rect 3329 18615 3387 18621
rect 3329 18612 3341 18615
rect 3108 18584 3341 18612
rect 3108 18572 3114 18584
rect 3329 18581 3341 18584
rect 3375 18581 3387 18615
rect 4246 18612 4252 18624
rect 4159 18584 4252 18612
rect 3329 18575 3387 18581
rect 4246 18572 4252 18584
rect 4304 18612 4310 18624
rect 4890 18612 4896 18624
rect 4304 18584 4896 18612
rect 4304 18572 4310 18584
rect 4890 18572 4896 18584
rect 4948 18572 4954 18624
rect 4985 18615 5043 18621
rect 4985 18581 4997 18615
rect 5031 18612 5043 18615
rect 5810 18612 5816 18624
rect 5031 18584 5816 18612
rect 5031 18581 5043 18584
rect 4985 18575 5043 18581
rect 5810 18572 5816 18584
rect 5868 18572 5874 18624
rect 6638 18612 6644 18624
rect 6599 18584 6644 18612
rect 6638 18572 6644 18584
rect 6696 18572 6702 18624
rect 7006 18612 7012 18624
rect 6967 18584 7012 18612
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 7466 18612 7472 18624
rect 7379 18584 7472 18612
rect 7466 18572 7472 18584
rect 7524 18612 7530 18624
rect 8018 18612 8024 18624
rect 7524 18584 8024 18612
rect 7524 18572 7530 18584
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 8570 18612 8576 18624
rect 8531 18584 8576 18612
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 8938 18612 8944 18624
rect 8899 18584 8944 18612
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 11333 18615 11391 18621
rect 11333 18612 11345 18615
rect 11204 18584 11345 18612
rect 11204 18572 11210 18584
rect 11333 18581 11345 18584
rect 11379 18612 11391 18615
rect 11974 18612 11980 18624
rect 11379 18584 11980 18612
rect 11379 18581 11391 18584
rect 11333 18575 11391 18581
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12713 18615 12771 18621
rect 12713 18581 12725 18615
rect 12759 18612 12771 18615
rect 12894 18612 12900 18624
rect 12759 18584 12900 18612
rect 12759 18581 12771 18584
rect 12713 18575 12771 18581
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 13630 18612 13636 18624
rect 13591 18584 13636 18612
rect 13630 18572 13636 18584
rect 13688 18572 13694 18624
rect 14366 18612 14372 18624
rect 14327 18584 14372 18612
rect 14366 18572 14372 18584
rect 14424 18612 14430 18624
rect 15013 18615 15071 18621
rect 15013 18612 15025 18615
rect 14424 18584 15025 18612
rect 14424 18572 14430 18584
rect 15013 18581 15025 18584
rect 15059 18581 15071 18615
rect 17954 18612 17960 18624
rect 17915 18584 17960 18612
rect 15013 18575 15071 18581
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18248 18621 18276 18720
rect 18414 18708 18420 18720
rect 18472 18708 18478 18760
rect 18690 18748 18696 18760
rect 18651 18720 18696 18748
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 19518 18748 19524 18760
rect 19479 18720 19524 18748
rect 19518 18708 19524 18720
rect 19576 18708 19582 18760
rect 19628 18680 19656 18856
rect 19705 18853 19717 18887
rect 19751 18853 19763 18887
rect 19705 18847 19763 18853
rect 19720 18748 19748 18847
rect 20165 18751 20223 18757
rect 20165 18748 20177 18751
rect 19720 18720 20177 18748
rect 20165 18717 20177 18720
rect 20211 18717 20223 18751
rect 20622 18748 20628 18760
rect 20583 18720 20628 18748
rect 20165 18711 20223 18717
rect 20622 18708 20628 18720
rect 20680 18708 20686 18760
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 21100 18680 21128 18711
rect 19628 18652 21128 18680
rect 18233 18615 18291 18621
rect 18233 18581 18245 18615
rect 18279 18581 18291 18615
rect 19978 18612 19984 18624
rect 19939 18584 19984 18612
rect 18233 18575 18291 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 20070 18572 20076 18624
rect 20128 18612 20134 18624
rect 20441 18615 20499 18621
rect 20441 18612 20453 18615
rect 20128 18584 20453 18612
rect 20128 18572 20134 18584
rect 20441 18581 20453 18584
rect 20487 18581 20499 18615
rect 21266 18612 21272 18624
rect 21227 18584 21272 18612
rect 20441 18575 20499 18581
rect 21266 18572 21272 18584
rect 21324 18572 21330 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 2130 18408 2136 18420
rect 2091 18380 2136 18408
rect 2130 18368 2136 18380
rect 2188 18368 2194 18420
rect 2409 18411 2467 18417
rect 2409 18377 2421 18411
rect 2455 18377 2467 18411
rect 2409 18371 2467 18377
rect 2424 18340 2452 18371
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 2869 18411 2927 18417
rect 2869 18408 2881 18411
rect 2832 18380 2881 18408
rect 2832 18368 2838 18380
rect 2869 18377 2881 18380
rect 2915 18377 2927 18411
rect 2869 18371 2927 18377
rect 4522 18368 4528 18420
rect 4580 18408 4586 18420
rect 4709 18411 4767 18417
rect 4709 18408 4721 18411
rect 4580 18380 4721 18408
rect 4580 18368 4586 18380
rect 4709 18377 4721 18380
rect 4755 18377 4767 18411
rect 4709 18371 4767 18377
rect 6917 18411 6975 18417
rect 6917 18377 6929 18411
rect 6963 18408 6975 18411
rect 7653 18411 7711 18417
rect 7653 18408 7665 18411
rect 6963 18380 7665 18408
rect 6963 18377 6975 18380
rect 6917 18371 6975 18377
rect 7653 18377 7665 18380
rect 7699 18377 7711 18411
rect 7653 18371 7711 18377
rect 8570 18368 8576 18420
rect 8628 18408 8634 18420
rect 9953 18411 10011 18417
rect 9953 18408 9965 18411
rect 8628 18380 9965 18408
rect 8628 18368 8634 18380
rect 9953 18377 9965 18380
rect 9999 18377 10011 18411
rect 9953 18371 10011 18377
rect 10134 18368 10140 18420
rect 10192 18408 10198 18420
rect 10597 18411 10655 18417
rect 10597 18408 10609 18411
rect 10192 18380 10609 18408
rect 10192 18368 10198 18380
rect 10597 18377 10609 18380
rect 10643 18377 10655 18411
rect 10597 18371 10655 18377
rect 11238 18368 11244 18420
rect 11296 18408 11302 18420
rect 11974 18408 11980 18420
rect 11296 18380 11980 18408
rect 11296 18368 11302 18380
rect 11974 18368 11980 18380
rect 12032 18368 12038 18420
rect 12802 18408 12808 18420
rect 12763 18380 12808 18408
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 13449 18411 13507 18417
rect 13449 18377 13461 18411
rect 13495 18408 13507 18411
rect 15105 18411 15163 18417
rect 15105 18408 15117 18411
rect 13495 18380 15117 18408
rect 13495 18377 13507 18380
rect 13449 18371 13507 18377
rect 15105 18377 15117 18380
rect 15151 18377 15163 18411
rect 15105 18371 15163 18377
rect 15473 18411 15531 18417
rect 15473 18377 15485 18411
rect 15519 18408 15531 18411
rect 15746 18408 15752 18420
rect 15519 18380 15752 18408
rect 15519 18377 15531 18380
rect 15473 18371 15531 18377
rect 15746 18368 15752 18380
rect 15804 18368 15810 18420
rect 16301 18411 16359 18417
rect 16301 18377 16313 18411
rect 16347 18408 16359 18411
rect 18601 18411 18659 18417
rect 16347 18380 17080 18408
rect 16347 18377 16359 18380
rect 16301 18371 16359 18377
rect 4614 18340 4620 18352
rect 1688 18312 2452 18340
rect 4575 18312 4620 18340
rect 1688 18281 1716 18312
rect 4614 18300 4620 18312
rect 4672 18300 4678 18352
rect 7006 18300 7012 18352
rect 7064 18340 7070 18352
rect 8021 18343 8079 18349
rect 8021 18340 8033 18343
rect 7064 18312 8033 18340
rect 7064 18300 7070 18312
rect 8021 18309 8033 18312
rect 8067 18309 8079 18343
rect 8021 18303 8079 18309
rect 8202 18300 8208 18352
rect 8260 18340 8266 18352
rect 9033 18343 9091 18349
rect 9033 18340 9045 18343
rect 8260 18312 9045 18340
rect 8260 18300 8266 18312
rect 9033 18309 9045 18312
rect 9079 18309 9091 18343
rect 9033 18303 9091 18309
rect 10042 18300 10048 18352
rect 10100 18340 10106 18352
rect 14369 18343 14427 18349
rect 14369 18340 14381 18343
rect 10100 18312 14381 18340
rect 10100 18300 10106 18312
rect 14369 18309 14381 18312
rect 14415 18309 14427 18343
rect 14369 18303 14427 18309
rect 15565 18343 15623 18349
rect 15565 18309 15577 18343
rect 15611 18340 15623 18343
rect 15654 18340 15660 18352
rect 15611 18312 15660 18340
rect 15611 18309 15623 18312
rect 15565 18303 15623 18309
rect 15654 18300 15660 18312
rect 15712 18300 15718 18352
rect 17052 18340 17080 18380
rect 18601 18377 18613 18411
rect 18647 18408 18659 18411
rect 19518 18408 19524 18420
rect 18647 18380 19524 18408
rect 18647 18377 18659 18380
rect 18601 18371 18659 18377
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 19889 18411 19947 18417
rect 19889 18377 19901 18411
rect 19935 18408 19947 18411
rect 20990 18408 20996 18420
rect 19935 18380 20996 18408
rect 19935 18377 19947 18380
rect 19889 18371 19947 18377
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 17052 18312 21128 18340
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 1946 18272 1952 18284
rect 1907 18244 1952 18272
rect 1673 18235 1731 18241
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 2593 18275 2651 18281
rect 2593 18241 2605 18275
rect 2639 18272 2651 18275
rect 2958 18272 2964 18284
rect 2639 18244 2964 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 3050 18232 3056 18284
rect 3108 18272 3114 18284
rect 6825 18275 6883 18281
rect 3108 18244 3153 18272
rect 3108 18232 3114 18244
rect 6825 18241 6837 18275
rect 6871 18272 6883 18275
rect 7558 18272 7564 18284
rect 6871 18244 7564 18272
rect 6871 18241 6883 18244
rect 6825 18235 6883 18241
rect 7558 18232 7564 18244
rect 7616 18232 7622 18284
rect 7742 18232 7748 18284
rect 7800 18272 7806 18284
rect 7800 18244 8340 18272
rect 7800 18232 7806 18244
rect 4525 18207 4583 18213
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 7101 18207 7159 18213
rect 7101 18204 7113 18207
rect 4571 18176 7113 18204
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 7101 18173 7113 18176
rect 7147 18173 7159 18207
rect 8110 18204 8116 18216
rect 8071 18176 8116 18204
rect 7101 18167 7159 18173
rect 5077 18139 5135 18145
rect 5077 18105 5089 18139
rect 5123 18136 5135 18139
rect 5626 18136 5632 18148
rect 5123 18108 5632 18136
rect 5123 18105 5135 18108
rect 5077 18099 5135 18105
rect 5626 18096 5632 18108
rect 5684 18096 5690 18148
rect 7116 18136 7144 18167
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 8312 18213 8340 18244
rect 9122 18232 9128 18284
rect 9180 18272 9186 18284
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 9180 18244 12449 18272
rect 9180 18232 9186 18244
rect 12437 18241 12449 18244
rect 12483 18272 12495 18275
rect 14458 18272 14464 18284
rect 12483 18244 14320 18272
rect 14419 18244 14464 18272
rect 12483 18241 12495 18244
rect 12437 18235 12495 18241
rect 8297 18207 8355 18213
rect 8297 18173 8309 18207
rect 8343 18204 8355 18207
rect 8570 18204 8576 18216
rect 8343 18176 8576 18204
rect 8343 18173 8355 18176
rect 8297 18167 8355 18173
rect 8570 18164 8576 18176
rect 8628 18204 8634 18216
rect 8938 18204 8944 18216
rect 8628 18176 8944 18204
rect 8628 18164 8634 18176
rect 8938 18164 8944 18176
rect 8996 18164 9002 18216
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18173 9735 18207
rect 9858 18204 9864 18216
rect 9819 18176 9864 18204
rect 9677 18167 9735 18173
rect 9692 18136 9720 18167
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 13170 18204 13176 18216
rect 13131 18176 13176 18204
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 13354 18204 13360 18216
rect 13315 18176 13360 18204
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 14182 18204 14188 18216
rect 14143 18176 14188 18204
rect 14182 18164 14188 18176
rect 14240 18164 14246 18216
rect 14292 18204 14320 18244
rect 14458 18232 14464 18244
rect 14516 18232 14522 18284
rect 15102 18232 15108 18284
rect 15160 18272 15166 18284
rect 16114 18272 16120 18284
rect 15160 18244 15700 18272
rect 16075 18244 16120 18272
rect 15160 18232 15166 18244
rect 15562 18204 15568 18216
rect 14292 18176 15568 18204
rect 15562 18164 15568 18176
rect 15620 18164 15626 18216
rect 15672 18213 15700 18244
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18241 17371 18275
rect 17313 18235 17371 18241
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18173 15715 18207
rect 15657 18167 15715 18173
rect 17037 18207 17095 18213
rect 17037 18173 17049 18207
rect 17083 18204 17095 18207
rect 17328 18204 17356 18235
rect 17402 18232 17408 18284
rect 17460 18272 17466 18284
rect 18233 18275 18291 18281
rect 18233 18272 18245 18275
rect 17460 18244 18245 18272
rect 17460 18232 17466 18244
rect 18233 18241 18245 18244
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 18322 18232 18328 18284
rect 18380 18272 18386 18284
rect 18877 18275 18935 18281
rect 18877 18272 18889 18275
rect 18380 18244 18889 18272
rect 18380 18232 18386 18244
rect 18877 18241 18889 18244
rect 18923 18241 18935 18275
rect 18877 18235 18935 18241
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19245 18275 19303 18281
rect 19245 18272 19257 18275
rect 19116 18244 19257 18272
rect 19116 18232 19122 18244
rect 19245 18241 19257 18244
rect 19291 18241 19303 18275
rect 19245 18235 19303 18241
rect 19705 18275 19763 18281
rect 19705 18241 19717 18275
rect 19751 18272 19763 18275
rect 20070 18272 20076 18284
rect 19751 18244 20076 18272
rect 19751 18241 19763 18244
rect 19705 18235 19763 18241
rect 20070 18232 20076 18244
rect 20128 18232 20134 18284
rect 20162 18232 20168 18284
rect 20220 18272 20226 18284
rect 20806 18272 20812 18284
rect 20220 18244 20265 18272
rect 20767 18244 20812 18272
rect 20220 18232 20226 18244
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 21100 18281 21128 18312
rect 21085 18275 21143 18281
rect 21085 18241 21097 18275
rect 21131 18241 21143 18275
rect 21085 18235 21143 18241
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17083 18176 18061 18204
rect 17083 18173 17095 18176
rect 17037 18167 17095 18173
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 18141 18207 18199 18213
rect 18141 18173 18153 18207
rect 18187 18204 18199 18207
rect 19518 18204 19524 18216
rect 18187 18176 19524 18204
rect 18187 18173 18199 18176
rect 18141 18167 18199 18173
rect 9766 18136 9772 18148
rect 7116 18108 8800 18136
rect 9692 18108 9772 18136
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 3234 18028 3240 18080
rect 3292 18068 3298 18080
rect 3329 18071 3387 18077
rect 3329 18068 3341 18071
rect 3292 18040 3341 18068
rect 3292 18028 3298 18040
rect 3329 18037 3341 18040
rect 3375 18037 3387 18071
rect 3329 18031 3387 18037
rect 3789 18071 3847 18077
rect 3789 18037 3801 18071
rect 3835 18068 3847 18071
rect 3970 18068 3976 18080
rect 3835 18040 3976 18068
rect 3835 18037 3847 18040
rect 3789 18031 3847 18037
rect 3970 18028 3976 18040
rect 4028 18028 4034 18080
rect 5350 18068 5356 18080
rect 5311 18040 5356 18068
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 5718 18068 5724 18080
rect 5679 18040 5724 18068
rect 5718 18028 5724 18040
rect 5776 18028 5782 18080
rect 5810 18028 5816 18080
rect 5868 18068 5874 18080
rect 6457 18071 6515 18077
rect 6457 18068 6469 18071
rect 5868 18040 6469 18068
rect 5868 18028 5874 18040
rect 6457 18037 6469 18040
rect 6503 18037 6515 18071
rect 6457 18031 6515 18037
rect 8570 18028 8576 18080
rect 8628 18068 8634 18080
rect 8665 18071 8723 18077
rect 8665 18068 8677 18071
rect 8628 18040 8677 18068
rect 8628 18028 8634 18040
rect 8665 18037 8677 18040
rect 8711 18037 8723 18071
rect 8772 18068 8800 18108
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 10321 18139 10379 18145
rect 10321 18105 10333 18139
rect 10367 18136 10379 18139
rect 11790 18136 11796 18148
rect 10367 18108 11796 18136
rect 10367 18105 10379 18108
rect 10321 18099 10379 18105
rect 11790 18096 11796 18108
rect 11848 18096 11854 18148
rect 14829 18139 14887 18145
rect 14829 18105 14841 18139
rect 14875 18136 14887 18139
rect 17402 18136 17408 18148
rect 14875 18108 17408 18136
rect 14875 18105 14887 18108
rect 14829 18099 14887 18105
rect 17402 18096 17408 18108
rect 17460 18096 17466 18148
rect 18064 18136 18092 18167
rect 19518 18164 19524 18176
rect 19576 18164 19582 18216
rect 20714 18204 20720 18216
rect 20272 18176 20720 18204
rect 18322 18136 18328 18148
rect 18064 18108 18328 18136
rect 18322 18096 18328 18108
rect 18380 18096 18386 18148
rect 19429 18139 19487 18145
rect 19429 18105 19441 18139
rect 19475 18136 19487 18139
rect 20272 18136 20300 18176
rect 20714 18164 20720 18176
rect 20772 18164 20778 18216
rect 19475 18108 20300 18136
rect 20349 18139 20407 18145
rect 19475 18105 19487 18108
rect 19429 18099 19487 18105
rect 20349 18105 20361 18139
rect 20395 18136 20407 18139
rect 21082 18136 21088 18148
rect 20395 18108 21088 18136
rect 20395 18105 20407 18108
rect 20349 18099 20407 18105
rect 21082 18096 21088 18108
rect 21140 18096 21146 18148
rect 12066 18068 12072 18080
rect 8772 18040 12072 18068
rect 8665 18031 8723 18037
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 13817 18071 13875 18077
rect 13817 18037 13829 18071
rect 13863 18068 13875 18071
rect 18414 18068 18420 18080
rect 13863 18040 18420 18068
rect 13863 18037 13875 18040
rect 13817 18031 13875 18037
rect 18414 18028 18420 18040
rect 18472 18028 18478 18080
rect 20254 18028 20260 18080
rect 20312 18068 20318 18080
rect 20625 18071 20683 18077
rect 20625 18068 20637 18071
rect 20312 18040 20637 18068
rect 20312 18028 20318 18040
rect 20625 18037 20637 18040
rect 20671 18037 20683 18071
rect 20625 18031 20683 18037
rect 21269 18071 21327 18077
rect 21269 18037 21281 18071
rect 21315 18068 21327 18071
rect 21358 18068 21364 18080
rect 21315 18040 21364 18068
rect 21315 18037 21327 18040
rect 21269 18031 21327 18037
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 14 17824 20 17876
rect 72 17864 78 17876
rect 1026 17864 1032 17876
rect 72 17836 1032 17864
rect 72 17824 78 17836
rect 1026 17824 1032 17836
rect 1084 17824 1090 17876
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 2961 17867 3019 17873
rect 2961 17864 2973 17867
rect 2832 17836 2973 17864
rect 2832 17824 2838 17836
rect 2961 17833 2973 17836
rect 3007 17833 3019 17867
rect 6822 17864 6828 17876
rect 6783 17836 6828 17864
rect 2961 17827 3019 17833
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 7469 17867 7527 17873
rect 7469 17864 7481 17867
rect 7432 17836 7481 17864
rect 7432 17824 7438 17836
rect 7469 17833 7481 17836
rect 7515 17833 7527 17867
rect 7469 17827 7527 17833
rect 7837 17867 7895 17873
rect 7837 17833 7849 17867
rect 7883 17864 7895 17867
rect 8110 17864 8116 17876
rect 7883 17836 8116 17864
rect 7883 17833 7895 17836
rect 7837 17827 7895 17833
rect 8110 17824 8116 17836
rect 8168 17824 8174 17876
rect 8386 17824 8392 17876
rect 8444 17864 8450 17876
rect 11054 17864 11060 17876
rect 8444 17836 11060 17864
rect 8444 17824 8450 17836
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 17218 17864 17224 17876
rect 12406 17836 17224 17864
rect 1854 17756 1860 17808
rect 1912 17796 1918 17808
rect 4062 17796 4068 17808
rect 1912 17768 4068 17796
rect 1912 17756 1918 17768
rect 4062 17756 4068 17768
rect 4120 17756 4126 17808
rect 8754 17756 8760 17808
rect 8812 17796 8818 17808
rect 12406 17796 12434 17836
rect 17218 17824 17224 17836
rect 17276 17864 17282 17876
rect 18230 17864 18236 17876
rect 17276 17836 18236 17864
rect 17276 17824 17282 17836
rect 18230 17824 18236 17836
rect 18288 17824 18294 17876
rect 18414 17864 18420 17876
rect 18375 17836 18420 17864
rect 18414 17824 18420 17836
rect 18472 17824 18478 17876
rect 19337 17867 19395 17873
rect 19337 17833 19349 17867
rect 19383 17864 19395 17867
rect 19518 17864 19524 17876
rect 19383 17836 19524 17864
rect 19383 17833 19395 17836
rect 19337 17827 19395 17833
rect 19518 17824 19524 17836
rect 19576 17824 19582 17876
rect 8812 17768 12434 17796
rect 8812 17756 8818 17768
rect 12526 17756 12532 17808
rect 12584 17796 12590 17808
rect 16114 17796 16120 17808
rect 12584 17768 16120 17796
rect 12584 17756 12590 17768
rect 16114 17756 16120 17768
rect 16172 17756 16178 17808
rect 16390 17756 16396 17808
rect 16448 17796 16454 17808
rect 16577 17799 16635 17805
rect 16577 17796 16589 17799
rect 16448 17768 16589 17796
rect 16448 17756 16454 17768
rect 16577 17765 16589 17768
rect 16623 17796 16635 17799
rect 16623 17768 17264 17796
rect 16623 17765 16635 17768
rect 16577 17759 16635 17765
rect 3970 17728 3976 17740
rect 2700 17700 3976 17728
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17629 1731 17663
rect 2222 17660 2228 17672
rect 2183 17632 2228 17660
rect 1673 17623 1731 17629
rect 1688 17592 1716 17623
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 2700 17669 2728 17700
rect 3970 17688 3976 17700
rect 4028 17688 4034 17740
rect 4617 17731 4675 17737
rect 4617 17697 4629 17731
rect 4663 17728 4675 17731
rect 5350 17728 5356 17740
rect 4663 17700 5356 17728
rect 4663 17697 4675 17700
rect 4617 17691 4675 17697
rect 5350 17688 5356 17700
rect 5408 17688 5414 17740
rect 5442 17688 5448 17740
rect 5500 17728 5506 17740
rect 8386 17728 8392 17740
rect 5500 17700 8392 17728
rect 5500 17688 5506 17700
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 10226 17728 10232 17740
rect 8527 17700 10232 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 10226 17688 10232 17700
rect 10284 17688 10290 17740
rect 10321 17731 10379 17737
rect 10321 17697 10333 17731
rect 10367 17728 10379 17731
rect 10410 17728 10416 17740
rect 10367 17700 10416 17728
rect 10367 17697 10379 17700
rect 10321 17691 10379 17697
rect 10410 17688 10416 17700
rect 10468 17688 10474 17740
rect 11054 17728 11060 17740
rect 11015 17700 11060 17728
rect 11054 17688 11060 17700
rect 11112 17728 11118 17740
rect 11885 17731 11943 17737
rect 11112 17700 11376 17728
rect 11112 17688 11118 17700
rect 2685 17663 2743 17669
rect 2685 17629 2697 17663
rect 2731 17629 2743 17663
rect 2685 17623 2743 17629
rect 3145 17663 3203 17669
rect 3145 17629 3157 17663
rect 3191 17660 3203 17663
rect 3234 17660 3240 17672
rect 3191 17632 3240 17660
rect 3191 17629 3203 17632
rect 3145 17623 3203 17629
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 5261 17663 5319 17669
rect 5261 17629 5273 17663
rect 5307 17660 5319 17663
rect 5721 17663 5779 17669
rect 5721 17660 5733 17663
rect 5307 17632 5733 17660
rect 5307 17629 5319 17632
rect 5261 17623 5319 17629
rect 5721 17629 5733 17632
rect 5767 17660 5779 17663
rect 5994 17660 6000 17672
rect 5767 17632 6000 17660
rect 5767 17629 5779 17632
rect 5721 17623 5779 17629
rect 5994 17620 6000 17632
rect 6052 17620 6058 17672
rect 7374 17620 7380 17672
rect 7432 17660 7438 17672
rect 11348 17669 11376 17700
rect 11885 17697 11897 17731
rect 11931 17728 11943 17731
rect 12710 17728 12716 17740
rect 11931 17700 12388 17728
rect 12671 17700 12716 17728
rect 11931 17697 11943 17700
rect 11885 17691 11943 17697
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7432 17632 8217 17660
rect 7432 17620 7438 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 9401 17663 9459 17669
rect 9401 17629 9413 17663
rect 9447 17660 9459 17663
rect 10045 17663 10103 17669
rect 10045 17660 10057 17663
rect 9447 17632 10057 17660
rect 9447 17629 9459 17632
rect 9401 17623 9459 17629
rect 10045 17629 10057 17632
rect 10091 17660 10103 17663
rect 11333 17663 11391 17669
rect 10091 17632 10916 17660
rect 10091 17629 10103 17632
rect 10045 17623 10103 17629
rect 4341 17595 4399 17601
rect 1688 17564 2544 17592
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 2038 17524 2044 17536
rect 1999 17496 2044 17524
rect 2038 17484 2044 17496
rect 2096 17484 2102 17536
rect 2516 17533 2544 17564
rect 4341 17561 4353 17595
rect 4387 17592 4399 17595
rect 4387 17564 5120 17592
rect 4387 17561 4399 17564
rect 4341 17555 4399 17561
rect 2501 17527 2559 17533
rect 2501 17493 2513 17527
rect 2547 17493 2559 17527
rect 3970 17524 3976 17536
rect 3931 17496 3976 17524
rect 2501 17487 2559 17493
rect 3970 17484 3976 17496
rect 4028 17484 4034 17536
rect 4430 17524 4436 17536
rect 4391 17496 4436 17524
rect 4430 17484 4436 17496
rect 4488 17484 4494 17536
rect 5092 17524 5120 17564
rect 7926 17552 7932 17604
rect 7984 17592 7990 17604
rect 9033 17595 9091 17601
rect 9033 17592 9045 17595
rect 7984 17564 9045 17592
rect 7984 17552 7990 17564
rect 9033 17561 9045 17564
rect 9079 17592 9091 17595
rect 10502 17592 10508 17604
rect 9079 17564 10508 17592
rect 9079 17561 9091 17564
rect 9033 17555 9091 17561
rect 10502 17552 10508 17564
rect 10560 17552 10566 17604
rect 10888 17592 10916 17632
rect 11333 17629 11345 17663
rect 11379 17660 11391 17663
rect 12250 17660 12256 17672
rect 11379 17632 12256 17660
rect 11379 17629 11391 17632
rect 11333 17623 11391 17629
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 12360 17604 12388 17700
rect 12710 17688 12716 17700
rect 12768 17688 12774 17740
rect 15657 17731 15715 17737
rect 15657 17697 15669 17731
rect 15703 17728 15715 17731
rect 15838 17728 15844 17740
rect 15703 17700 15844 17728
rect 15703 17697 15715 17700
rect 15657 17691 15715 17697
rect 15838 17688 15844 17700
rect 15896 17688 15902 17740
rect 17129 17731 17187 17737
rect 17129 17697 17141 17731
rect 17175 17697 17187 17731
rect 17236 17728 17264 17768
rect 17954 17756 17960 17808
rect 18012 17796 18018 17808
rect 18012 17768 21128 17796
rect 18012 17756 18018 17768
rect 18138 17728 18144 17740
rect 17236 17700 18144 17728
rect 17129 17691 17187 17697
rect 12434 17620 12440 17672
rect 12492 17660 12498 17672
rect 14550 17660 14556 17672
rect 12492 17632 14556 17660
rect 12492 17620 12498 17632
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 15013 17663 15071 17669
rect 15013 17660 15025 17663
rect 14936 17632 15025 17660
rect 11974 17592 11980 17604
rect 10888 17564 11980 17592
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 12342 17552 12348 17604
rect 12400 17592 12406 17604
rect 12621 17595 12679 17601
rect 12621 17592 12633 17595
rect 12400 17564 12633 17592
rect 12400 17552 12406 17564
rect 12621 17561 12633 17564
rect 12667 17561 12679 17595
rect 12621 17555 12679 17561
rect 14936 17536 14964 17632
rect 15013 17629 15025 17632
rect 15059 17629 15071 17663
rect 15013 17623 15071 17629
rect 15841 17595 15899 17601
rect 15841 17561 15853 17595
rect 15887 17592 15899 17595
rect 17034 17592 17040 17604
rect 15887 17564 17040 17592
rect 15887 17561 15899 17564
rect 15841 17555 15899 17561
rect 17034 17552 17040 17564
rect 17092 17552 17098 17604
rect 17144 17592 17172 17691
rect 18138 17688 18144 17700
rect 18196 17688 18202 17740
rect 19610 17728 19616 17740
rect 18248 17700 19616 17728
rect 17313 17663 17371 17669
rect 17313 17629 17325 17663
rect 17359 17660 17371 17663
rect 17862 17660 17868 17672
rect 17359 17632 17868 17660
rect 17359 17629 17371 17632
rect 17313 17623 17371 17629
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 18248 17669 18276 17700
rect 19610 17688 19616 17700
rect 19668 17688 19674 17740
rect 19794 17688 19800 17740
rect 19852 17728 19858 17740
rect 19889 17731 19947 17737
rect 19889 17728 19901 17731
rect 19852 17700 19901 17728
rect 19852 17688 19858 17700
rect 19889 17697 19901 17700
rect 19935 17728 19947 17731
rect 20438 17728 20444 17740
rect 19935 17700 20444 17728
rect 19935 17697 19947 17700
rect 19889 17691 19947 17697
rect 20438 17688 20444 17700
rect 20496 17688 20502 17740
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18506 17620 18512 17672
rect 18564 17660 18570 17672
rect 21100 17669 21128 17768
rect 18693 17663 18751 17669
rect 18693 17660 18705 17663
rect 18564 17632 18705 17660
rect 18564 17620 18570 17632
rect 18693 17629 18705 17632
rect 18739 17629 18751 17663
rect 20533 17663 20591 17669
rect 20533 17660 20545 17663
rect 18693 17623 18751 17629
rect 18892 17632 20545 17660
rect 17586 17592 17592 17604
rect 17144 17564 17592 17592
rect 17586 17552 17592 17564
rect 17644 17592 17650 17604
rect 18598 17592 18604 17604
rect 17644 17564 18604 17592
rect 17644 17552 17650 17564
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 6089 17527 6147 17533
rect 6089 17524 6101 17527
rect 5092 17496 6101 17524
rect 6089 17493 6101 17496
rect 6135 17493 6147 17527
rect 6089 17487 6147 17493
rect 7006 17484 7012 17536
rect 7064 17524 7070 17536
rect 7101 17527 7159 17533
rect 7101 17524 7113 17527
rect 7064 17496 7113 17524
rect 7064 17484 7070 17496
rect 7101 17493 7113 17496
rect 7147 17493 7159 17527
rect 7101 17487 7159 17493
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 8202 17524 8208 17536
rect 7432 17496 8208 17524
rect 7432 17484 7438 17496
rect 8202 17484 8208 17496
rect 8260 17524 8266 17536
rect 8297 17527 8355 17533
rect 8297 17524 8309 17527
rect 8260 17496 8309 17524
rect 8260 17484 8266 17496
rect 8297 17493 8309 17496
rect 8343 17493 8355 17527
rect 9674 17524 9680 17536
rect 9635 17496 9680 17524
rect 8297 17487 8355 17493
rect 9674 17484 9680 17496
rect 9732 17484 9738 17536
rect 10134 17524 10140 17536
rect 10095 17496 10140 17524
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 12158 17524 12164 17536
rect 12119 17496 12164 17524
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12529 17527 12587 17533
rect 12529 17493 12541 17527
rect 12575 17524 12587 17527
rect 13173 17527 13231 17533
rect 13173 17524 13185 17527
rect 12575 17496 13185 17524
rect 12575 17493 12587 17496
rect 12529 17487 12587 17493
rect 13173 17493 13185 17496
rect 13219 17493 13231 17527
rect 13173 17487 13231 17493
rect 13538 17484 13544 17536
rect 13596 17524 13602 17536
rect 13633 17527 13691 17533
rect 13633 17524 13645 17527
rect 13596 17496 13645 17524
rect 13596 17484 13602 17496
rect 13633 17493 13645 17496
rect 13679 17493 13691 17527
rect 14366 17524 14372 17536
rect 14327 17496 14372 17524
rect 13633 17487 13691 17493
rect 14366 17484 14372 17496
rect 14424 17524 14430 17536
rect 14642 17524 14648 17536
rect 14424 17496 14648 17524
rect 14424 17484 14430 17496
rect 14642 17484 14648 17496
rect 14700 17484 14706 17536
rect 14737 17527 14795 17533
rect 14737 17493 14749 17527
rect 14783 17524 14795 17527
rect 14918 17524 14924 17536
rect 14783 17496 14924 17524
rect 14783 17493 14795 17496
rect 14737 17487 14795 17493
rect 14918 17484 14924 17496
rect 14976 17484 14982 17536
rect 15194 17524 15200 17536
rect 15155 17496 15200 17524
rect 15194 17484 15200 17496
rect 15252 17484 15258 17536
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 15749 17527 15807 17533
rect 15749 17524 15761 17527
rect 15620 17496 15761 17524
rect 15620 17484 15626 17496
rect 15749 17493 15761 17496
rect 15795 17493 15807 17527
rect 15749 17487 15807 17493
rect 16209 17527 16267 17533
rect 16209 17493 16221 17527
rect 16255 17524 16267 17527
rect 16390 17524 16396 17536
rect 16255 17496 16396 17524
rect 16255 17493 16267 17496
rect 16209 17487 16267 17493
rect 16390 17484 16396 17496
rect 16448 17484 16454 17536
rect 17218 17524 17224 17536
rect 17179 17496 17224 17524
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 17678 17524 17684 17536
rect 17639 17496 17684 17524
rect 17678 17484 17684 17496
rect 17736 17484 17742 17536
rect 18892 17533 18920 17632
rect 20533 17629 20545 17632
rect 20579 17629 20591 17663
rect 20533 17623 20591 17629
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 19702 17592 19708 17604
rect 19663 17564 19708 17592
rect 19702 17552 19708 17564
rect 19760 17552 19766 17604
rect 18877 17527 18935 17533
rect 18877 17493 18889 17527
rect 18923 17493 18935 17527
rect 18877 17487 18935 17493
rect 19797 17527 19855 17533
rect 19797 17493 19809 17527
rect 19843 17524 19855 17527
rect 20346 17524 20352 17536
rect 19843 17496 20352 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 20714 17524 20720 17536
rect 20675 17496 20720 17524
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 21269 17527 21327 17533
rect 21269 17493 21281 17527
rect 21315 17524 21327 17527
rect 21450 17524 21456 17536
rect 21315 17496 21456 17524
rect 21315 17493 21327 17496
rect 21269 17487 21327 17493
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1946 17280 1952 17332
rect 2004 17320 2010 17332
rect 2317 17323 2375 17329
rect 2317 17320 2329 17323
rect 2004 17292 2329 17320
rect 2004 17280 2010 17292
rect 2317 17289 2329 17292
rect 2363 17289 2375 17323
rect 2317 17283 2375 17289
rect 2777 17323 2835 17329
rect 2777 17289 2789 17323
rect 2823 17320 2835 17323
rect 3329 17323 3387 17329
rect 3329 17320 3341 17323
rect 2823 17292 3341 17320
rect 2823 17289 2835 17292
rect 2777 17283 2835 17289
rect 3329 17289 3341 17292
rect 3375 17289 3387 17323
rect 5442 17320 5448 17332
rect 3329 17283 3387 17289
rect 3620 17292 5448 17320
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 2498 17184 2504 17196
rect 1719 17156 2504 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 2682 17184 2688 17196
rect 2643 17156 2688 17184
rect 2682 17144 2688 17156
rect 2740 17144 2746 17196
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17116 3019 17119
rect 3620 17116 3648 17292
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 5626 17320 5632 17332
rect 5587 17292 5632 17320
rect 5626 17280 5632 17292
rect 5684 17280 5690 17332
rect 5721 17323 5779 17329
rect 5721 17289 5733 17323
rect 5767 17320 5779 17323
rect 5810 17320 5816 17332
rect 5767 17292 5816 17320
rect 5767 17289 5779 17292
rect 5721 17283 5779 17289
rect 5810 17280 5816 17292
rect 5868 17280 5874 17332
rect 6733 17323 6791 17329
rect 6733 17289 6745 17323
rect 6779 17320 6791 17323
rect 6822 17320 6828 17332
rect 6779 17292 6828 17320
rect 6779 17289 6791 17292
rect 6733 17283 6791 17289
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 7558 17320 7564 17332
rect 7519 17292 7564 17320
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 7926 17320 7932 17332
rect 7887 17292 7932 17320
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 9217 17323 9275 17329
rect 9217 17289 9229 17323
rect 9263 17320 9275 17323
rect 9674 17320 9680 17332
rect 9263 17292 9680 17320
rect 9263 17289 9275 17292
rect 9217 17283 9275 17289
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 10318 17320 10324 17332
rect 10279 17292 10324 17320
rect 10318 17280 10324 17292
rect 10376 17280 10382 17332
rect 10413 17323 10471 17329
rect 10413 17289 10425 17323
rect 10459 17320 10471 17323
rect 12158 17320 12164 17332
rect 10459 17292 12164 17320
rect 10459 17289 10471 17292
rect 10413 17283 10471 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 13173 17323 13231 17329
rect 13173 17289 13185 17323
rect 13219 17320 13231 17323
rect 13262 17320 13268 17332
rect 13219 17292 13268 17320
rect 13219 17289 13231 17292
rect 13173 17283 13231 17289
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 13814 17320 13820 17332
rect 13775 17292 13820 17320
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 14458 17320 14464 17332
rect 14419 17292 14464 17320
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 15562 17320 15568 17332
rect 15523 17292 15568 17320
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 17678 17320 17684 17332
rect 17639 17292 17684 17320
rect 17678 17280 17684 17292
rect 17736 17280 17742 17332
rect 17770 17280 17776 17332
rect 17828 17320 17834 17332
rect 19058 17320 19064 17332
rect 17828 17292 19064 17320
rect 17828 17280 17834 17292
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 19245 17323 19303 17329
rect 19245 17289 19257 17323
rect 19291 17320 19303 17323
rect 20622 17320 20628 17332
rect 19291 17292 20628 17320
rect 19291 17289 19303 17292
rect 19245 17283 19303 17289
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 4062 17212 4068 17264
rect 4120 17252 4126 17264
rect 8573 17255 8631 17261
rect 8573 17252 8585 17255
rect 4120 17224 8585 17252
rect 4120 17212 4126 17224
rect 8573 17221 8585 17224
rect 8619 17252 8631 17255
rect 9309 17255 9367 17261
rect 9309 17252 9321 17255
rect 8619 17224 9321 17252
rect 8619 17221 8631 17224
rect 8573 17215 8631 17221
rect 9309 17221 9321 17224
rect 9355 17252 9367 17255
rect 13630 17252 13636 17264
rect 9355 17224 13636 17252
rect 9355 17221 9367 17224
rect 9309 17215 9367 17221
rect 13630 17212 13636 17224
rect 13688 17212 13694 17264
rect 13725 17255 13783 17261
rect 13725 17221 13737 17255
rect 13771 17252 13783 17255
rect 14274 17252 14280 17264
rect 13771 17224 14280 17252
rect 13771 17221 13783 17224
rect 13725 17215 13783 17221
rect 14274 17212 14280 17224
rect 14332 17212 14338 17264
rect 14550 17212 14556 17264
rect 14608 17252 14614 17264
rect 14608 17224 15056 17252
rect 14608 17212 14614 17224
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 3007 17088 3648 17116
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 2041 16983 2099 16989
rect 2041 16949 2053 16983
rect 2087 16980 2099 16983
rect 3234 16980 3240 16992
rect 2087 16952 3240 16980
rect 2087 16949 2099 16952
rect 2041 16943 2099 16949
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 3712 16980 3740 17147
rect 3878 17144 3884 17196
rect 3936 17184 3942 17196
rect 6825 17187 6883 17193
rect 3936 17156 6500 17184
rect 3936 17144 3942 17156
rect 3789 17119 3847 17125
rect 3789 17085 3801 17119
rect 3835 17085 3847 17119
rect 3789 17079 3847 17085
rect 3973 17119 4031 17125
rect 3973 17085 3985 17119
rect 4019 17116 4031 17119
rect 4154 17116 4160 17128
rect 4019 17088 4160 17116
rect 4019 17085 4031 17088
rect 3973 17079 4031 17085
rect 3804 17048 3832 17079
rect 4154 17076 4160 17088
rect 4212 17076 4218 17128
rect 4982 17116 4988 17128
rect 4943 17088 4988 17116
rect 4982 17076 4988 17088
rect 5040 17076 5046 17128
rect 5905 17119 5963 17125
rect 5905 17085 5917 17119
rect 5951 17116 5963 17119
rect 5994 17116 6000 17128
rect 5951 17088 6000 17116
rect 5951 17085 5963 17088
rect 5905 17079 5963 17085
rect 5994 17076 6000 17088
rect 6052 17076 6058 17128
rect 6365 17051 6423 17057
rect 6365 17048 6377 17051
rect 3804 17020 6377 17048
rect 6365 17017 6377 17020
rect 6411 17017 6423 17051
rect 6472 17048 6500 17156
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 7006 17184 7012 17196
rect 6871 17156 7012 17184
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 7006 17144 7012 17156
rect 7064 17144 7070 17196
rect 7466 17144 7472 17196
rect 7524 17184 7530 17196
rect 9490 17184 9496 17196
rect 7524 17156 9496 17184
rect 7524 17144 7530 17156
rect 9490 17144 9496 17156
rect 9548 17144 9554 17196
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17184 12311 17187
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 12299 17156 12633 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 12621 17153 12633 17156
rect 12667 17184 12679 17187
rect 14458 17184 14464 17196
rect 12667 17156 14464 17184
rect 12667 17153 12679 17156
rect 12621 17147 12679 17153
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 14826 17184 14832 17196
rect 14787 17156 14832 17184
rect 14826 17144 14832 17156
rect 14884 17144 14890 17196
rect 6917 17119 6975 17125
rect 6917 17085 6929 17119
rect 6963 17116 6975 17119
rect 7190 17116 7196 17128
rect 6963 17088 7196 17116
rect 6963 17085 6975 17088
rect 6917 17079 6975 17085
rect 7190 17076 7196 17088
rect 7248 17076 7254 17128
rect 8018 17116 8024 17128
rect 7979 17088 8024 17116
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 8570 17116 8576 17128
rect 8251 17088 8576 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 8662 17076 8668 17128
rect 8720 17116 8726 17128
rect 9033 17119 9091 17125
rect 9033 17116 9045 17119
rect 8720 17088 9045 17116
rect 8720 17076 8726 17088
rect 9033 17085 9045 17088
rect 9079 17085 9091 17119
rect 10134 17116 10140 17128
rect 9033 17079 9091 17085
rect 9140 17088 9996 17116
rect 10095 17088 10140 17116
rect 9140 17048 9168 17088
rect 6472 17020 9168 17048
rect 9677 17051 9735 17057
rect 6365 17011 6423 17017
rect 9677 17017 9689 17051
rect 9723 17048 9735 17051
rect 9858 17048 9864 17060
rect 9723 17020 9864 17048
rect 9723 17017 9735 17020
rect 9677 17011 9735 17017
rect 9858 17008 9864 17020
rect 9916 17008 9922 17060
rect 9968 17048 9996 17088
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 11514 17116 11520 17128
rect 11475 17088 11520 17116
rect 11514 17076 11520 17088
rect 11572 17076 11578 17128
rect 13633 17119 13691 17125
rect 13633 17085 13645 17119
rect 13679 17085 13691 17119
rect 13633 17079 13691 17085
rect 11149 17051 11207 17057
rect 11149 17048 11161 17051
rect 9968 17020 11161 17048
rect 11149 17017 11161 17020
rect 11195 17048 11207 17051
rect 12526 17048 12532 17060
rect 11195 17020 12532 17048
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 13648 17048 13676 17079
rect 14366 17076 14372 17128
rect 14424 17116 14430 17128
rect 15028 17125 15056 17224
rect 15194 17212 15200 17264
rect 15252 17252 15258 17264
rect 15252 17224 20576 17252
rect 15252 17212 15258 17224
rect 15930 17184 15936 17196
rect 15891 17156 15936 17184
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17184 16083 17187
rect 17678 17184 17684 17196
rect 16071 17156 17684 17184
rect 16071 17153 16083 17156
rect 16025 17147 16083 17153
rect 17678 17144 17684 17156
rect 17736 17144 17742 17196
rect 18138 17144 18144 17196
rect 18196 17184 18202 17196
rect 18414 17184 18420 17196
rect 18196 17156 18420 17184
rect 18196 17144 18202 17156
rect 18414 17144 18420 17156
rect 18472 17144 18478 17196
rect 18874 17184 18880 17196
rect 18835 17156 18880 17184
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 19794 17144 19800 17196
rect 19852 17184 19858 17196
rect 20548 17193 20576 17224
rect 19889 17187 19947 17193
rect 19889 17184 19901 17187
rect 19852 17156 19901 17184
rect 19852 17144 19858 17156
rect 19889 17153 19901 17156
rect 19935 17153 19947 17187
rect 19889 17147 19947 17153
rect 20533 17187 20591 17193
rect 20533 17153 20545 17187
rect 20579 17153 20591 17187
rect 21082 17184 21088 17196
rect 21043 17156 21088 17184
rect 20533 17147 20591 17153
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 14424 17088 14933 17116
rect 14424 17076 14430 17088
rect 14921 17085 14933 17088
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17116 15071 17119
rect 16206 17116 16212 17128
rect 15059 17088 16077 17116
rect 16167 17088 16212 17116
rect 15059 17085 15071 17088
rect 15013 17079 15071 17085
rect 13814 17048 13820 17060
rect 13648 17020 13820 17048
rect 13814 17008 13820 17020
rect 13872 17008 13878 17060
rect 14936 17048 14964 17079
rect 15562 17048 15568 17060
rect 14936 17020 15568 17048
rect 15562 17008 15568 17020
rect 15620 17008 15626 17060
rect 16049 17048 16077 17088
rect 16206 17076 16212 17088
rect 16264 17076 16270 17128
rect 17497 17119 17555 17125
rect 17497 17085 17509 17119
rect 17543 17085 17555 17119
rect 17497 17079 17555 17085
rect 17589 17119 17647 17125
rect 17589 17085 17601 17119
rect 17635 17085 17647 17119
rect 18690 17116 18696 17128
rect 18651 17088 18696 17116
rect 17589 17079 17647 17085
rect 16669 17051 16727 17057
rect 16669 17048 16681 17051
rect 16049 17020 16681 17048
rect 16669 17017 16681 17020
rect 16715 17048 16727 17051
rect 17402 17048 17408 17060
rect 16715 17020 17408 17048
rect 16715 17017 16727 17020
rect 16669 17011 16727 17017
rect 17402 17008 17408 17020
rect 17460 17008 17466 17060
rect 4433 16983 4491 16989
rect 4433 16980 4445 16983
rect 3712 16952 4445 16980
rect 4433 16949 4445 16952
rect 4479 16980 4491 16983
rect 4522 16980 4528 16992
rect 4479 16952 4528 16980
rect 4479 16949 4491 16952
rect 4433 16943 4491 16949
rect 4522 16940 4528 16952
rect 4580 16940 4586 16992
rect 5258 16980 5264 16992
rect 5219 16952 5264 16980
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 5442 16940 5448 16992
rect 5500 16980 5506 16992
rect 8754 16980 8760 16992
rect 5500 16952 8760 16980
rect 5500 16940 5506 16952
rect 8754 16940 8760 16952
rect 8812 16940 8818 16992
rect 10778 16980 10784 16992
rect 10739 16952 10784 16980
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 14185 16983 14243 16989
rect 14185 16949 14197 16983
rect 14231 16980 14243 16983
rect 15746 16980 15752 16992
rect 14231 16952 15752 16980
rect 14231 16949 14243 16952
rect 14185 16943 14243 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 17512 16980 17540 17079
rect 17604 17048 17632 17079
rect 18690 17076 18696 17088
rect 18748 17076 18754 17128
rect 18785 17119 18843 17125
rect 18785 17085 18797 17119
rect 18831 17116 18843 17119
rect 19610 17116 19616 17128
rect 18831 17088 19616 17116
rect 18831 17085 18843 17088
rect 18785 17079 18843 17085
rect 19610 17076 19616 17088
rect 19668 17076 19674 17128
rect 19702 17076 19708 17128
rect 19760 17116 19766 17128
rect 19981 17119 20039 17125
rect 19981 17116 19993 17119
rect 19760 17088 19993 17116
rect 19760 17076 19766 17088
rect 19981 17085 19993 17088
rect 20027 17085 20039 17119
rect 19981 17079 20039 17085
rect 20073 17119 20131 17125
rect 20073 17085 20085 17119
rect 20119 17085 20131 17119
rect 20073 17079 20131 17085
rect 19521 17051 19579 17057
rect 19521 17048 19533 17051
rect 17604 17020 19533 17048
rect 19521 17017 19533 17020
rect 19567 17017 19579 17051
rect 19521 17011 19579 17017
rect 17954 16980 17960 16992
rect 17512 16952 17960 16980
rect 17954 16940 17960 16952
rect 18012 16940 18018 16992
rect 18049 16983 18107 16989
rect 18049 16949 18061 16983
rect 18095 16980 18107 16983
rect 18506 16980 18512 16992
rect 18095 16952 18512 16980
rect 18095 16949 18107 16952
rect 18049 16943 18107 16949
rect 18506 16940 18512 16952
rect 18564 16940 18570 16992
rect 18598 16940 18604 16992
rect 18656 16980 18662 16992
rect 20088 16980 20116 17079
rect 20714 16980 20720 16992
rect 18656 16952 20116 16980
rect 20675 16952 20720 16980
rect 18656 16940 18662 16952
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 21266 16980 21272 16992
rect 21227 16952 21272 16980
rect 21266 16940 21272 16952
rect 21324 16940 21330 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 4525 16779 4583 16785
rect 4525 16745 4537 16779
rect 4571 16776 4583 16779
rect 5074 16776 5080 16788
rect 4571 16748 5080 16776
rect 4571 16745 4583 16748
rect 4525 16739 4583 16745
rect 1578 16668 1584 16720
rect 1636 16708 1642 16720
rect 4540 16708 4568 16739
rect 5074 16736 5080 16748
rect 5132 16736 5138 16788
rect 6181 16779 6239 16785
rect 6181 16745 6193 16779
rect 6227 16776 6239 16779
rect 7190 16776 7196 16788
rect 6227 16748 7196 16776
rect 6227 16745 6239 16748
rect 6181 16739 6239 16745
rect 7190 16736 7196 16748
rect 7248 16776 7254 16788
rect 10042 16776 10048 16788
rect 7248 16748 10048 16776
rect 7248 16736 7254 16748
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 11146 16776 11152 16788
rect 10612 16748 11152 16776
rect 6822 16708 6828 16720
rect 1636 16680 4568 16708
rect 4816 16680 6828 16708
rect 1636 16668 1642 16680
rect 4154 16640 4160 16652
rect 4067 16612 4160 16640
rect 4154 16600 4160 16612
rect 4212 16640 4218 16652
rect 4816 16640 4844 16680
rect 6822 16668 6828 16680
rect 6880 16668 6886 16720
rect 6917 16711 6975 16717
rect 6917 16677 6929 16711
rect 6963 16708 6975 16711
rect 7098 16708 7104 16720
rect 6963 16680 7104 16708
rect 6963 16677 6975 16680
rect 6917 16671 6975 16677
rect 7098 16668 7104 16680
rect 7156 16708 7162 16720
rect 7926 16708 7932 16720
rect 7156 16680 7932 16708
rect 7156 16668 7162 16680
rect 7926 16668 7932 16680
rect 7984 16668 7990 16720
rect 9950 16708 9956 16720
rect 9911 16680 9956 16708
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 10612 16652 10640 16748
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 12158 16736 12164 16788
rect 12216 16776 12222 16788
rect 12342 16776 12348 16788
rect 12216 16748 12348 16776
rect 12216 16736 12222 16748
rect 12342 16736 12348 16748
rect 12400 16776 12406 16788
rect 15286 16776 15292 16788
rect 12400 16748 15292 16776
rect 12400 16736 12406 16748
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 16022 16736 16028 16788
rect 16080 16776 16086 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 16080 16748 16405 16776
rect 16080 16736 16086 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 16393 16739 16451 16745
rect 17221 16779 17279 16785
rect 17221 16745 17233 16779
rect 17267 16776 17279 16779
rect 17310 16776 17316 16788
rect 17267 16748 17316 16776
rect 17267 16745 17279 16748
rect 17221 16739 17279 16745
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 17770 16776 17776 16788
rect 17512 16748 17776 16776
rect 17512 16720 17540 16748
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 18233 16779 18291 16785
rect 18233 16745 18245 16779
rect 18279 16776 18291 16779
rect 18874 16776 18880 16788
rect 18279 16748 18880 16776
rect 18279 16745 18291 16748
rect 18233 16739 18291 16745
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 19610 16776 19616 16788
rect 19571 16748 19616 16776
rect 19610 16736 19616 16748
rect 19668 16736 19674 16788
rect 10686 16668 10692 16720
rect 10744 16708 10750 16720
rect 10744 16680 12434 16708
rect 10744 16668 10750 16680
rect 4212 16612 4844 16640
rect 4893 16643 4951 16649
rect 4212 16600 4218 16612
rect 4893 16609 4905 16643
rect 4939 16640 4951 16643
rect 7837 16643 7895 16649
rect 7837 16640 7849 16643
rect 4939 16612 7849 16640
rect 4939 16609 4951 16612
rect 4893 16603 4951 16609
rect 7837 16609 7849 16612
rect 7883 16640 7895 16643
rect 9214 16640 9220 16652
rect 7883 16612 9220 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 9490 16640 9496 16652
rect 9451 16612 9496 16640
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 10318 16640 10324 16652
rect 10279 16612 10324 16640
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 10594 16600 10600 16652
rect 10652 16640 10658 16652
rect 10781 16643 10839 16649
rect 10781 16640 10793 16643
rect 10652 16612 10793 16640
rect 10652 16600 10658 16612
rect 10781 16609 10793 16612
rect 10827 16609 10839 16643
rect 11054 16640 11060 16652
rect 11015 16612 11060 16640
rect 10781 16603 10839 16609
rect 11054 16600 11060 16612
rect 11112 16600 11118 16652
rect 12406 16640 12434 16680
rect 13538 16668 13544 16720
rect 13596 16708 13602 16720
rect 17494 16708 17500 16720
rect 13596 16680 17500 16708
rect 13596 16668 13602 16680
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 17604 16680 18736 16708
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 12406 16612 12633 16640
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 13078 16640 13084 16652
rect 13039 16612 13084 16640
rect 12621 16603 12679 16609
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 13630 16640 13636 16652
rect 13591 16612 13636 16640
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 14553 16643 14611 16649
rect 14553 16609 14565 16643
rect 14599 16640 14611 16643
rect 14826 16640 14832 16652
rect 14599 16612 14832 16640
rect 14599 16609 14611 16612
rect 14553 16603 14611 16609
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 15105 16643 15163 16649
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 15470 16640 15476 16652
rect 15151 16612 15476 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 15470 16600 15476 16612
rect 15528 16640 15534 16652
rect 16025 16643 16083 16649
rect 16025 16640 16037 16643
rect 15528 16612 16037 16640
rect 15528 16600 15534 16612
rect 16025 16609 16037 16612
rect 16071 16640 16083 16643
rect 16853 16643 16911 16649
rect 16071 16612 16804 16640
rect 16071 16609 16083 16612
rect 16025 16603 16083 16609
rect 1670 16572 1676 16584
rect 1631 16544 1676 16572
rect 1670 16532 1676 16544
rect 1728 16532 1734 16584
rect 2317 16575 2375 16581
rect 2317 16541 2329 16575
rect 2363 16541 2375 16575
rect 2317 16535 2375 16541
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 3234 16572 3240 16584
rect 3007 16544 3240 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 106 16464 112 16516
rect 164 16504 170 16516
rect 1394 16504 1400 16516
rect 164 16476 1400 16504
rect 164 16464 170 16476
rect 1394 16464 1400 16476
rect 1452 16464 1458 16516
rect 2332 16504 2360 16535
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 3326 16532 3332 16584
rect 3384 16572 3390 16584
rect 3421 16575 3479 16581
rect 3421 16572 3433 16575
rect 3384 16544 3433 16572
rect 3384 16532 3390 16544
rect 3421 16541 3433 16544
rect 3467 16541 3479 16575
rect 3421 16535 3479 16541
rect 4982 16532 4988 16584
rect 5040 16572 5046 16584
rect 5169 16575 5227 16581
rect 5169 16572 5181 16575
rect 5040 16544 5181 16572
rect 5040 16532 5046 16544
rect 5169 16541 5181 16544
rect 5215 16541 5227 16575
rect 5169 16535 5227 16541
rect 7653 16575 7711 16581
rect 7653 16541 7665 16575
rect 7699 16572 7711 16575
rect 7926 16572 7932 16584
rect 7699 16544 7932 16572
rect 7699 16541 7711 16544
rect 7653 16535 7711 16541
rect 7926 16532 7932 16544
rect 7984 16532 7990 16584
rect 9306 16572 9312 16584
rect 9267 16544 9312 16572
rect 9306 16532 9312 16544
rect 9364 16532 9370 16584
rect 11885 16575 11943 16581
rect 11885 16541 11897 16575
rect 11931 16572 11943 16575
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 11931 16544 12265 16572
rect 11931 16541 11943 16544
rect 11885 16535 11943 16541
rect 12253 16541 12265 16544
rect 12299 16572 12311 16575
rect 13170 16572 13176 16584
rect 12299 16544 13176 16572
rect 12299 16541 12311 16544
rect 12253 16535 12311 16541
rect 13170 16532 13176 16544
rect 13228 16572 13234 16584
rect 13722 16572 13728 16584
rect 13228 16544 13728 16572
rect 13228 16532 13234 16544
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 5258 16504 5264 16516
rect 2332 16476 5264 16504
rect 5258 16464 5264 16476
rect 5316 16464 5322 16516
rect 6549 16507 6607 16513
rect 6549 16473 6561 16507
rect 6595 16504 6607 16507
rect 7561 16507 7619 16513
rect 7561 16504 7573 16507
rect 6595 16476 7573 16504
rect 6595 16473 6607 16476
rect 6549 16467 6607 16473
rect 7561 16473 7573 16476
rect 7607 16504 7619 16507
rect 7742 16504 7748 16516
rect 7607 16476 7748 16504
rect 7607 16473 7619 16476
rect 7561 16467 7619 16473
rect 7742 16464 7748 16476
rect 7800 16504 7806 16516
rect 12618 16504 12624 16516
rect 7800 16476 12624 16504
rect 7800 16464 7806 16476
rect 12618 16464 12624 16476
rect 12676 16464 12682 16516
rect 14918 16464 14924 16516
rect 14976 16504 14982 16516
rect 15289 16507 15347 16513
rect 15289 16504 15301 16507
rect 14976 16476 15301 16504
rect 14976 16464 14982 16476
rect 15289 16473 15301 16476
rect 15335 16473 15347 16507
rect 16776 16504 16804 16612
rect 16853 16609 16865 16643
rect 16899 16640 16911 16643
rect 17218 16640 17224 16652
rect 16899 16612 17224 16640
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 17604 16649 17632 16680
rect 17589 16643 17647 16649
rect 17589 16609 17601 16643
rect 17635 16609 17647 16643
rect 17770 16640 17776 16652
rect 17731 16612 17776 16640
rect 17589 16603 17647 16609
rect 17770 16600 17776 16612
rect 17828 16600 17834 16652
rect 18708 16640 18736 16680
rect 18782 16640 18788 16652
rect 18708 16612 18788 16640
rect 18782 16600 18788 16612
rect 18840 16640 18846 16652
rect 20165 16643 20223 16649
rect 20165 16640 20177 16643
rect 18840 16612 20177 16640
rect 18840 16600 18846 16612
rect 20165 16609 20177 16612
rect 20211 16609 20223 16643
rect 20165 16603 20223 16609
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 21174 16640 21180 16652
rect 20956 16612 21036 16640
rect 21135 16612 21180 16640
rect 20956 16600 20962 16612
rect 18506 16572 18512 16584
rect 18467 16544 18512 16572
rect 18506 16532 18512 16544
rect 18564 16532 18570 16584
rect 20806 16572 20812 16584
rect 18708 16544 20812 16572
rect 17770 16504 17776 16516
rect 16776 16476 17776 16504
rect 15289 16467 15347 16473
rect 17770 16464 17776 16476
rect 17828 16464 17834 16516
rect 17865 16507 17923 16513
rect 17865 16473 17877 16507
rect 17911 16473 17923 16507
rect 17865 16467 17923 16473
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 2130 16436 2136 16448
rect 2091 16408 2136 16436
rect 2130 16396 2136 16408
rect 2188 16396 2194 16448
rect 2590 16396 2596 16448
rect 2648 16436 2654 16448
rect 2777 16439 2835 16445
rect 2777 16436 2789 16439
rect 2648 16408 2789 16436
rect 2648 16396 2654 16408
rect 2777 16405 2789 16408
rect 2823 16405 2835 16439
rect 2777 16399 2835 16405
rect 2958 16396 2964 16448
rect 3016 16436 3022 16448
rect 3237 16439 3295 16445
rect 3237 16436 3249 16439
rect 3016 16408 3249 16436
rect 3016 16396 3022 16408
rect 3237 16405 3249 16408
rect 3283 16405 3295 16439
rect 5074 16436 5080 16448
rect 5035 16408 5080 16436
rect 3237 16399 3295 16405
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 5534 16436 5540 16448
rect 5495 16408 5540 16436
rect 5534 16396 5540 16408
rect 5592 16396 5598 16448
rect 7190 16436 7196 16448
rect 7151 16408 7196 16436
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 8202 16436 8208 16448
rect 8163 16408 8208 16436
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 8386 16396 8392 16448
rect 8444 16436 8450 16448
rect 8941 16439 8999 16445
rect 8941 16436 8953 16439
rect 8444 16408 8953 16436
rect 8444 16396 8450 16408
rect 8941 16405 8953 16408
rect 8987 16405 8999 16439
rect 8941 16399 8999 16405
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 9456 16408 9501 16436
rect 9456 16396 9462 16408
rect 14642 16396 14648 16448
rect 14700 16436 14706 16448
rect 15197 16439 15255 16445
rect 15197 16436 15209 16439
rect 14700 16408 15209 16436
rect 14700 16396 14706 16408
rect 15197 16405 15209 16408
rect 15243 16405 15255 16439
rect 15654 16436 15660 16448
rect 15615 16408 15660 16436
rect 15197 16399 15255 16405
rect 15654 16396 15660 16408
rect 15712 16396 15718 16448
rect 17880 16436 17908 16467
rect 18506 16436 18512 16448
rect 17880 16408 18512 16436
rect 18506 16396 18512 16408
rect 18564 16396 18570 16448
rect 18708 16445 18736 16544
rect 20806 16532 20812 16544
rect 20864 16532 20870 16584
rect 21008 16572 21036 16612
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 21008 16544 21097 16572
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 18693 16439 18751 16445
rect 18693 16405 18705 16439
rect 18739 16405 18751 16439
rect 18693 16399 18751 16405
rect 19058 16396 19064 16448
rect 19116 16436 19122 16448
rect 19245 16439 19303 16445
rect 19245 16436 19257 16439
rect 19116 16408 19257 16436
rect 19116 16396 19122 16408
rect 19245 16405 19257 16408
rect 19291 16405 19303 16439
rect 19245 16399 19303 16405
rect 19610 16396 19616 16448
rect 19668 16436 19674 16448
rect 19981 16439 20039 16445
rect 19981 16436 19993 16439
rect 19668 16408 19993 16436
rect 19668 16396 19674 16408
rect 19981 16405 19993 16408
rect 20027 16405 20039 16439
rect 19981 16399 20039 16405
rect 20073 16439 20131 16445
rect 20073 16405 20085 16439
rect 20119 16436 20131 16439
rect 20162 16436 20168 16448
rect 20119 16408 20168 16436
rect 20119 16405 20131 16408
rect 20073 16399 20131 16405
rect 20162 16396 20168 16408
rect 20220 16396 20226 16448
rect 20622 16436 20628 16448
rect 20583 16408 20628 16436
rect 20622 16396 20628 16408
rect 20680 16396 20686 16448
rect 20993 16439 21051 16445
rect 20993 16405 21005 16439
rect 21039 16436 21051 16439
rect 21082 16436 21088 16448
rect 21039 16408 21088 16436
rect 21039 16405 21051 16408
rect 20993 16399 21051 16405
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 2498 16232 2504 16244
rect 2459 16204 2504 16232
rect 2498 16192 2504 16204
rect 2556 16192 2562 16244
rect 3326 16232 3332 16244
rect 3287 16204 3332 16232
rect 3326 16192 3332 16204
rect 3384 16192 3390 16244
rect 3620 16204 4016 16232
rect 3620 16164 3648 16204
rect 2700 16136 3648 16164
rect 3697 16167 3755 16173
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 2225 16099 2283 16105
rect 2225 16065 2237 16099
rect 2271 16096 2283 16099
rect 2590 16096 2596 16108
rect 2271 16068 2596 16096
rect 2271 16065 2283 16068
rect 2225 16059 2283 16065
rect 1688 16028 1716 16059
rect 2590 16056 2596 16068
rect 2648 16056 2654 16108
rect 2700 16105 2728 16136
rect 3697 16133 3709 16167
rect 3743 16164 3755 16167
rect 3878 16164 3884 16176
rect 3743 16136 3884 16164
rect 3743 16133 3755 16136
rect 3697 16127 3755 16133
rect 3878 16124 3884 16136
rect 3936 16124 3942 16176
rect 3988 16164 4016 16204
rect 5350 16192 5356 16244
rect 5408 16232 5414 16244
rect 5813 16235 5871 16241
rect 5813 16232 5825 16235
rect 5408 16204 5825 16232
rect 5408 16192 5414 16204
rect 5813 16201 5825 16204
rect 5859 16201 5871 16235
rect 5813 16195 5871 16201
rect 7653 16235 7711 16241
rect 7653 16201 7665 16235
rect 7699 16232 7711 16235
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 7699 16204 8217 16232
rect 7699 16201 7711 16204
rect 7653 16195 7711 16201
rect 8205 16201 8217 16204
rect 8251 16201 8263 16235
rect 8205 16195 8263 16201
rect 8665 16235 8723 16241
rect 8665 16201 8677 16235
rect 8711 16232 8723 16235
rect 9398 16232 9404 16244
rect 8711 16204 9404 16232
rect 8711 16201 8723 16204
rect 8665 16195 8723 16201
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 10870 16192 10876 16244
rect 10928 16232 10934 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 10928 16204 11529 16232
rect 10928 16192 10934 16204
rect 11517 16201 11529 16204
rect 11563 16232 11575 16235
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 11563 16204 11897 16232
rect 11563 16201 11575 16204
rect 11517 16195 11575 16201
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 12618 16232 12624 16244
rect 12579 16204 12624 16232
rect 11885 16195 11943 16201
rect 5445 16167 5503 16173
rect 5445 16164 5457 16167
rect 3988 16136 5457 16164
rect 5445 16133 5457 16136
rect 5491 16164 5503 16167
rect 7006 16164 7012 16176
rect 5491 16136 7012 16164
rect 5491 16133 5503 16136
rect 5445 16127 5503 16133
rect 7006 16124 7012 16136
rect 7064 16164 7070 16176
rect 7193 16167 7251 16173
rect 7193 16164 7205 16167
rect 7064 16136 7205 16164
rect 7064 16124 7070 16136
rect 7193 16133 7205 16136
rect 7239 16164 7251 16167
rect 8110 16164 8116 16176
rect 7239 16136 8116 16164
rect 7239 16133 7251 16136
rect 7193 16127 7251 16133
rect 8110 16124 8116 16136
rect 8168 16124 8174 16176
rect 11422 16164 11428 16176
rect 8220 16136 11428 16164
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16065 2743 16099
rect 2685 16059 2743 16065
rect 3789 16099 3847 16105
rect 3789 16065 3801 16099
rect 3835 16096 3847 16099
rect 4062 16096 4068 16108
rect 3835 16068 4068 16096
rect 3835 16065 3847 16068
rect 3789 16059 3847 16065
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 6748 16068 7297 16096
rect 6748 16040 6776 16068
rect 7285 16065 7297 16068
rect 7331 16096 7343 16099
rect 8220 16096 8248 16136
rect 11422 16124 11428 16136
rect 11480 16124 11486 16176
rect 11900 16164 11928 16195
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 15470 16232 15476 16244
rect 15383 16204 15476 16232
rect 15470 16192 15476 16204
rect 15528 16232 15534 16244
rect 15930 16232 15936 16244
rect 15528 16204 15936 16232
rect 15528 16192 15534 16204
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 17221 16235 17279 16241
rect 17221 16201 17233 16235
rect 17267 16232 17279 16235
rect 18046 16232 18052 16244
rect 17267 16204 18052 16232
rect 17267 16201 17279 16204
rect 17221 16195 17279 16201
rect 18046 16192 18052 16204
rect 18104 16192 18110 16244
rect 18969 16235 19027 16241
rect 18969 16201 18981 16235
rect 19015 16201 19027 16235
rect 18969 16195 19027 16201
rect 12989 16167 13047 16173
rect 12989 16164 13001 16167
rect 11900 16136 13001 16164
rect 12989 16133 13001 16136
rect 13035 16164 13047 16167
rect 13170 16164 13176 16176
rect 13035 16136 13176 16164
rect 13035 16133 13047 16136
rect 12989 16127 13047 16133
rect 13170 16124 13176 16136
rect 13228 16124 13234 16176
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 15841 16167 15899 16173
rect 15841 16164 15853 16167
rect 15344 16136 15853 16164
rect 15344 16124 15350 16136
rect 15841 16133 15853 16136
rect 15887 16164 15899 16167
rect 16209 16167 16267 16173
rect 16209 16164 16221 16167
rect 15887 16136 16221 16164
rect 15887 16133 15899 16136
rect 15841 16127 15899 16133
rect 16209 16133 16221 16136
rect 16255 16133 16267 16167
rect 17494 16164 17500 16176
rect 17455 16136 17500 16164
rect 16209 16127 16267 16133
rect 17494 16124 17500 16136
rect 17552 16124 17558 16176
rect 7331 16068 8248 16096
rect 8297 16099 8355 16105
rect 7331 16065 7343 16068
rect 7285 16059 7343 16065
rect 8297 16065 8309 16099
rect 8343 16096 8355 16099
rect 8343 16068 8432 16096
rect 8343 16065 8355 16068
rect 8297 16059 8355 16065
rect 2498 16028 2504 16040
rect 1688 16000 2504 16028
rect 2498 15988 2504 16000
rect 2556 15988 2562 16040
rect 3694 15988 3700 16040
rect 3752 16028 3758 16040
rect 3881 16031 3939 16037
rect 3881 16028 3893 16031
rect 3752 16000 3893 16028
rect 3752 15988 3758 16000
rect 3881 15997 3893 16000
rect 3927 15997 3939 16031
rect 3881 15991 3939 15997
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 16028 6699 16031
rect 6730 16028 6736 16040
rect 6687 16000 6736 16028
rect 6687 15997 6699 16000
rect 6641 15991 6699 15997
rect 6730 15988 6736 16000
rect 6788 15988 6794 16040
rect 7098 16028 7104 16040
rect 7059 16000 7104 16028
rect 7098 15988 7104 16000
rect 7156 15988 7162 16040
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 16028 8171 16031
rect 8202 16028 8208 16040
rect 8159 16000 8208 16028
rect 8159 15997 8171 16000
rect 8113 15991 8171 15997
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 2038 15960 2044 15972
rect 1999 15932 2044 15960
rect 2038 15920 2044 15932
rect 2096 15920 2102 15972
rect 2774 15920 2780 15972
rect 2832 15960 2838 15972
rect 4985 15963 5043 15969
rect 4985 15960 4997 15963
rect 2832 15932 4997 15960
rect 2832 15920 2838 15932
rect 4985 15929 4997 15932
rect 5031 15960 5043 15963
rect 7558 15960 7564 15972
rect 5031 15932 7564 15960
rect 5031 15929 5043 15932
rect 4985 15923 5043 15929
rect 7558 15920 7564 15932
rect 7616 15920 7622 15972
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 2866 15852 2872 15904
rect 2924 15892 2930 15904
rect 2961 15895 3019 15901
rect 2961 15892 2973 15895
rect 2924 15864 2973 15892
rect 2924 15852 2930 15864
rect 2961 15861 2973 15864
rect 3007 15861 3019 15895
rect 2961 15855 3019 15861
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15892 4767 15895
rect 4798 15892 4804 15904
rect 4755 15864 4804 15892
rect 4755 15861 4767 15864
rect 4709 15855 4767 15861
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 7926 15892 7932 15904
rect 5224 15864 7932 15892
rect 5224 15852 5230 15864
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 8202 15852 8208 15904
rect 8260 15892 8266 15904
rect 8404 15892 8432 16068
rect 10042 16056 10048 16108
rect 10100 16096 10106 16108
rect 10870 16096 10876 16108
rect 10100 16068 10876 16096
rect 10100 16056 10106 16068
rect 10870 16056 10876 16068
rect 10928 16056 10934 16108
rect 14918 16096 14924 16108
rect 13924 16068 14924 16096
rect 13924 16028 13952 16068
rect 14918 16056 14924 16068
rect 14976 16056 14982 16108
rect 15562 16056 15568 16108
rect 15620 16096 15626 16108
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 15620 16068 16681 16096
rect 15620 16056 15626 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 18785 16099 18843 16105
rect 18785 16096 18797 16099
rect 16669 16059 16727 16065
rect 18432 16068 18797 16096
rect 8956 16000 13952 16028
rect 14277 16031 14335 16037
rect 8956 15901 8984 16000
rect 14277 15997 14289 16031
rect 14323 16028 14335 16031
rect 14550 16028 14556 16040
rect 14323 16000 14556 16028
rect 14323 15997 14335 16000
rect 14277 15991 14335 15997
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 9769 15963 9827 15969
rect 9769 15929 9781 15963
rect 9815 15960 9827 15963
rect 10318 15960 10324 15972
rect 9815 15932 10324 15960
rect 9815 15929 9827 15932
rect 9769 15923 9827 15929
rect 10318 15920 10324 15932
rect 10376 15920 10382 15972
rect 10505 15963 10563 15969
rect 10505 15929 10517 15963
rect 10551 15960 10563 15963
rect 10962 15960 10968 15972
rect 10551 15932 10968 15960
rect 10551 15929 10563 15932
rect 10505 15923 10563 15929
rect 10962 15920 10968 15932
rect 11020 15920 11026 15972
rect 13909 15963 13967 15969
rect 13909 15929 13921 15963
rect 13955 15960 13967 15963
rect 16942 15960 16948 15972
rect 13955 15932 16948 15960
rect 13955 15929 13967 15932
rect 13909 15923 13967 15929
rect 16942 15920 16948 15932
rect 17000 15920 17006 15972
rect 18138 15960 18144 15972
rect 18099 15932 18144 15960
rect 18138 15920 18144 15932
rect 18196 15960 18202 15972
rect 18432 15969 18460 16068
rect 18785 16065 18797 16068
rect 18831 16096 18843 16099
rect 18874 16096 18880 16108
rect 18831 16068 18880 16096
rect 18831 16065 18843 16068
rect 18785 16059 18843 16065
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 18984 16096 19012 16195
rect 20622 16192 20628 16244
rect 20680 16232 20686 16244
rect 20717 16235 20775 16241
rect 20717 16232 20729 16235
rect 20680 16204 20729 16232
rect 20680 16192 20686 16204
rect 20717 16201 20729 16204
rect 20763 16201 20775 16235
rect 20717 16195 20775 16201
rect 19429 16167 19487 16173
rect 19429 16133 19441 16167
rect 19475 16164 19487 16167
rect 19475 16136 20668 16164
rect 19475 16133 19487 16136
rect 19429 16127 19487 16133
rect 20640 16105 20668 16136
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 18984 16068 19717 16096
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19705 16059 19763 16065
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 19518 15988 19524 16040
rect 19576 16028 19582 16040
rect 20809 16031 20867 16037
rect 20809 16028 20821 16031
rect 19576 16000 20821 16028
rect 19576 15988 19582 16000
rect 20809 15997 20821 16000
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 18417 15963 18475 15969
rect 18417 15960 18429 15963
rect 18196 15932 18429 15960
rect 18196 15920 18202 15932
rect 18417 15929 18429 15932
rect 18463 15929 18475 15963
rect 18417 15923 18475 15929
rect 18506 15920 18512 15972
rect 18564 15960 18570 15972
rect 20257 15963 20315 15969
rect 20257 15960 20269 15963
rect 18564 15932 20269 15960
rect 18564 15920 18570 15932
rect 20257 15929 20269 15932
rect 20303 15929 20315 15963
rect 20257 15923 20315 15929
rect 8941 15895 8999 15901
rect 8941 15892 8953 15895
rect 8260 15864 8953 15892
rect 8260 15852 8266 15864
rect 8941 15861 8953 15864
rect 8987 15861 8999 15895
rect 9398 15892 9404 15904
rect 9359 15864 9404 15892
rect 8941 15855 8999 15861
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 10042 15892 10048 15904
rect 10003 15864 10048 15892
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 10870 15892 10876 15904
rect 10831 15864 10876 15892
rect 10870 15852 10876 15864
rect 10928 15852 10934 15904
rect 12342 15892 12348 15904
rect 12303 15864 12348 15892
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 13354 15892 13360 15904
rect 13315 15864 13360 15892
rect 13354 15852 13360 15864
rect 13412 15852 13418 15904
rect 14642 15892 14648 15904
rect 14603 15864 14648 15892
rect 14642 15852 14648 15864
rect 14700 15852 14706 15904
rect 19886 15892 19892 15904
rect 19847 15864 19892 15892
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 21266 15892 21272 15904
rect 21227 15864 21272 15892
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 2222 15688 2228 15700
rect 2183 15660 2228 15688
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 2498 15648 2504 15700
rect 2556 15688 2562 15700
rect 2685 15691 2743 15697
rect 2685 15688 2697 15691
rect 2556 15660 2697 15688
rect 2556 15648 2562 15660
rect 2685 15657 2697 15660
rect 2731 15657 2743 15691
rect 2685 15651 2743 15657
rect 5902 15648 5908 15700
rect 5960 15688 5966 15700
rect 6089 15691 6147 15697
rect 6089 15688 6101 15691
rect 5960 15660 6101 15688
rect 5960 15648 5966 15660
rect 6089 15657 6101 15660
rect 6135 15657 6147 15691
rect 6089 15651 6147 15657
rect 8662 15648 8668 15700
rect 8720 15688 8726 15700
rect 9309 15691 9367 15697
rect 9309 15688 9321 15691
rect 8720 15660 9321 15688
rect 8720 15648 8726 15660
rect 9309 15657 9321 15660
rect 9355 15657 9367 15691
rect 11146 15688 11152 15700
rect 9309 15651 9367 15657
rect 9784 15660 11152 15688
rect 1394 15580 1400 15632
rect 1452 15620 1458 15632
rect 8202 15620 8208 15632
rect 1452 15592 8208 15620
rect 1452 15580 1458 15592
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 8294 15580 8300 15632
rect 8352 15620 8358 15632
rect 9784 15620 9812 15660
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 11330 15688 11336 15700
rect 11291 15660 11336 15688
rect 11330 15648 11336 15660
rect 11388 15648 11394 15700
rect 11698 15688 11704 15700
rect 11659 15660 11704 15688
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 17494 15688 17500 15700
rect 15948 15660 17500 15688
rect 15948 15620 15976 15660
rect 17494 15648 17500 15660
rect 17552 15648 17558 15700
rect 17678 15688 17684 15700
rect 17639 15660 17684 15688
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 8352 15592 9812 15620
rect 11348 15592 15976 15620
rect 8352 15580 8358 15592
rect 3881 15555 3939 15561
rect 3881 15521 3893 15555
rect 3927 15552 3939 15555
rect 4798 15552 4804 15564
rect 3927 15524 4804 15552
rect 3927 15521 3939 15524
rect 3881 15515 3939 15521
rect 4798 15512 4804 15524
rect 4856 15512 4862 15564
rect 5074 15512 5080 15564
rect 5132 15552 5138 15564
rect 5350 15552 5356 15564
rect 5132 15524 5356 15552
rect 5132 15512 5138 15524
rect 5350 15512 5356 15524
rect 5408 15552 5414 15564
rect 5537 15555 5595 15561
rect 5537 15552 5549 15555
rect 5408 15524 5549 15552
rect 5408 15512 5414 15524
rect 5537 15521 5549 15524
rect 5583 15521 5595 15555
rect 5537 15515 5595 15521
rect 6362 15512 6368 15564
rect 6420 15552 6426 15564
rect 6733 15555 6791 15561
rect 6733 15552 6745 15555
rect 6420 15524 6745 15552
rect 6420 15512 6426 15524
rect 6733 15521 6745 15524
rect 6779 15552 6791 15555
rect 7006 15552 7012 15564
rect 6779 15524 7012 15552
rect 6779 15521 6791 15524
rect 6733 15515 6791 15521
rect 7006 15512 7012 15524
rect 7064 15512 7070 15564
rect 7558 15552 7564 15564
rect 7519 15524 7564 15552
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 7745 15555 7803 15561
rect 7745 15521 7757 15555
rect 7791 15552 7803 15555
rect 8110 15552 8116 15564
rect 7791 15524 8116 15552
rect 7791 15521 7803 15524
rect 7745 15515 7803 15521
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 8389 15555 8447 15561
rect 8389 15552 8401 15555
rect 8220 15524 8401 15552
rect 842 15444 848 15496
rect 900 15484 906 15496
rect 1486 15484 1492 15496
rect 900 15456 1492 15484
rect 900 15444 906 15456
rect 1486 15444 1492 15456
rect 1544 15444 1550 15496
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15444 1734 15496
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15484 2467 15487
rect 2774 15484 2780 15496
rect 2455 15456 2780 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 2774 15444 2780 15456
rect 2832 15444 2838 15496
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15484 2927 15487
rect 2915 15456 3280 15484
rect 2915 15453 2927 15456
rect 2869 15447 2927 15453
rect 3252 15360 3280 15456
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 4157 15487 4215 15493
rect 4157 15484 4169 15487
rect 4028 15456 4169 15484
rect 4028 15444 4034 15456
rect 4157 15453 4169 15456
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15484 6515 15487
rect 6546 15484 6552 15496
rect 6503 15456 6552 15484
rect 6503 15453 6515 15456
rect 6457 15447 6515 15453
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 8220 15484 8248 15524
rect 8389 15521 8401 15524
rect 8435 15552 8447 15555
rect 8754 15552 8760 15564
rect 8435 15524 8760 15552
rect 8435 15521 8447 15524
rect 8389 15515 8447 15521
rect 8754 15512 8760 15524
rect 8812 15512 8818 15564
rect 7515 15456 8248 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 8294 15444 8300 15496
rect 8352 15484 8358 15496
rect 8478 15484 8484 15496
rect 8352 15456 8484 15484
rect 8352 15444 8358 15456
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 9732 15456 10701 15484
rect 9732 15444 9738 15456
rect 10689 15453 10701 15456
rect 10735 15484 10747 15487
rect 10965 15487 11023 15493
rect 10965 15484 10977 15487
rect 10735 15456 10977 15484
rect 10735 15453 10747 15456
rect 10689 15447 10747 15453
rect 10965 15453 10977 15456
rect 11011 15484 11023 15487
rect 11238 15484 11244 15496
rect 11011 15456 11244 15484
rect 11011 15453 11023 15456
rect 10965 15447 11023 15453
rect 11238 15444 11244 15456
rect 11296 15444 11302 15496
rect 3326 15376 3332 15428
rect 3384 15416 3390 15428
rect 5445 15419 5503 15425
rect 5445 15416 5457 15419
rect 3384 15388 5457 15416
rect 3384 15376 3390 15388
rect 5445 15385 5457 15388
rect 5491 15385 5503 15419
rect 5445 15379 5503 15385
rect 7558 15376 7564 15428
rect 7616 15416 7622 15428
rect 8941 15419 8999 15425
rect 8941 15416 8953 15419
rect 7616 15388 8953 15416
rect 7616 15376 7622 15388
rect 8941 15385 8953 15388
rect 8987 15385 8999 15419
rect 8941 15379 8999 15385
rect 10410 15376 10416 15428
rect 10468 15425 10474 15428
rect 10468 15416 10480 15425
rect 11348 15416 11376 15592
rect 17402 15580 17408 15632
rect 17460 15620 17466 15632
rect 17862 15620 17868 15632
rect 17460 15592 17868 15620
rect 17460 15580 17466 15592
rect 17862 15580 17868 15592
rect 17920 15580 17926 15632
rect 11422 15512 11428 15564
rect 11480 15552 11486 15564
rect 13265 15555 13323 15561
rect 11480 15524 12434 15552
rect 11480 15512 11486 15524
rect 11698 15444 11704 15496
rect 11756 15484 11762 15496
rect 12158 15484 12164 15496
rect 11756 15456 12164 15484
rect 11756 15444 11762 15456
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 12406 15484 12434 15524
rect 13265 15521 13277 15555
rect 13311 15552 13323 15555
rect 15470 15552 15476 15564
rect 13311 15524 15476 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 13280 15484 13308 15515
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 17034 15512 17040 15564
rect 17092 15552 17098 15564
rect 18233 15555 18291 15561
rect 18233 15552 18245 15555
rect 17092 15524 18245 15552
rect 17092 15512 17098 15524
rect 18233 15521 18245 15524
rect 18279 15521 18291 15555
rect 18233 15515 18291 15521
rect 19610 15512 19616 15564
rect 19668 15552 19674 15564
rect 20070 15552 20076 15564
rect 19668 15524 20076 15552
rect 19668 15512 19674 15524
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 12406 15456 13308 15484
rect 13446 15444 13452 15496
rect 13504 15484 13510 15496
rect 16586 15487 16644 15493
rect 16586 15484 16598 15487
rect 13504 15456 16598 15484
rect 13504 15444 13510 15456
rect 16586 15453 16598 15456
rect 16632 15453 16644 15487
rect 16586 15447 16644 15453
rect 16853 15487 16911 15493
rect 16853 15453 16865 15487
rect 16899 15484 16911 15487
rect 16899 15456 17264 15484
rect 16899 15453 16911 15456
rect 16853 15447 16911 15453
rect 10468 15388 10513 15416
rect 11072 15388 11376 15416
rect 10468 15379 10480 15388
rect 10468 15376 10474 15379
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 3234 15348 3240 15360
rect 3195 15320 3240 15348
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 4065 15351 4123 15357
rect 4065 15317 4077 15351
rect 4111 15348 4123 15351
rect 4154 15348 4160 15360
rect 4111 15320 4160 15348
rect 4111 15317 4123 15320
rect 4065 15311 4123 15317
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 4522 15348 4528 15360
rect 4483 15320 4528 15348
rect 4522 15308 4528 15320
rect 4580 15308 4586 15360
rect 4982 15348 4988 15360
rect 4943 15320 4988 15348
rect 4982 15308 4988 15320
rect 5040 15308 5046 15360
rect 5350 15348 5356 15360
rect 5311 15320 5356 15348
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 6549 15351 6607 15357
rect 6549 15317 6561 15351
rect 6595 15348 6607 15351
rect 7101 15351 7159 15357
rect 7101 15348 7113 15351
rect 6595 15320 7113 15348
rect 6595 15317 6607 15320
rect 6549 15311 6607 15317
rect 7101 15317 7113 15320
rect 7147 15317 7159 15351
rect 7101 15311 7159 15317
rect 7926 15308 7932 15360
rect 7984 15348 7990 15360
rect 11072 15348 11100 15388
rect 12342 15376 12348 15428
rect 12400 15416 12406 15428
rect 13633 15419 13691 15425
rect 13633 15416 13645 15419
rect 12400 15388 13645 15416
rect 12400 15376 12406 15388
rect 13633 15385 13645 15388
rect 13679 15416 13691 15419
rect 14093 15419 14151 15425
rect 14093 15416 14105 15419
rect 13679 15388 14105 15416
rect 13679 15385 13691 15388
rect 13633 15379 13691 15385
rect 14093 15385 14105 15388
rect 14139 15416 14151 15419
rect 14274 15416 14280 15428
rect 14139 15388 14280 15416
rect 14139 15385 14151 15388
rect 14093 15379 14151 15385
rect 14274 15376 14280 15388
rect 14332 15416 14338 15428
rect 14829 15419 14887 15425
rect 14829 15416 14841 15419
rect 14332 15388 14841 15416
rect 14332 15376 14338 15388
rect 14829 15385 14841 15388
rect 14875 15385 14887 15419
rect 14829 15379 14887 15385
rect 7984 15320 11100 15348
rect 7984 15308 7990 15320
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 12032 15320 12081 15348
rect 12032 15308 12038 15320
rect 12069 15317 12081 15320
rect 12115 15317 12127 15351
rect 12069 15311 12127 15317
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 12492 15320 12537 15348
rect 12492 15308 12498 15320
rect 12618 15308 12624 15360
rect 12676 15348 12682 15360
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 12676 15320 12817 15348
rect 12676 15308 12682 15320
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 12805 15311 12863 15317
rect 12894 15308 12900 15360
rect 12952 15348 12958 15360
rect 14461 15351 14519 15357
rect 14461 15348 14473 15351
rect 12952 15320 14473 15348
rect 12952 15308 12958 15320
rect 14461 15317 14473 15320
rect 14507 15348 14519 15351
rect 15102 15348 15108 15360
rect 14507 15320 15108 15348
rect 14507 15317 14519 15320
rect 14461 15311 14519 15317
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 15378 15308 15384 15360
rect 15436 15348 15442 15360
rect 17236 15357 17264 15456
rect 17494 15444 17500 15496
rect 17552 15484 17558 15496
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 17552 15456 18153 15484
rect 17552 15444 17558 15456
rect 18141 15453 18153 15456
rect 18187 15484 18199 15487
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18187 15456 18705 15484
rect 18187 15453 18199 15456
rect 18141 15447 18199 15453
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 18693 15447 18751 15453
rect 18966 15444 18972 15496
rect 19024 15484 19030 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19024 15456 19441 15484
rect 19024 15444 19030 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19978 15484 19984 15496
rect 19939 15456 19984 15484
rect 19429 15447 19487 15453
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 20530 15484 20536 15496
rect 20491 15456 20536 15484
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 20990 15444 20996 15496
rect 21048 15484 21054 15496
rect 21085 15487 21143 15493
rect 21085 15484 21097 15487
rect 21048 15456 21097 15484
rect 21048 15444 21054 15456
rect 21085 15453 21097 15456
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 15473 15351 15531 15357
rect 15473 15348 15485 15351
rect 15436 15320 15485 15348
rect 15436 15308 15442 15320
rect 15473 15317 15485 15320
rect 15519 15317 15531 15351
rect 15473 15311 15531 15317
rect 17221 15351 17279 15357
rect 17221 15317 17233 15351
rect 17267 15348 17279 15351
rect 17402 15348 17408 15360
rect 17267 15320 17408 15348
rect 17267 15317 17279 15320
rect 17221 15311 17279 15317
rect 17402 15308 17408 15320
rect 17460 15308 17466 15360
rect 18046 15348 18052 15360
rect 18007 15320 18052 15348
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 19610 15348 19616 15360
rect 19571 15320 19616 15348
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 20162 15348 20168 15360
rect 20123 15320 20168 15348
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 20714 15348 20720 15360
rect 20675 15320 20720 15348
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 21269 15351 21327 15357
rect 21269 15317 21281 15351
rect 21315 15348 21327 15351
rect 21358 15348 21364 15360
rect 21315 15320 21364 15348
rect 21315 15317 21327 15320
rect 21269 15311 21327 15317
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15113 2007 15147
rect 1949 15107 2007 15113
rect 2777 15147 2835 15153
rect 2777 15113 2789 15147
rect 2823 15144 2835 15147
rect 3326 15144 3332 15156
rect 2823 15116 3332 15144
rect 2823 15113 2835 15116
rect 2777 15107 2835 15113
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 1964 15008 1992 15107
rect 3326 15104 3332 15116
rect 3384 15104 3390 15156
rect 3418 15104 3424 15156
rect 3476 15144 3482 15156
rect 3789 15147 3847 15153
rect 3789 15144 3801 15147
rect 3476 15116 3801 15144
rect 3476 15104 3482 15116
rect 3789 15113 3801 15116
rect 3835 15113 3847 15147
rect 3789 15107 3847 15113
rect 4617 15147 4675 15153
rect 4617 15113 4629 15147
rect 4663 15144 4675 15147
rect 4982 15144 4988 15156
rect 4663 15116 4988 15144
rect 4663 15113 4675 15116
rect 4617 15107 4675 15113
rect 4982 15104 4988 15116
rect 5040 15104 5046 15156
rect 11057 15147 11115 15153
rect 7024 15116 10824 15144
rect 2406 15036 2412 15088
rect 2464 15076 2470 15088
rect 5442 15076 5448 15088
rect 2464 15048 5448 15076
rect 2464 15036 2470 15048
rect 5442 15036 5448 15048
rect 5500 15036 5506 15088
rect 5994 15036 6000 15088
rect 6052 15076 6058 15088
rect 7024 15076 7052 15116
rect 10796 15088 10824 15116
rect 11057 15113 11069 15147
rect 11103 15144 11115 15147
rect 11146 15144 11152 15156
rect 11103 15116 11152 15144
rect 11103 15113 11115 15116
rect 11057 15107 11115 15113
rect 11146 15104 11152 15116
rect 11204 15104 11210 15156
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 11296 15116 11529 15144
rect 11296 15104 11302 15116
rect 11517 15113 11529 15116
rect 11563 15144 11575 15147
rect 12342 15144 12348 15156
rect 11563 15116 12348 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 12342 15104 12348 15116
rect 12400 15144 12406 15156
rect 12529 15147 12587 15153
rect 12529 15144 12541 15147
rect 12400 15116 12541 15144
rect 12400 15104 12406 15116
rect 12529 15113 12541 15116
rect 12575 15113 12587 15147
rect 12529 15107 12587 15113
rect 12897 15147 12955 15153
rect 12897 15113 12909 15147
rect 12943 15144 12955 15147
rect 13446 15144 13452 15156
rect 12943 15116 13452 15144
rect 12943 15113 12955 15116
rect 12897 15107 12955 15113
rect 13446 15104 13452 15116
rect 13504 15104 13510 15156
rect 15102 15104 15108 15156
rect 15160 15144 15166 15156
rect 17218 15144 17224 15156
rect 15160 15116 17224 15144
rect 15160 15104 15166 15116
rect 17218 15104 17224 15116
rect 17276 15104 17282 15156
rect 19613 15147 19671 15153
rect 19613 15113 19625 15147
rect 19659 15144 19671 15147
rect 20622 15144 20628 15156
rect 19659 15116 20628 15144
rect 19659 15113 19671 15116
rect 19613 15107 19671 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 6052 15048 7052 15076
rect 6052 15036 6058 15048
rect 7098 15036 7104 15088
rect 7156 15076 7162 15088
rect 9922 15079 9980 15085
rect 9922 15076 9934 15079
rect 7156 15048 9934 15076
rect 7156 15036 7162 15048
rect 2130 15008 2136 15020
rect 1719 14980 1992 15008
rect 2091 14980 2136 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 6914 15008 6920 15020
rect 5675 14980 6920 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 15008 7435 15011
rect 7926 15008 7932 15020
rect 7423 14980 7932 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 7926 14968 7932 14980
rect 7984 15008 7990 15020
rect 8389 15011 8447 15017
rect 8389 15008 8401 15011
rect 7984 14980 8401 15008
rect 7984 14968 7990 14980
rect 8389 14977 8401 14980
rect 8435 14977 8447 15011
rect 8389 14971 8447 14977
rect 9582 14968 9588 15020
rect 9640 15008 9646 15020
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 9640 14980 9689 15008
rect 9640 14968 9646 14980
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 2593 14943 2651 14949
rect 2593 14909 2605 14943
rect 2639 14909 2651 14943
rect 2593 14903 2651 14909
rect 2685 14943 2743 14949
rect 2685 14909 2697 14943
rect 2731 14940 2743 14943
rect 4706 14940 4712 14952
rect 2731 14912 3556 14940
rect 4667 14912 4712 14940
rect 2731 14909 2743 14912
rect 2685 14903 2743 14909
rect 2608 14872 2636 14903
rect 3528 14884 3556 14912
rect 4706 14900 4712 14912
rect 4764 14900 4770 14952
rect 4798 14900 4804 14952
rect 4856 14940 4862 14952
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 4856 14912 4905 14940
rect 4856 14900 4862 14912
rect 4893 14909 4905 14912
rect 4939 14940 4951 14943
rect 5442 14940 5448 14952
rect 4939 14912 5448 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14909 5779 14943
rect 5721 14903 5779 14909
rect 5905 14943 5963 14949
rect 5905 14909 5917 14943
rect 5951 14940 5963 14943
rect 5994 14940 6000 14952
rect 5951 14912 6000 14940
rect 5951 14909 5963 14912
rect 5905 14903 5963 14909
rect 2958 14872 2964 14884
rect 2608 14844 2964 14872
rect 2958 14832 2964 14844
rect 3016 14832 3022 14884
rect 3510 14872 3516 14884
rect 3471 14844 3516 14872
rect 3510 14832 3516 14844
rect 3568 14832 3574 14884
rect 4062 14832 4068 14884
rect 4120 14872 4126 14884
rect 5261 14875 5319 14881
rect 5261 14872 5273 14875
rect 4120 14844 5273 14872
rect 4120 14832 4126 14844
rect 5261 14841 5273 14844
rect 5307 14841 5319 14875
rect 5261 14835 5319 14841
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 3142 14804 3148 14816
rect 3103 14776 3148 14804
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 4246 14804 4252 14816
rect 4207 14776 4252 14804
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 5736 14804 5764 14903
rect 5994 14900 6000 14912
rect 6052 14900 6058 14952
rect 7006 14900 7012 14952
rect 7064 14900 7070 14952
rect 7466 14940 7472 14952
rect 7427 14912 7472 14940
rect 7466 14900 7472 14912
rect 7524 14900 7530 14952
rect 7558 14900 7564 14952
rect 7616 14940 7622 14952
rect 9784 14940 9812 15048
rect 9922 15045 9934 15048
rect 9968 15045 9980 15079
rect 9922 15039 9980 15045
rect 10778 15036 10784 15088
rect 10836 15076 10842 15088
rect 10836 15048 14412 15076
rect 10836 15036 10842 15048
rect 13998 14968 14004 15020
rect 14056 15017 14062 15020
rect 14056 15008 14068 15017
rect 14274 15008 14280 15020
rect 14056 14980 14101 15008
rect 14235 14980 14280 15008
rect 14056 14971 14068 14980
rect 14056 14968 14062 14971
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 14384 15008 14412 15048
rect 15562 15036 15568 15088
rect 15620 15076 15626 15088
rect 19058 15076 19064 15088
rect 15620 15048 16068 15076
rect 15620 15036 15626 15048
rect 16040 15017 16068 15048
rect 17420 15048 19064 15076
rect 17420 15020 17448 15048
rect 19058 15036 19064 15048
rect 19116 15076 19122 15088
rect 21542 15076 21548 15088
rect 19116 15048 19196 15076
rect 19116 15036 19122 15048
rect 15758 15011 15816 15017
rect 15758 15008 15770 15011
rect 14384 14980 15770 15008
rect 15758 14977 15770 14980
rect 15804 14977 15816 15011
rect 15758 14971 15816 14977
rect 16025 15011 16083 15017
rect 16025 14977 16037 15011
rect 16071 15008 16083 15011
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16071 14980 16681 15008
rect 16071 14977 16083 14980
rect 16025 14971 16083 14977
rect 16669 14977 16681 14980
rect 16715 15008 16727 15011
rect 17218 15008 17224 15020
rect 16715 14980 17224 15008
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 17218 14968 17224 14980
rect 17276 15008 17282 15020
rect 17402 15008 17408 15020
rect 17276 14980 17408 15008
rect 17276 14968 17282 14980
rect 17402 14968 17408 14980
rect 17460 14968 17466 15020
rect 18322 14968 18328 15020
rect 18380 15008 18386 15020
rect 18874 15008 18880 15020
rect 18932 15017 18938 15020
rect 19168 15017 19196 15048
rect 20824 15048 21548 15076
rect 18380 14980 18880 15008
rect 18380 14968 18386 14980
rect 18874 14968 18880 14980
rect 18932 15008 18944 15017
rect 19153 15011 19211 15017
rect 18932 14980 18977 15008
rect 18932 14971 18944 14980
rect 19153 14977 19165 15011
rect 19199 14977 19211 15011
rect 20726 15011 20784 15017
rect 20726 15008 20738 15011
rect 19153 14971 19211 14977
rect 19260 14980 20738 15008
rect 18932 14968 18938 14971
rect 7616 14912 7661 14940
rect 8036 14912 9628 14940
rect 7616 14900 7622 14912
rect 6733 14875 6791 14881
rect 6733 14841 6745 14875
rect 6779 14872 6791 14875
rect 7024 14872 7052 14900
rect 8036 14872 8064 14912
rect 6779 14844 8064 14872
rect 6779 14841 6791 14844
rect 6733 14835 6791 14841
rect 8110 14832 8116 14884
rect 8168 14872 8174 14884
rect 8757 14875 8815 14881
rect 8757 14872 8769 14875
rect 8168 14844 8769 14872
rect 8168 14832 8174 14844
rect 8757 14841 8769 14844
rect 8803 14841 8815 14875
rect 8757 14835 8815 14841
rect 7009 14807 7067 14813
rect 7009 14804 7021 14807
rect 5736 14776 7021 14804
rect 7009 14773 7021 14776
rect 7055 14773 7067 14807
rect 7009 14767 7067 14773
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 8021 14807 8079 14813
rect 8021 14804 8033 14807
rect 7524 14776 8033 14804
rect 7524 14764 7530 14776
rect 8021 14773 8033 14776
rect 8067 14804 8079 14807
rect 8202 14804 8208 14816
rect 8067 14776 8208 14804
rect 8067 14773 8079 14776
rect 8021 14767 8079 14773
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 8478 14764 8484 14816
rect 8536 14804 8542 14816
rect 9030 14804 9036 14816
rect 8536 14776 9036 14804
rect 8536 14764 8542 14776
rect 9030 14764 9036 14776
rect 9088 14804 9094 14816
rect 9125 14807 9183 14813
rect 9125 14804 9137 14807
rect 9088 14776 9137 14804
rect 9088 14764 9094 14776
rect 9125 14773 9137 14776
rect 9171 14773 9183 14807
rect 9600 14804 9628 14912
rect 9692 14912 9812 14940
rect 9692 14884 9720 14912
rect 9674 14832 9680 14884
rect 9732 14832 9738 14884
rect 11146 14832 11152 14884
rect 11204 14872 11210 14884
rect 12710 14872 12716 14884
rect 11204 14844 12716 14872
rect 11204 14832 11210 14844
rect 12710 14832 12716 14844
rect 12768 14832 12774 14884
rect 17328 14844 18276 14872
rect 11330 14804 11336 14816
rect 9600 14776 11336 14804
rect 9125 14767 9183 14773
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 11977 14807 12035 14813
rect 11977 14773 11989 14807
rect 12023 14804 12035 14807
rect 12158 14804 12164 14816
rect 12023 14776 12164 14804
rect 12023 14773 12035 14776
rect 11977 14767 12035 14773
rect 12158 14764 12164 14776
rect 12216 14804 12222 14816
rect 14645 14807 14703 14813
rect 14645 14804 14657 14807
rect 12216 14776 14657 14804
rect 12216 14764 12222 14776
rect 14645 14773 14657 14776
rect 14691 14773 14703 14807
rect 14645 14767 14703 14773
rect 16022 14764 16028 14816
rect 16080 14804 16086 14816
rect 17328 14813 17356 14844
rect 17313 14807 17371 14813
rect 17313 14804 17325 14807
rect 16080 14776 17325 14804
rect 16080 14764 16086 14776
rect 17313 14773 17325 14776
rect 17359 14773 17371 14807
rect 17770 14804 17776 14816
rect 17731 14776 17776 14804
rect 17313 14767 17371 14773
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 18248 14804 18276 14844
rect 19260 14804 19288 14980
rect 20726 14977 20738 14980
rect 20772 15008 20784 15011
rect 20824 15008 20852 15048
rect 21542 15036 21548 15048
rect 21600 15036 21606 15088
rect 20772 14980 20852 15008
rect 20772 14977 20784 14980
rect 20726 14971 20784 14977
rect 20898 14968 20904 15020
rect 20956 15008 20962 15020
rect 20993 15011 21051 15017
rect 20993 15008 21005 15011
rect 20956 14980 21005 15008
rect 20956 14968 20962 14980
rect 20993 14977 21005 14980
rect 21039 15008 21051 15011
rect 21266 15008 21272 15020
rect 21039 14980 21272 15008
rect 21039 14977 21051 14980
rect 20993 14971 21051 14977
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 18248 14776 19288 14804
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 7098 14600 7104 14612
rect 3988 14572 7104 14600
rect 3053 14535 3111 14541
rect 3053 14501 3065 14535
rect 3099 14532 3111 14535
rect 3988 14532 4016 14572
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 10410 14600 10416 14612
rect 7524 14572 10272 14600
rect 10371 14572 10416 14600
rect 7524 14560 7530 14572
rect 3099 14504 4016 14532
rect 3099 14501 3111 14504
rect 3053 14495 3111 14501
rect 3068 14464 3096 14495
rect 4062 14492 4068 14544
rect 4120 14532 4126 14544
rect 7837 14535 7895 14541
rect 7837 14532 7849 14535
rect 4120 14504 7849 14532
rect 4120 14492 4126 14504
rect 7837 14501 7849 14504
rect 7883 14501 7895 14535
rect 10244 14532 10272 14572
rect 10410 14560 10416 14572
rect 10468 14560 10474 14612
rect 10689 14603 10747 14609
rect 10689 14569 10701 14603
rect 10735 14600 10747 14603
rect 10778 14600 10784 14612
rect 10735 14572 10784 14600
rect 10735 14569 10747 14572
rect 10689 14563 10747 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 11146 14560 11152 14612
rect 11204 14600 11210 14612
rect 11882 14600 11888 14612
rect 11204 14572 11888 14600
rect 11204 14560 11210 14572
rect 11882 14560 11888 14572
rect 11940 14600 11946 14612
rect 11940 14572 13860 14600
rect 11940 14560 11946 14572
rect 10594 14532 10600 14544
rect 10244 14504 10600 14532
rect 7837 14495 7895 14501
rect 10594 14492 10600 14504
rect 10652 14492 10658 14544
rect 4246 14464 4252 14476
rect 2700 14436 3096 14464
rect 4207 14436 4252 14464
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1946 14396 1952 14408
rect 1719 14368 1952 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2700 14405 2728 14436
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 6086 14464 6092 14476
rect 4479 14436 4936 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4908 14408 4936 14436
rect 5092 14436 6092 14464
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2677 14399 2735 14405
rect 2271 14368 2544 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2038 14260 2044 14272
rect 1999 14232 2044 14260
rect 2038 14220 2044 14232
rect 2096 14220 2102 14272
rect 2516 14269 2544 14368
rect 2677 14365 2689 14399
rect 2723 14365 2735 14399
rect 2677 14359 2735 14365
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 3786 14396 3792 14408
rect 3467 14368 3792 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 4157 14399 4215 14405
rect 4157 14365 4169 14399
rect 4203 14396 4215 14399
rect 4522 14396 4528 14408
rect 4203 14368 4528 14396
rect 4203 14365 4215 14368
rect 4157 14359 4215 14365
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 4890 14396 4896 14408
rect 4851 14368 4896 14396
rect 4890 14356 4896 14368
rect 4948 14356 4954 14408
rect 2746 14300 3832 14328
rect 2746 14272 2774 14300
rect 2501 14263 2559 14269
rect 2501 14229 2513 14263
rect 2547 14229 2559 14263
rect 2501 14223 2559 14229
rect 2682 14220 2688 14272
rect 2740 14232 2774 14272
rect 3804 14269 3832 14300
rect 4798 14288 4804 14340
rect 4856 14328 4862 14340
rect 5092 14328 5120 14436
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 6917 14467 6975 14473
rect 6917 14433 6929 14467
rect 6963 14433 6975 14467
rect 6917 14427 6975 14433
rect 7101 14467 7159 14473
rect 7101 14433 7113 14467
rect 7147 14464 7159 14467
rect 7190 14464 7196 14476
rect 7147 14436 7196 14464
rect 7147 14433 7159 14436
rect 7101 14427 7159 14433
rect 5166 14356 5172 14408
rect 5224 14396 5230 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 5224 14368 6469 14396
rect 5224 14356 5230 14368
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 6932 14396 6960 14427
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 12069 14467 12127 14473
rect 12069 14433 12081 14467
rect 12115 14464 12127 14467
rect 12342 14464 12348 14476
rect 12115 14436 12348 14464
rect 12115 14433 12127 14436
rect 12069 14427 12127 14433
rect 12342 14424 12348 14436
rect 12400 14424 12406 14476
rect 6932 14392 7052 14396
rect 7116 14392 7328 14396
rect 6932 14368 7328 14392
rect 6457 14359 6515 14365
rect 7024 14364 7144 14368
rect 4856 14300 5120 14328
rect 4856 14288 4862 14300
rect 5534 14288 5540 14340
rect 5592 14328 5598 14340
rect 7300 14328 7328 14368
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 9033 14399 9091 14405
rect 9033 14396 9045 14399
rect 8536 14368 9045 14396
rect 8536 14356 8542 14368
rect 9033 14365 9045 14368
rect 9079 14365 9091 14399
rect 11238 14396 11244 14408
rect 9033 14359 9091 14365
rect 9140 14368 11244 14396
rect 9140 14328 9168 14368
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 12612 14399 12670 14405
rect 12612 14365 12624 14399
rect 12658 14396 12670 14399
rect 12894 14396 12900 14408
rect 12658 14368 12900 14396
rect 12658 14365 12670 14368
rect 12612 14359 12670 14365
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 13832 14396 13860 14572
rect 13906 14560 13912 14612
rect 13964 14600 13970 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13964 14572 14105 14600
rect 13964 14560 13970 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 14093 14563 14151 14569
rect 15841 14603 15899 14609
rect 15841 14569 15853 14603
rect 15887 14600 15899 14603
rect 16206 14600 16212 14612
rect 15887 14572 16212 14600
rect 15887 14569 15899 14572
rect 15841 14563 15899 14569
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 16316 14572 18828 14600
rect 15746 14492 15752 14544
rect 15804 14532 15810 14544
rect 16316 14532 16344 14572
rect 15804 14504 16344 14532
rect 15804 14492 15810 14504
rect 15206 14399 15264 14405
rect 15206 14396 15218 14399
rect 13832 14368 15218 14396
rect 15206 14365 15218 14368
rect 15252 14365 15264 14399
rect 15206 14359 15264 14365
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14396 15531 14399
rect 15562 14396 15568 14408
rect 15519 14368 15568 14396
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 16954 14399 17012 14405
rect 16954 14365 16966 14399
rect 17000 14365 17012 14399
rect 17218 14396 17224 14408
rect 17179 14368 17224 14396
rect 16954 14359 17012 14365
rect 9306 14337 9312 14340
rect 9300 14328 9312 14337
rect 5592 14300 7144 14328
rect 7300 14300 9168 14328
rect 9267 14300 9312 14328
rect 5592 14288 5598 14300
rect 3789 14263 3847 14269
rect 2740 14220 2746 14232
rect 3789 14229 3801 14263
rect 3835 14229 3847 14263
rect 5258 14260 5264 14272
rect 5219 14232 5264 14260
rect 3789 14223 3847 14229
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 5442 14220 5448 14272
rect 5500 14260 5506 14272
rect 5813 14263 5871 14269
rect 5813 14260 5825 14263
rect 5500 14232 5825 14260
rect 5500 14220 5506 14232
rect 5813 14229 5825 14232
rect 5859 14260 5871 14263
rect 5902 14260 5908 14272
rect 5859 14232 5908 14260
rect 5859 14229 5871 14232
rect 5813 14223 5871 14229
rect 5902 14220 5908 14232
rect 5960 14220 5966 14272
rect 7116 14260 7144 14300
rect 9300 14291 9312 14300
rect 9306 14288 9312 14291
rect 9364 14288 9370 14340
rect 9416 14300 10824 14328
rect 9416 14272 9444 14300
rect 7193 14263 7251 14269
rect 7193 14260 7205 14263
rect 7116 14232 7205 14260
rect 7193 14229 7205 14232
rect 7239 14229 7251 14263
rect 7558 14260 7564 14272
rect 7519 14232 7564 14260
rect 7193 14223 7251 14229
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 8297 14263 8355 14269
rect 8297 14229 8309 14263
rect 8343 14260 8355 14263
rect 8570 14260 8576 14272
rect 8343 14232 8576 14260
rect 8343 14229 8355 14232
rect 8297 14223 8355 14229
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 9398 14220 9404 14272
rect 9456 14220 9462 14272
rect 10796 14260 10824 14300
rect 11054 14288 11060 14340
rect 11112 14328 11118 14340
rect 11330 14328 11336 14340
rect 11112 14300 11336 14328
rect 11112 14288 11118 14300
rect 11330 14288 11336 14300
rect 11388 14288 11394 14340
rect 11824 14331 11882 14337
rect 11824 14297 11836 14331
rect 11870 14328 11882 14331
rect 12066 14328 12072 14340
rect 11870 14300 12072 14328
rect 11870 14297 11882 14300
rect 11824 14291 11882 14297
rect 12066 14288 12072 14300
rect 12124 14288 12130 14340
rect 16960 14328 16988 14359
rect 17218 14356 17224 14368
rect 17276 14396 17282 14408
rect 17402 14396 17408 14408
rect 17276 14368 17408 14396
rect 17276 14356 17282 14368
rect 17402 14356 17408 14368
rect 17460 14396 17466 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 17460 14368 17509 14396
rect 17460 14356 17466 14368
rect 17497 14365 17509 14368
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 17753 14399 17811 14405
rect 17753 14396 17765 14399
rect 17644 14368 17765 14396
rect 17644 14356 17650 14368
rect 17753 14365 17765 14368
rect 17799 14396 17811 14399
rect 18138 14396 18144 14408
rect 17799 14368 18144 14396
rect 17799 14365 17811 14368
rect 17753 14359 17811 14365
rect 18138 14356 18144 14368
rect 18196 14356 18202 14408
rect 18800 14396 18828 14572
rect 18874 14560 18880 14612
rect 18932 14600 18938 14612
rect 19429 14603 19487 14609
rect 19429 14600 19441 14603
rect 18932 14572 19441 14600
rect 18932 14560 18938 14572
rect 19429 14569 19441 14572
rect 19475 14569 19487 14603
rect 19429 14563 19487 14569
rect 20162 14396 20168 14408
rect 18800 14368 20168 14396
rect 20162 14356 20168 14368
rect 20220 14356 20226 14408
rect 20806 14396 20812 14408
rect 20767 14368 20812 14396
rect 20806 14356 20812 14368
rect 20864 14356 20870 14408
rect 21082 14396 21088 14408
rect 21043 14368 21088 14396
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 17034 14328 17040 14340
rect 12728 14300 14780 14328
rect 16960 14300 17040 14328
rect 12728 14260 12756 14300
rect 13722 14260 13728 14272
rect 10796 14232 12756 14260
rect 13635 14232 13728 14260
rect 13722 14220 13728 14232
rect 13780 14260 13786 14272
rect 13998 14260 14004 14272
rect 13780 14232 14004 14260
rect 13780 14220 13786 14232
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14752 14260 14780 14300
rect 17034 14288 17040 14300
rect 17092 14288 17098 14340
rect 20438 14288 20444 14340
rect 20496 14328 20502 14340
rect 20542 14331 20600 14337
rect 20542 14328 20554 14331
rect 20496 14300 20554 14328
rect 20496 14288 20502 14300
rect 20542 14297 20554 14300
rect 20588 14297 20600 14331
rect 20542 14291 20600 14297
rect 17218 14260 17224 14272
rect 14752 14232 17224 14260
rect 17218 14220 17224 14232
rect 17276 14220 17282 14272
rect 17310 14220 17316 14272
rect 17368 14260 17374 14272
rect 17586 14260 17592 14272
rect 17368 14232 17592 14260
rect 17368 14220 17374 14232
rect 17586 14220 17592 14232
rect 17644 14220 17650 14272
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 18874 14260 18880 14272
rect 18012 14232 18880 14260
rect 18012 14220 18018 14232
rect 18874 14220 18880 14232
rect 18932 14220 18938 14272
rect 21266 14260 21272 14272
rect 21227 14232 21272 14260
rect 21266 14220 21272 14232
rect 21324 14220 21330 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 1946 14056 1952 14068
rect 1907 14028 1952 14056
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 2409 14059 2467 14065
rect 2409 14025 2421 14059
rect 2455 14025 2467 14059
rect 2409 14019 2467 14025
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 2424 13920 2452 14019
rect 3878 14016 3884 14068
rect 3936 14056 3942 14068
rect 3973 14059 4031 14065
rect 3973 14056 3985 14059
rect 3936 14028 3985 14056
rect 3936 14016 3942 14028
rect 3973 14025 3985 14028
rect 4019 14025 4031 14059
rect 3973 14019 4031 14025
rect 4433 14059 4491 14065
rect 4433 14025 4445 14059
rect 4479 14056 4491 14059
rect 5077 14059 5135 14065
rect 5077 14056 5089 14059
rect 4479 14028 5089 14056
rect 4479 14025 4491 14028
rect 4433 14019 4491 14025
rect 5077 14025 5089 14028
rect 5123 14025 5135 14059
rect 5077 14019 5135 14025
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 5537 14059 5595 14065
rect 5537 14056 5549 14059
rect 5500 14028 5549 14056
rect 5500 14016 5506 14028
rect 5537 14025 5549 14028
rect 5583 14025 5595 14059
rect 7098 14056 7104 14068
rect 7059 14028 7104 14056
rect 5537 14019 5595 14025
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 9398 14056 9404 14068
rect 7208 14028 9404 14056
rect 2774 13948 2780 14000
rect 2832 13988 2838 14000
rect 4062 13988 4068 14000
rect 2832 13960 4068 13988
rect 2832 13948 2838 13960
rect 4062 13948 4068 13960
rect 4120 13948 4126 14000
rect 5902 13948 5908 14000
rect 5960 13988 5966 14000
rect 7208 13988 7236 14028
rect 9398 14016 9404 14028
rect 9456 14016 9462 14068
rect 9493 14059 9551 14065
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 9766 14056 9772 14068
rect 9539 14028 9772 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 9766 14016 9772 14028
rect 9824 14056 9830 14068
rect 10594 14056 10600 14068
rect 9824 14028 10600 14056
rect 9824 14016 9830 14028
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 11146 14056 11152 14068
rect 11107 14028 11152 14056
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 14185 14059 14243 14065
rect 14185 14056 14197 14059
rect 12124 14028 14197 14056
rect 12124 14016 12130 14028
rect 14185 14025 14197 14028
rect 14231 14025 14243 14059
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 14185 14019 14243 14025
rect 17402 14016 17408 14028
rect 17460 14056 17466 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 17460 14028 17693 14056
rect 17460 14016 17466 14028
rect 17681 14025 17693 14028
rect 17727 14056 17739 14059
rect 18785 14059 18843 14065
rect 18785 14056 18797 14059
rect 17727 14028 18797 14056
rect 17727 14025 17739 14028
rect 17681 14019 17739 14025
rect 18785 14025 18797 14028
rect 18831 14056 18843 14059
rect 19058 14056 19064 14068
rect 18831 14028 19064 14056
rect 18831 14025 18843 14028
rect 18785 14019 18843 14025
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 19521 14059 19579 14065
rect 19521 14025 19533 14059
rect 19567 14056 19579 14059
rect 20438 14056 20444 14068
rect 19567 14028 20444 14056
rect 19567 14025 19579 14028
rect 19521 14019 19579 14025
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 21177 14059 21235 14065
rect 21177 14056 21189 14059
rect 20548 14028 21189 14056
rect 5960 13960 7236 13988
rect 7377 13991 7435 13997
rect 5960 13948 5966 13960
rect 7377 13957 7389 13991
rect 7423 13988 7435 13991
rect 7834 13988 7840 14000
rect 7423 13960 7840 13988
rect 7423 13957 7435 13960
rect 7377 13951 7435 13957
rect 7834 13948 7840 13960
rect 7892 13948 7898 14000
rect 8380 13991 8438 13997
rect 8380 13957 8392 13991
rect 8426 13988 8438 13991
rect 8846 13988 8852 14000
rect 8426 13960 8852 13988
rect 8426 13957 8438 13960
rect 8380 13951 8438 13957
rect 8846 13948 8852 13960
rect 8904 13948 8910 14000
rect 10036 13991 10094 13997
rect 10036 13957 10048 13991
rect 10082 13988 10094 13991
rect 10134 13988 10140 14000
rect 10082 13960 10140 13988
rect 10082 13957 10094 13960
rect 10036 13951 10094 13957
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 11609 13991 11667 13997
rect 11609 13957 11621 13991
rect 11655 13988 11667 13991
rect 12161 13991 12219 13997
rect 12161 13988 12173 13991
rect 11655 13960 12173 13988
rect 11655 13957 11667 13960
rect 11609 13951 11667 13957
rect 12161 13957 12173 13960
rect 12207 13988 12219 13991
rect 12342 13988 12348 14000
rect 12207 13960 12348 13988
rect 12207 13957 12219 13960
rect 12161 13951 12219 13957
rect 12342 13948 12348 13960
rect 12400 13988 12406 14000
rect 12400 13960 13952 13988
rect 12400 13948 12406 13960
rect 2590 13920 2596 13932
rect 2179 13892 2452 13920
rect 2551 13892 2596 13920
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 1688 13852 1716 13883
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 3050 13920 3056 13932
rect 3011 13892 3056 13920
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 4338 13920 4344 13932
rect 4299 13892 4344 13920
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 4614 13880 4620 13932
rect 4672 13920 4678 13932
rect 5350 13920 5356 13932
rect 4672 13892 5356 13920
rect 4672 13880 4678 13892
rect 5350 13880 5356 13892
rect 5408 13920 5414 13932
rect 5445 13923 5503 13929
rect 5445 13920 5457 13923
rect 5408 13892 5457 13920
rect 5408 13880 5414 13892
rect 5445 13889 5457 13892
rect 5491 13889 5503 13923
rect 5718 13920 5724 13932
rect 5631 13892 5724 13920
rect 5445 13883 5503 13889
rect 5644 13861 5672 13892
rect 5718 13880 5724 13892
rect 5776 13920 5782 13932
rect 5776 13892 6500 13920
rect 5776 13880 5782 13892
rect 4525 13855 4583 13861
rect 1688 13824 2912 13852
rect 2884 13793 2912 13824
rect 4525 13821 4537 13855
rect 4571 13821 4583 13855
rect 4525 13815 4583 13821
rect 5629 13855 5687 13861
rect 5629 13821 5641 13855
rect 5675 13821 5687 13855
rect 5629 13815 5687 13821
rect 2869 13787 2927 13793
rect 2869 13753 2881 13787
rect 2915 13753 2927 13787
rect 2869 13747 2927 13753
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 3326 13676 3332 13728
rect 3384 13716 3390 13728
rect 3421 13719 3479 13725
rect 3421 13716 3433 13719
rect 3384 13688 3433 13716
rect 3384 13676 3390 13688
rect 3421 13685 3433 13688
rect 3467 13685 3479 13719
rect 4540 13716 4568 13815
rect 5902 13812 5908 13864
rect 5960 13852 5966 13864
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 5960 13824 6377 13852
rect 5960 13812 5966 13824
rect 6365 13821 6377 13824
rect 6411 13821 6423 13855
rect 6472 13852 6500 13892
rect 7190 13880 7196 13932
rect 7248 13920 7254 13932
rect 7742 13920 7748 13932
rect 7248 13892 7748 13920
rect 7248 13880 7254 13892
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 9364 13892 12572 13920
rect 9364 13880 9370 13892
rect 7466 13852 7472 13864
rect 6472 13824 7472 13852
rect 6365 13815 6423 13821
rect 7466 13812 7472 13824
rect 7524 13812 7530 13864
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 7883 13824 8125 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 8113 13821 8125 13824
rect 8159 13821 8171 13855
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 8113 13815 8171 13821
rect 9416 13824 9781 13852
rect 5994 13716 6000 13728
rect 4540 13688 6000 13716
rect 3421 13679 3479 13685
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 8128 13716 8156 13815
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 9306 13784 9312 13796
rect 9180 13756 9312 13784
rect 9180 13744 9186 13756
rect 9306 13744 9312 13756
rect 9364 13744 9370 13796
rect 8478 13716 8484 13728
rect 8128 13688 8484 13716
rect 8478 13676 8484 13688
rect 8536 13716 8542 13728
rect 9416 13716 9444 13824
rect 9769 13821 9781 13824
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 12342 13852 12348 13864
rect 11112 13824 12348 13852
rect 11112 13812 11118 13824
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 12544 13793 12572 13892
rect 12710 13880 12716 13932
rect 12768 13920 12774 13932
rect 13642 13923 13700 13929
rect 13642 13920 13654 13923
rect 12768 13892 13654 13920
rect 12768 13880 12774 13892
rect 13642 13889 13654 13892
rect 13688 13889 13700 13923
rect 13642 13883 13700 13889
rect 13814 13880 13820 13932
rect 13872 13920 13878 13932
rect 13924 13929 13952 13960
rect 13998 13948 14004 14000
rect 14056 13988 14062 14000
rect 17310 13988 17316 14000
rect 14056 13960 17316 13988
rect 14056 13948 14062 13960
rect 17310 13948 17316 13960
rect 17368 13948 17374 14000
rect 18046 13948 18052 14000
rect 18104 13988 18110 14000
rect 20548 13988 20576 14028
rect 21177 14025 21189 14028
rect 21223 14025 21235 14059
rect 21177 14019 21235 14025
rect 18104 13960 20576 13988
rect 18104 13948 18110 13960
rect 20622 13948 20628 14000
rect 20680 13997 20686 14000
rect 20680 13988 20692 13997
rect 20680 13960 20725 13988
rect 20680 13951 20692 13960
rect 20680 13948 20686 13951
rect 13909 13923 13967 13929
rect 13909 13920 13921 13923
rect 13872 13892 13921 13920
rect 13872 13880 13878 13892
rect 13909 13889 13921 13892
rect 13955 13889 13967 13923
rect 13909 13883 13967 13889
rect 15286 13880 15292 13932
rect 15344 13929 15350 13932
rect 15344 13920 15356 13929
rect 15344 13892 15389 13920
rect 15344 13883 15356 13892
rect 15344 13880 15350 13883
rect 16114 13880 16120 13932
rect 16172 13920 16178 13932
rect 17037 13923 17095 13929
rect 16172 13892 16896 13920
rect 16172 13880 16178 13892
rect 15562 13852 15568 13864
rect 15523 13824 15568 13852
rect 15562 13812 15568 13824
rect 15620 13852 15626 13864
rect 15841 13855 15899 13861
rect 15841 13852 15853 13855
rect 15620 13824 15853 13852
rect 15620 13812 15626 13824
rect 15841 13821 15853 13824
rect 15887 13852 15899 13855
rect 16209 13855 16267 13861
rect 16209 13852 16221 13855
rect 15887 13824 16221 13852
rect 15887 13821 15899 13824
rect 15841 13815 15899 13821
rect 16209 13821 16221 13824
rect 16255 13821 16267 13855
rect 16868 13852 16896 13892
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 20732 13920 20852 13924
rect 17083 13896 20852 13920
rect 17083 13892 20760 13896
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 16868 13824 18061 13852
rect 16209 13815 16267 13821
rect 18049 13821 18061 13824
rect 18095 13852 18107 13855
rect 19886 13852 19892 13864
rect 18095 13824 19892 13852
rect 18095 13821 18107 13824
rect 18049 13815 18107 13821
rect 19886 13812 19892 13824
rect 19944 13812 19950 13864
rect 20824 13852 20852 13896
rect 20898 13880 20904 13932
rect 20956 13920 20962 13932
rect 21361 13923 21419 13929
rect 21361 13920 21373 13923
rect 20956 13892 21001 13920
rect 21100 13892 21373 13920
rect 20956 13880 20962 13892
rect 21100 13852 21128 13892
rect 21361 13889 21373 13892
rect 21407 13920 21419 13923
rect 21542 13920 21548 13932
rect 21407 13892 21548 13920
rect 21407 13889 21419 13892
rect 21361 13883 21419 13889
rect 21542 13880 21548 13892
rect 21600 13880 21606 13932
rect 20824 13824 21128 13852
rect 12529 13787 12587 13793
rect 12529 13753 12541 13787
rect 12575 13753 12587 13787
rect 12529 13747 12587 13753
rect 17862 13744 17868 13796
rect 17920 13784 17926 13796
rect 18417 13787 18475 13793
rect 18417 13784 18429 13787
rect 17920 13756 18429 13784
rect 17920 13744 17926 13756
rect 18417 13753 18429 13756
rect 18463 13784 18475 13787
rect 19153 13787 19211 13793
rect 19153 13784 19165 13787
rect 18463 13756 19165 13784
rect 18463 13753 18475 13756
rect 18417 13747 18475 13753
rect 19153 13753 19165 13756
rect 19199 13784 19211 13787
rect 19610 13784 19616 13796
rect 19199 13756 19616 13784
rect 19199 13753 19211 13756
rect 19153 13747 19211 13753
rect 19610 13744 19616 13756
rect 19668 13744 19674 13796
rect 20898 13744 20904 13796
rect 20956 13784 20962 13796
rect 21634 13784 21640 13796
rect 20956 13756 21640 13784
rect 20956 13744 20962 13756
rect 21634 13744 21640 13756
rect 21692 13744 21698 13796
rect 8536 13688 9444 13716
rect 8536 13676 8542 13688
rect 9490 13676 9496 13728
rect 9548 13716 9554 13728
rect 11882 13716 11888 13728
rect 9548 13688 11888 13716
rect 9548 13676 9554 13688
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 2556 13484 2820 13512
rect 2556 13472 2562 13484
rect 2225 13447 2283 13453
rect 2225 13413 2237 13447
rect 2271 13444 2283 13447
rect 2406 13444 2412 13456
rect 2271 13416 2412 13444
rect 2271 13413 2283 13416
rect 2225 13407 2283 13413
rect 2406 13404 2412 13416
rect 2464 13404 2470 13456
rect 2682 13404 2688 13456
rect 2740 13404 2746 13456
rect 2700 13317 2728 13404
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 2685 13311 2743 13317
rect 1719 13280 2544 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 2041 13243 2099 13249
rect 2041 13209 2053 13243
rect 2087 13209 2099 13243
rect 2516 13240 2544 13280
rect 2685 13277 2697 13311
rect 2731 13277 2743 13311
rect 2792 13308 2820 13484
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 3145 13515 3203 13521
rect 3145 13512 3157 13515
rect 3108 13484 3157 13512
rect 3108 13472 3114 13484
rect 3145 13481 3157 13484
rect 3191 13481 3203 13515
rect 3145 13475 3203 13481
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4396 13484 4813 13512
rect 4396 13472 4402 13484
rect 4801 13481 4813 13484
rect 4847 13481 4859 13515
rect 4801 13475 4859 13481
rect 5994 13472 6000 13524
rect 6052 13512 6058 13524
rect 6052 13484 9904 13512
rect 6052 13472 6058 13484
rect 5626 13404 5632 13456
rect 5684 13444 5690 13456
rect 7193 13447 7251 13453
rect 7193 13444 7205 13447
rect 5684 13416 7205 13444
rect 5684 13404 5690 13416
rect 7193 13413 7205 13416
rect 7239 13413 7251 13447
rect 9876 13444 9904 13484
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10321 13515 10379 13521
rect 10321 13512 10333 13515
rect 10192 13484 10333 13512
rect 10192 13472 10198 13484
rect 10321 13481 10333 13484
rect 10367 13481 10379 13515
rect 10321 13475 10379 13481
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 13872 13484 14105 13512
rect 13872 13472 13878 13484
rect 14093 13481 14105 13484
rect 14139 13512 14151 13515
rect 15105 13515 15163 13521
rect 15105 13512 15117 13515
rect 14139 13484 15117 13512
rect 14139 13481 14151 13484
rect 14093 13475 14151 13481
rect 15105 13481 15117 13484
rect 15151 13512 15163 13515
rect 15562 13512 15568 13524
rect 15151 13484 15568 13512
rect 15151 13481 15163 13484
rect 15105 13475 15163 13481
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 15838 13512 15844 13524
rect 15799 13484 15844 13512
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 18138 13472 18144 13524
rect 18196 13512 18202 13524
rect 18414 13512 18420 13524
rect 18196 13484 18420 13512
rect 18196 13472 18202 13484
rect 18414 13472 18420 13484
rect 18472 13472 18478 13524
rect 18782 13472 18788 13524
rect 18840 13512 18846 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 18840 13484 18889 13512
rect 18840 13472 18846 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 19058 13472 19064 13524
rect 19116 13512 19122 13524
rect 19337 13515 19395 13521
rect 19337 13512 19349 13515
rect 19116 13484 19349 13512
rect 19116 13472 19122 13484
rect 19337 13481 19349 13484
rect 19383 13512 19395 13515
rect 19426 13512 19432 13524
rect 19383 13484 19432 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19426 13472 19432 13484
rect 19484 13512 19490 13524
rect 20806 13512 20812 13524
rect 19484 13484 20812 13512
rect 19484 13472 19490 13484
rect 20806 13472 20812 13484
rect 20864 13512 20870 13524
rect 20990 13512 20996 13524
rect 20864 13484 20996 13512
rect 20864 13472 20870 13484
rect 20990 13472 20996 13484
rect 21048 13472 21054 13524
rect 11698 13444 11704 13456
rect 9876 13416 11704 13444
rect 7193 13407 7251 13413
rect 11698 13404 11704 13416
rect 11756 13404 11762 13456
rect 11882 13404 11888 13456
rect 11940 13444 11946 13456
rect 14461 13447 14519 13453
rect 14461 13444 14473 13447
rect 11940 13416 14473 13444
rect 11940 13404 11946 13416
rect 14461 13413 14473 13416
rect 14507 13444 14519 13447
rect 15286 13444 15292 13456
rect 14507 13416 15292 13444
rect 14507 13413 14519 13416
rect 14461 13407 14519 13413
rect 15286 13404 15292 13416
rect 15344 13404 15350 13456
rect 20346 13444 20352 13456
rect 20307 13416 20352 13444
rect 20346 13404 20352 13416
rect 20404 13404 20410 13456
rect 5445 13379 5503 13385
rect 5445 13345 5457 13379
rect 5491 13376 5503 13379
rect 5718 13376 5724 13388
rect 5491 13348 5724 13376
rect 5491 13345 5503 13348
rect 5445 13339 5503 13345
rect 5718 13336 5724 13348
rect 5776 13336 5782 13388
rect 6457 13379 6515 13385
rect 6457 13345 6469 13379
rect 6503 13376 6515 13379
rect 6638 13376 6644 13388
rect 6503 13348 6644 13376
rect 6503 13345 6515 13348
rect 6457 13339 6515 13345
rect 6638 13336 6644 13348
rect 6696 13336 6702 13388
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 7006 13376 7012 13388
rect 6963 13348 7012 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 7006 13336 7012 13348
rect 7064 13376 7070 13388
rect 7837 13379 7895 13385
rect 7064 13348 7604 13376
rect 7064 13336 7070 13348
rect 3329 13311 3387 13317
rect 3329 13308 3341 13311
rect 2792 13280 3341 13308
rect 2685 13271 2743 13277
rect 3329 13277 3341 13280
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 3418 13268 3424 13320
rect 3476 13308 3482 13320
rect 5169 13311 5227 13317
rect 3476 13280 4384 13308
rect 3476 13268 3482 13280
rect 3602 13240 3608 13252
rect 2516 13212 3608 13240
rect 2041 13203 2099 13209
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 2056 13172 2084 13203
rect 3602 13200 3608 13212
rect 3660 13200 3666 13252
rect 4356 13249 4384 13280
rect 5169 13277 5181 13311
rect 5215 13308 5227 13311
rect 5258 13308 5264 13320
rect 5215 13280 5264 13308
rect 5215 13277 5227 13280
rect 5169 13271 5227 13277
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13308 6331 13311
rect 7098 13308 7104 13320
rect 6319 13280 7104 13308
rect 6319 13277 6331 13280
rect 6273 13271 6331 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 7576 13317 7604 13348
rect 7837 13345 7849 13379
rect 7883 13345 7895 13379
rect 7837 13339 7895 13345
rect 7561 13311 7619 13317
rect 7561 13277 7573 13311
rect 7607 13308 7619 13311
rect 7650 13308 7656 13320
rect 7607 13280 7656 13308
rect 7607 13277 7619 13280
rect 7561 13271 7619 13277
rect 7650 13268 7656 13280
rect 7708 13268 7714 13320
rect 7852 13308 7880 13339
rect 8478 13336 8484 13388
rect 8536 13376 8542 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8536 13348 8953 13376
rect 8536 13336 8542 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 8956 13308 8984 13339
rect 9950 13336 9956 13388
rect 10008 13376 10014 13388
rect 15470 13376 15476 13388
rect 10008 13348 15476 13376
rect 10008 13336 10014 13348
rect 15470 13336 15476 13348
rect 15528 13336 15534 13388
rect 19610 13336 19616 13388
rect 19668 13376 19674 13388
rect 20622 13376 20628 13388
rect 19668 13348 20628 13376
rect 19668 13336 19674 13348
rect 20622 13336 20628 13348
rect 20680 13376 20686 13388
rect 20901 13379 20959 13385
rect 20901 13376 20913 13379
rect 20680 13348 20913 13376
rect 20680 13336 20686 13348
rect 20901 13345 20913 13348
rect 20947 13345 20959 13379
rect 20901 13339 20959 13345
rect 9030 13308 9036 13320
rect 7852 13280 8524 13308
rect 8943 13280 9036 13308
rect 8496 13252 8524 13280
rect 9030 13268 9036 13280
rect 9088 13308 9094 13320
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 9088 13280 10609 13308
rect 9088 13268 9094 13280
rect 10597 13277 10609 13280
rect 10643 13308 10655 13311
rect 10778 13308 10784 13320
rect 10643 13280 10784 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 10778 13268 10784 13280
rect 10836 13308 10842 13320
rect 10965 13311 11023 13317
rect 10965 13308 10977 13311
rect 10836 13280 10977 13308
rect 10836 13268 10842 13280
rect 10965 13277 10977 13280
rect 11011 13277 11023 13311
rect 12618 13308 12624 13320
rect 10965 13271 11023 13277
rect 11072 13280 12624 13308
rect 4341 13243 4399 13249
rect 4341 13209 4353 13243
rect 4387 13240 4399 13243
rect 5994 13240 6000 13252
rect 4387 13212 6000 13240
rect 4387 13209 4399 13212
rect 4341 13203 4399 13209
rect 5994 13200 6000 13212
rect 6052 13200 6058 13252
rect 6181 13243 6239 13249
rect 6181 13209 6193 13243
rect 6227 13240 6239 13243
rect 7834 13240 7840 13252
rect 6227 13212 7840 13240
rect 6227 13209 6239 13212
rect 6181 13203 6239 13209
rect 7834 13200 7840 13212
rect 7892 13200 7898 13252
rect 8202 13240 8208 13252
rect 8163 13212 8208 13240
rect 8202 13200 8208 13212
rect 8260 13200 8266 13252
rect 8478 13200 8484 13252
rect 8536 13200 8542 13252
rect 9208 13243 9266 13249
rect 9208 13209 9220 13243
rect 9254 13240 9266 13243
rect 11072 13240 11100 13280
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 16206 13268 16212 13320
rect 16264 13308 16270 13320
rect 17221 13311 17279 13317
rect 16264 13280 16896 13308
rect 16264 13268 16270 13280
rect 9254 13212 11100 13240
rect 9254 13209 9266 13212
rect 9208 13203 9266 13209
rect 11146 13200 11152 13252
rect 11204 13240 11210 13252
rect 12805 13243 12863 13249
rect 12805 13240 12817 13243
rect 11204 13212 12817 13240
rect 11204 13200 11210 13212
rect 12805 13209 12817 13212
rect 12851 13209 12863 13243
rect 12805 13203 12863 13209
rect 13725 13243 13783 13249
rect 13725 13209 13737 13243
rect 13771 13240 13783 13243
rect 16868 13240 16896 13280
rect 17221 13277 17233 13311
rect 17267 13308 17279 13311
rect 17402 13308 17408 13320
rect 17267 13280 17408 13308
rect 17267 13277 17279 13280
rect 17221 13271 17279 13277
rect 17402 13268 17408 13280
rect 17460 13308 17466 13320
rect 17497 13311 17555 13317
rect 17497 13308 17509 13311
rect 17460 13280 17509 13308
rect 17460 13268 17466 13280
rect 17497 13277 17509 13280
rect 17543 13277 17555 13311
rect 17497 13271 17555 13277
rect 20073 13311 20131 13317
rect 20073 13277 20085 13311
rect 20119 13308 20131 13311
rect 20254 13308 20260 13320
rect 20119 13280 20260 13308
rect 20119 13277 20131 13280
rect 20073 13271 20131 13277
rect 20254 13268 20260 13280
rect 20312 13268 20318 13320
rect 16954 13243 17012 13249
rect 16954 13240 16966 13243
rect 13771 13212 16804 13240
rect 16868 13212 16966 13240
rect 13771 13209 13783 13212
rect 13725 13203 13783 13209
rect 2774 13172 2780 13184
rect 2056 13144 2780 13172
rect 2774 13132 2780 13144
rect 2832 13132 2838 13184
rect 2869 13175 2927 13181
rect 2869 13141 2881 13175
rect 2915 13172 2927 13175
rect 3786 13172 3792 13184
rect 2915 13144 3792 13172
rect 2915 13141 2927 13144
rect 2869 13135 2927 13141
rect 3786 13132 3792 13144
rect 3844 13132 3850 13184
rect 3973 13175 4031 13181
rect 3973 13141 3985 13175
rect 4019 13172 4031 13175
rect 4062 13172 4068 13184
rect 4019 13144 4068 13172
rect 4019 13141 4031 13144
rect 3973 13135 4031 13141
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 4890 13132 4896 13184
rect 4948 13172 4954 13184
rect 5261 13175 5319 13181
rect 5261 13172 5273 13175
rect 4948 13144 5273 13172
rect 4948 13132 4954 13144
rect 5261 13141 5273 13144
rect 5307 13141 5319 13175
rect 5261 13135 5319 13141
rect 5718 13132 5724 13184
rect 5776 13172 5782 13184
rect 5813 13175 5871 13181
rect 5813 13172 5825 13175
rect 5776 13144 5825 13172
rect 5776 13132 5782 13144
rect 5813 13141 5825 13144
rect 5859 13141 5871 13175
rect 5813 13135 5871 13141
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 7852 13172 7880 13200
rect 9950 13172 9956 13184
rect 7708 13144 7753 13172
rect 7852 13144 9956 13172
rect 7708 13132 7714 13144
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11333 13175 11391 13181
rect 11333 13172 11345 13175
rect 11112 13144 11345 13172
rect 11112 13132 11118 13144
rect 11333 13141 11345 13144
rect 11379 13141 11391 13175
rect 11333 13135 11391 13141
rect 11793 13175 11851 13181
rect 11793 13141 11805 13175
rect 11839 13172 11851 13175
rect 11882 13172 11888 13184
rect 11839 13144 11888 13172
rect 11839 13141 11851 13144
rect 11793 13135 11851 13141
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 12161 13175 12219 13181
rect 12161 13141 12173 13175
rect 12207 13172 12219 13175
rect 12434 13172 12440 13184
rect 12207 13144 12440 13172
rect 12207 13141 12219 13144
rect 12161 13135 12219 13141
rect 12434 13132 12440 13144
rect 12492 13132 12498 13184
rect 12529 13175 12587 13181
rect 12529 13141 12541 13175
rect 12575 13172 12587 13175
rect 12710 13172 12716 13184
rect 12575 13144 12716 13172
rect 12575 13141 12587 13144
rect 12529 13135 12587 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 13265 13175 13323 13181
rect 13265 13172 13277 13175
rect 13136 13144 13277 13172
rect 13136 13132 13142 13144
rect 13265 13141 13277 13144
rect 13311 13141 13323 13175
rect 15562 13172 15568 13184
rect 15523 13144 15568 13172
rect 13265 13135 13323 13141
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 16776 13172 16804 13212
rect 16954 13209 16966 13212
rect 17000 13209 17012 13243
rect 16954 13203 17012 13209
rect 17764 13243 17822 13249
rect 17764 13209 17776 13243
rect 17810 13240 17822 13243
rect 18414 13240 18420 13252
rect 17810 13212 18420 13240
rect 17810 13209 17822 13212
rect 17764 13203 17822 13209
rect 18414 13200 18420 13212
rect 18472 13240 18478 13252
rect 19518 13240 19524 13252
rect 18472 13212 19524 13240
rect 18472 13200 18478 13212
rect 19518 13200 19524 13212
rect 19576 13200 19582 13252
rect 18322 13172 18328 13184
rect 16776 13144 18328 13172
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 19886 13172 19892 13184
rect 19847 13144 19892 13172
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 20622 13132 20628 13184
rect 20680 13172 20686 13184
rect 20717 13175 20775 13181
rect 20717 13172 20729 13175
rect 20680 13144 20729 13172
rect 20680 13132 20686 13144
rect 20717 13141 20729 13144
rect 20763 13141 20775 13175
rect 20717 13135 20775 13141
rect 20806 13132 20812 13184
rect 20864 13172 20870 13184
rect 20864 13144 20909 13172
rect 20864 13132 20870 13144
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 2317 12971 2375 12977
rect 2317 12937 2329 12971
rect 2363 12968 2375 12971
rect 2590 12968 2596 12980
rect 2363 12940 2596 12968
rect 2363 12937 2375 12940
rect 2317 12931 2375 12937
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 2869 12971 2927 12977
rect 2869 12937 2881 12971
rect 2915 12968 2927 12971
rect 3418 12968 3424 12980
rect 2915 12940 3424 12968
rect 2915 12937 2927 12940
rect 2869 12931 2927 12937
rect 3418 12928 3424 12940
rect 3476 12928 3482 12980
rect 3602 12968 3608 12980
rect 3563 12940 3608 12968
rect 3602 12928 3608 12940
rect 3660 12928 3666 12980
rect 4522 12968 4528 12980
rect 4483 12940 4528 12968
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 4706 12928 4712 12980
rect 4764 12968 4770 12980
rect 5261 12971 5319 12977
rect 5261 12968 5273 12971
rect 4764 12940 5273 12968
rect 4764 12928 4770 12940
rect 5261 12937 5273 12940
rect 5307 12937 5319 12971
rect 5718 12968 5724 12980
rect 5679 12940 5724 12968
rect 5261 12931 5319 12937
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 10778 12968 10784 12980
rect 5828 12940 10456 12968
rect 10739 12940 10784 12968
rect 5828 12900 5856 12940
rect 2746 12872 5856 12900
rect 7469 12903 7527 12909
rect 1946 12832 1952 12844
rect 1907 12804 1952 12832
rect 1946 12792 1952 12804
rect 2004 12792 2010 12844
rect 2038 12792 2044 12844
rect 2096 12832 2102 12844
rect 2746 12832 2774 12872
rect 7469 12869 7481 12903
rect 7515 12900 7527 12903
rect 7650 12900 7656 12912
rect 7515 12872 7656 12900
rect 7515 12869 7527 12872
rect 7469 12863 7527 12869
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 9766 12860 9772 12912
rect 9824 12900 9830 12912
rect 10226 12900 10232 12912
rect 10284 12909 10290 12912
rect 9824 12872 10232 12900
rect 9824 12860 9830 12872
rect 10226 12860 10232 12872
rect 10284 12900 10296 12909
rect 10284 12872 10329 12900
rect 10284 12863 10296 12872
rect 10284 12860 10290 12863
rect 2096 12804 2774 12832
rect 2961 12835 3019 12841
rect 2096 12792 2102 12804
rect 2961 12801 2973 12835
rect 3007 12832 3019 12835
rect 3050 12832 3056 12844
rect 3007 12804 3056 12832
rect 3007 12801 3019 12804
rect 2961 12795 3019 12801
rect 3050 12792 3056 12804
rect 3108 12832 3114 12844
rect 3510 12832 3516 12844
rect 3108 12804 3516 12832
rect 3108 12792 3114 12804
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 3786 12832 3792 12844
rect 3747 12804 3792 12832
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 4062 12832 4068 12844
rect 4023 12804 4068 12832
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12832 5043 12835
rect 5074 12832 5080 12844
rect 5031 12804 5080 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12832 5687 12835
rect 5718 12832 5724 12844
rect 5675 12804 5724 12832
rect 5675 12801 5687 12804
rect 5629 12795 5687 12801
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 7834 12832 7840 12844
rect 7607 12804 7840 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 7834 12792 7840 12804
rect 7892 12832 7898 12844
rect 8113 12835 8171 12841
rect 8113 12832 8125 12835
rect 7892 12804 8125 12832
rect 7892 12792 7898 12804
rect 8113 12801 8125 12804
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 1673 12767 1731 12773
rect 1673 12733 1685 12767
rect 1719 12733 1731 12767
rect 1854 12764 1860 12776
rect 1815 12736 1860 12764
rect 1673 12727 1731 12733
rect 1688 12628 1716 12727
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 2866 12764 2872 12776
rect 2823 12736 2872 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 2866 12724 2872 12736
rect 2924 12724 2930 12776
rect 3326 12724 3332 12776
rect 3384 12764 3390 12776
rect 4338 12764 4344 12776
rect 3384 12736 4344 12764
rect 3384 12724 3390 12736
rect 4338 12724 4344 12736
rect 4396 12724 4402 12776
rect 5092 12764 5120 12792
rect 5442 12764 5448 12776
rect 5092 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12764 5506 12776
rect 5813 12767 5871 12773
rect 5813 12764 5825 12767
rect 5500 12736 5825 12764
rect 5500 12724 5506 12736
rect 5813 12733 5825 12736
rect 5859 12733 5871 12767
rect 7282 12764 7288 12776
rect 5813 12727 5871 12733
rect 5920 12736 7288 12764
rect 5534 12696 5540 12708
rect 2746 12668 5540 12696
rect 2746 12628 2774 12668
rect 5534 12656 5540 12668
rect 5592 12656 5598 12708
rect 3326 12628 3332 12640
rect 1688 12600 2774 12628
rect 3287 12600 3332 12628
rect 3326 12588 3332 12600
rect 3384 12588 3390 12640
rect 4249 12631 4307 12637
rect 4249 12597 4261 12631
rect 4295 12628 4307 12631
rect 5920 12628 5948 12736
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12764 7803 12767
rect 9306 12764 9312 12776
rect 7791 12736 9312 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 5994 12656 6000 12708
rect 6052 12696 6058 12708
rect 7760 12696 7788 12727
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 10428 12764 10456 12940
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 12618 12928 12624 12980
rect 12676 12968 12682 12980
rect 13081 12971 13139 12977
rect 13081 12968 13093 12971
rect 12676 12940 13093 12968
rect 12676 12928 12682 12940
rect 13081 12937 13093 12940
rect 13127 12937 13139 12971
rect 13081 12931 13139 12937
rect 14921 12971 14979 12977
rect 14921 12937 14933 12971
rect 14967 12937 14979 12971
rect 14921 12931 14979 12937
rect 10505 12835 10563 12841
rect 10505 12801 10517 12835
rect 10551 12832 10563 12835
rect 10796 12832 10824 12928
rect 13357 12903 13415 12909
rect 13357 12900 13369 12903
rect 11716 12872 13369 12900
rect 11716 12841 11744 12872
rect 13357 12869 13369 12872
rect 13403 12900 13415 12903
rect 13814 12900 13820 12912
rect 13403 12872 13820 12900
rect 13403 12869 13415 12872
rect 13357 12863 13415 12869
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 11701 12835 11759 12841
rect 11701 12832 11713 12835
rect 10551 12804 11713 12832
rect 10551 12801 10563 12804
rect 10505 12795 10563 12801
rect 11701 12801 11713 12804
rect 11747 12801 11759 12835
rect 11957 12835 12015 12841
rect 11957 12832 11969 12835
rect 11701 12795 11759 12801
rect 11808 12804 11969 12832
rect 11146 12764 11152 12776
rect 10428 12736 11152 12764
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 11238 12724 11244 12776
rect 11296 12764 11302 12776
rect 11808 12764 11836 12804
rect 11957 12801 11969 12804
rect 12003 12801 12015 12835
rect 11957 12795 12015 12801
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 14936 12832 14964 12931
rect 15470 12928 15476 12980
rect 15528 12968 15534 12980
rect 18506 12968 18512 12980
rect 15528 12940 18512 12968
rect 15528 12928 15534 12940
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 19153 12971 19211 12977
rect 19153 12968 19165 12971
rect 18748 12940 19165 12968
rect 18748 12928 18754 12940
rect 19153 12937 19165 12940
rect 19199 12937 19211 12971
rect 19426 12968 19432 12980
rect 19387 12940 19432 12968
rect 19153 12931 19211 12937
rect 17034 12860 17040 12912
rect 17092 12900 17098 12912
rect 17218 12900 17224 12912
rect 17092 12872 17224 12900
rect 17092 12860 17098 12872
rect 17218 12860 17224 12872
rect 17276 12860 17282 12912
rect 18040 12903 18098 12909
rect 18040 12869 18052 12903
rect 18086 12900 18098 12903
rect 18782 12900 18788 12912
rect 18086 12872 18788 12900
rect 18086 12869 18098 12872
rect 18040 12863 18098 12869
rect 18782 12860 18788 12872
rect 18840 12860 18846 12912
rect 19168 12900 19196 12931
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 20257 12971 20315 12977
rect 20257 12937 20269 12971
rect 20303 12968 20315 12971
rect 20530 12968 20536 12980
rect 20303 12940 20536 12968
rect 20303 12937 20315 12940
rect 20257 12931 20315 12937
rect 20530 12928 20536 12940
rect 20588 12928 20594 12980
rect 19610 12900 19616 12912
rect 19168 12872 19616 12900
rect 19610 12860 19616 12872
rect 19668 12860 19674 12912
rect 19720 12872 20852 12900
rect 16034 12835 16092 12841
rect 16034 12832 16046 12835
rect 12400 12804 14964 12832
rect 15111 12804 16046 12832
rect 12400 12792 12406 12804
rect 14642 12764 14648 12776
rect 11296 12736 11836 12764
rect 14555 12736 14648 12764
rect 11296 12724 11302 12736
rect 14642 12724 14648 12736
rect 14700 12764 14706 12776
rect 15111 12764 15139 12804
rect 16034 12801 16046 12804
rect 16080 12801 16092 12835
rect 16034 12795 16092 12801
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 19720 12832 19748 12872
rect 17552 12804 19748 12832
rect 17552 12792 17558 12804
rect 19978 12792 19984 12844
rect 20036 12832 20042 12844
rect 20824 12841 20852 12872
rect 20073 12835 20131 12841
rect 20073 12832 20085 12835
rect 20036 12804 20085 12832
rect 20036 12792 20042 12804
rect 20073 12801 20085 12804
rect 20119 12801 20131 12835
rect 20073 12795 20131 12801
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12801 20867 12835
rect 20809 12795 20867 12801
rect 14700 12736 15139 12764
rect 16301 12767 16359 12773
rect 14700 12724 14706 12736
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 17773 12767 17831 12773
rect 17773 12764 17785 12767
rect 16347 12736 16620 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 6052 12668 7788 12696
rect 8573 12699 8631 12705
rect 6052 12656 6058 12668
rect 8573 12665 8585 12699
rect 8619 12696 8631 12699
rect 8619 12668 9628 12696
rect 8619 12665 8631 12668
rect 8573 12659 8631 12665
rect 6638 12628 6644 12640
rect 4295 12600 5948 12628
rect 6599 12600 6644 12628
rect 4295 12597 4307 12600
rect 4249 12591 4307 12597
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 7098 12628 7104 12640
rect 7059 12600 7104 12628
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 9125 12631 9183 12637
rect 9125 12628 9137 12631
rect 8720 12600 9137 12628
rect 8720 12588 8726 12600
rect 9125 12597 9137 12600
rect 9171 12628 9183 12631
rect 9490 12628 9496 12640
rect 9171 12600 9496 12628
rect 9171 12597 9183 12600
rect 9125 12591 9183 12597
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 9600 12628 9628 12668
rect 13722 12656 13728 12708
rect 13780 12696 13786 12708
rect 14185 12699 14243 12705
rect 14185 12696 14197 12699
rect 13780 12668 14197 12696
rect 13780 12656 13786 12668
rect 14185 12665 14197 12668
rect 14231 12696 14243 12699
rect 14274 12696 14280 12708
rect 14231 12668 14280 12696
rect 14231 12665 14243 12668
rect 14185 12659 14243 12665
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 16592 12640 16620 12736
rect 17420 12736 17785 12764
rect 17420 12640 17448 12736
rect 17773 12733 17785 12736
rect 17819 12733 17831 12767
rect 17773 12727 17831 12733
rect 18782 12724 18788 12776
rect 18840 12764 18846 12776
rect 20530 12764 20536 12776
rect 18840 12736 20536 12764
rect 18840 12724 18846 12736
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 19518 12656 19524 12708
rect 19576 12696 19582 12708
rect 19978 12696 19984 12708
rect 19576 12668 19984 12696
rect 19576 12656 19582 12668
rect 19978 12656 19984 12668
rect 20036 12656 20042 12708
rect 16482 12628 16488 12640
rect 9600 12600 16488 12628
rect 16482 12588 16488 12600
rect 16540 12588 16546 12640
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 16761 12631 16819 12637
rect 16761 12628 16773 12631
rect 16632 12600 16773 12628
rect 16632 12588 16638 12600
rect 16761 12597 16773 12600
rect 16807 12628 16819 12631
rect 17313 12631 17371 12637
rect 17313 12628 17325 12631
rect 16807 12600 17325 12628
rect 16807 12597 16819 12600
rect 16761 12591 16819 12597
rect 17313 12597 17325 12600
rect 17359 12628 17371 12631
rect 17402 12628 17408 12640
rect 17359 12600 17408 12628
rect 17359 12597 17371 12600
rect 17313 12591 17371 12597
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 4522 12424 4528 12436
rect 1728 12396 4528 12424
rect 1728 12384 1734 12396
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 8021 12427 8079 12433
rect 8021 12424 8033 12427
rect 6880 12396 8033 12424
rect 6880 12384 6886 12396
rect 8021 12393 8033 12396
rect 8067 12393 8079 12427
rect 8021 12387 8079 12393
rect 8110 12384 8116 12436
rect 8168 12424 8174 12436
rect 8168 12396 10180 12424
rect 8168 12384 8174 12396
rect 2866 12356 2872 12368
rect 1872 12328 2872 12356
rect 1872 12220 1900 12328
rect 2866 12316 2872 12328
rect 2924 12356 2930 12368
rect 7653 12359 7711 12365
rect 7653 12356 7665 12359
rect 2924 12328 7665 12356
rect 2924 12316 2930 12328
rect 7653 12325 7665 12328
rect 7699 12325 7711 12359
rect 7653 12319 7711 12325
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 8389 12359 8447 12365
rect 8389 12356 8401 12359
rect 8352 12328 8401 12356
rect 8352 12316 8358 12328
rect 8389 12325 8401 12328
rect 8435 12325 8447 12359
rect 8389 12319 8447 12325
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2130 12288 2136 12300
rect 1995 12260 2136 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 2406 12248 2412 12300
rect 2464 12288 2470 12300
rect 2593 12291 2651 12297
rect 2593 12288 2605 12291
rect 2464 12260 2605 12288
rect 2464 12248 2470 12260
rect 2593 12257 2605 12260
rect 2639 12257 2651 12291
rect 2593 12251 2651 12257
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 3142 12288 3148 12300
rect 2823 12260 3148 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 4341 12291 4399 12297
rect 4341 12288 4353 12291
rect 3252 12260 4353 12288
rect 2225 12223 2283 12229
rect 2225 12220 2237 12223
rect 1872 12192 2237 12220
rect 2225 12189 2237 12192
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 3252 12220 3280 12260
rect 4341 12257 4353 12260
rect 4387 12257 4399 12291
rect 4341 12251 4399 12257
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 5994 12288 6000 12300
rect 5307 12260 6000 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12257 6883 12291
rect 6825 12251 6883 12257
rect 6917 12291 6975 12297
rect 6917 12257 6929 12291
rect 6963 12288 6975 12291
rect 7098 12288 7104 12300
rect 6963 12260 7104 12288
rect 6963 12257 6975 12260
rect 6917 12251 6975 12257
rect 3016 12192 3280 12220
rect 4157 12223 4215 12229
rect 3016 12180 3022 12192
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4798 12220 4804 12232
rect 4203 12192 4804 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 6840 12220 6868 12251
rect 7098 12248 7104 12260
rect 7156 12248 7162 12300
rect 10152 12288 10180 12396
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 11149 12427 11207 12433
rect 11149 12424 11161 12427
rect 10928 12396 11161 12424
rect 10928 12384 10934 12396
rect 11149 12393 11161 12396
rect 11195 12393 11207 12427
rect 11149 12387 11207 12393
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 11882 12424 11888 12436
rect 11664 12396 11888 12424
rect 11664 12384 11670 12396
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 13725 12427 13783 12433
rect 13725 12393 13737 12427
rect 13771 12424 13783 12427
rect 14458 12424 14464 12436
rect 13771 12396 14464 12424
rect 13771 12393 13783 12396
rect 13725 12387 13783 12393
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 16574 12424 16580 12436
rect 14844 12396 16580 12424
rect 10505 12359 10563 12365
rect 10505 12325 10517 12359
rect 10551 12356 10563 12359
rect 12158 12356 12164 12368
rect 10551 12328 12164 12356
rect 10551 12325 10563 12328
rect 10505 12319 10563 12325
rect 12158 12316 12164 12328
rect 12216 12316 12222 12368
rect 13814 12356 13820 12368
rect 12406 12328 13820 12356
rect 12406 12288 12434 12328
rect 13814 12316 13820 12328
rect 13872 12356 13878 12368
rect 14642 12356 14648 12368
rect 13872 12328 14648 12356
rect 13872 12316 13878 12328
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 10152 12260 12434 12288
rect 12989 12291 13047 12297
rect 12989 12257 13001 12291
rect 13035 12288 13047 12291
rect 13446 12288 13452 12300
rect 13035 12260 13452 12288
rect 13035 12257 13047 12260
rect 12989 12251 13047 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 13722 12248 13728 12300
rect 13780 12288 13786 12300
rect 14844 12297 14872 12396
rect 16574 12384 16580 12396
rect 16632 12384 16638 12436
rect 17402 12384 17408 12436
rect 17460 12384 17466 12436
rect 18138 12384 18144 12436
rect 18196 12424 18202 12436
rect 18785 12427 18843 12433
rect 18785 12424 18797 12427
rect 18196 12396 18797 12424
rect 18196 12384 18202 12396
rect 18785 12393 18797 12396
rect 18831 12424 18843 12427
rect 19058 12424 19064 12436
rect 18831 12396 19064 12424
rect 18831 12393 18843 12396
rect 18785 12387 18843 12393
rect 19058 12384 19064 12396
rect 19116 12384 19122 12436
rect 19705 12427 19763 12433
rect 19705 12393 19717 12427
rect 19751 12424 19763 12427
rect 19794 12424 19800 12436
rect 19751 12396 19800 12424
rect 19751 12393 19763 12396
rect 19705 12387 19763 12393
rect 19794 12384 19800 12396
rect 19852 12384 19858 12436
rect 20070 12384 20076 12436
rect 20128 12424 20134 12436
rect 20346 12424 20352 12436
rect 20128 12396 20352 12424
rect 20128 12384 20134 12396
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 20809 12427 20867 12433
rect 20809 12393 20821 12427
rect 20855 12424 20867 12427
rect 20990 12424 20996 12436
rect 20855 12396 20996 12424
rect 20855 12393 20867 12396
rect 20809 12387 20867 12393
rect 20990 12384 20996 12396
rect 21048 12384 21054 12436
rect 21174 12424 21180 12436
rect 21135 12396 21180 12424
rect 21174 12384 21180 12396
rect 21232 12384 21238 12436
rect 16209 12359 16267 12365
rect 16209 12325 16221 12359
rect 16255 12356 16267 12359
rect 16942 12356 16948 12368
rect 16255 12328 16948 12356
rect 16255 12325 16267 12328
rect 16209 12319 16267 12325
rect 16942 12316 16948 12328
rect 17000 12316 17006 12368
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 13780 12260 14197 12288
rect 13780 12248 13786 12260
rect 14185 12257 14197 12260
rect 14231 12288 14243 12291
rect 14553 12291 14611 12297
rect 14553 12288 14565 12291
rect 14231 12260 14565 12288
rect 14231 12257 14243 12260
rect 14185 12251 14243 12257
rect 14553 12257 14565 12260
rect 14599 12288 14611 12291
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 14599 12260 14841 12288
rect 14599 12257 14611 12260
rect 14553 12251 14611 12257
rect 14829 12257 14841 12260
rect 14875 12257 14887 12291
rect 14829 12251 14887 12257
rect 9122 12220 9128 12232
rect 6840 12192 8984 12220
rect 9083 12192 9128 12220
rect 2869 12155 2927 12161
rect 2869 12152 2881 12155
rect 2746 12124 2881 12152
rect 2590 12044 2596 12096
rect 2648 12084 2654 12096
rect 2746 12084 2774 12124
rect 2869 12121 2881 12124
rect 2915 12121 2927 12155
rect 2869 12115 2927 12121
rect 5445 12155 5503 12161
rect 5445 12121 5457 12155
rect 5491 12152 5503 12155
rect 6089 12155 6147 12161
rect 6089 12152 6101 12155
rect 5491 12124 6101 12152
rect 5491 12121 5503 12124
rect 5445 12115 5503 12121
rect 6089 12121 6101 12124
rect 6135 12121 6147 12155
rect 7009 12155 7067 12161
rect 7009 12152 7021 12155
rect 6089 12115 6147 12121
rect 6472 12124 7021 12152
rect 3234 12084 3240 12096
rect 2648 12056 2774 12084
rect 3195 12056 3240 12084
rect 2648 12044 2654 12056
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12084 3847 12087
rect 4062 12084 4068 12096
rect 3835 12056 4068 12084
rect 3835 12053 3847 12056
rect 3789 12047 3847 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 4249 12087 4307 12093
rect 4249 12053 4261 12087
rect 4295 12084 4307 12087
rect 4338 12084 4344 12096
rect 4295 12056 4344 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 5350 12084 5356 12096
rect 5311 12056 5356 12084
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5813 12087 5871 12093
rect 5813 12053 5825 12087
rect 5859 12084 5871 12087
rect 6472 12084 6500 12124
rect 7009 12121 7021 12124
rect 7055 12121 7067 12155
rect 7009 12115 7067 12121
rect 7190 12112 7196 12164
rect 7248 12152 7254 12164
rect 7558 12152 7564 12164
rect 7248 12124 7564 12152
rect 7248 12112 7254 12124
rect 7558 12112 7564 12124
rect 7616 12112 7622 12164
rect 5859 12056 6500 12084
rect 7377 12087 7435 12093
rect 5859 12053 5871 12056
rect 5813 12047 5871 12053
rect 7377 12053 7389 12087
rect 7423 12084 7435 12087
rect 7926 12084 7932 12096
rect 7423 12056 7932 12084
rect 7423 12053 7435 12056
rect 7377 12047 7435 12053
rect 7926 12044 7932 12056
rect 7984 12044 7990 12096
rect 8956 12084 8984 12192
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 13262 12220 13268 12232
rect 9223 12192 13268 12220
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 9223 12152 9251 12192
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 13630 12180 13636 12232
rect 13688 12180 13694 12232
rect 15096 12223 15154 12229
rect 15096 12189 15108 12223
rect 15142 12220 15154 12223
rect 15378 12220 15384 12232
rect 15142 12192 15384 12220
rect 15142 12189 15154 12192
rect 15096 12183 15154 12189
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 17420 12229 17448 12384
rect 19429 12359 19487 12365
rect 19429 12325 19441 12359
rect 19475 12356 19487 12359
rect 21082 12356 21088 12368
rect 19475 12328 21088 12356
rect 19475 12325 19487 12328
rect 19429 12319 19487 12325
rect 21082 12316 21088 12328
rect 21140 12316 21146 12368
rect 18782 12248 18788 12300
rect 18840 12288 18846 12300
rect 20349 12291 20407 12297
rect 18840 12260 20024 12288
rect 18840 12248 18846 12260
rect 17405 12223 17463 12229
rect 17405 12189 17417 12223
rect 17451 12220 17463 12223
rect 19245 12223 19303 12229
rect 17451 12192 17908 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 9088 12124 9251 12152
rect 9392 12155 9450 12161
rect 9088 12112 9094 12124
rect 9392 12121 9404 12155
rect 9438 12152 9450 12155
rect 9858 12152 9864 12164
rect 9438 12124 9864 12152
rect 9438 12121 9450 12124
rect 9392 12115 9450 12121
rect 9858 12112 9864 12124
rect 9916 12152 9922 12164
rect 10781 12155 10839 12161
rect 10781 12152 10793 12155
rect 9916 12124 10793 12152
rect 9916 12112 9922 12124
rect 10781 12121 10793 12124
rect 10827 12121 10839 12155
rect 10781 12115 10839 12121
rect 11606 12112 11612 12164
rect 11664 12152 11670 12164
rect 12066 12152 12072 12164
rect 11664 12124 12072 12152
rect 11664 12112 11670 12124
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 12621 12155 12679 12161
rect 12621 12121 12633 12155
rect 12667 12152 12679 12155
rect 13648 12152 13676 12180
rect 17880 12164 17908 12192
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 19886 12220 19892 12232
rect 19291 12192 19892 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 19886 12180 19892 12192
rect 19944 12180 19950 12232
rect 19996 12220 20024 12260
rect 20349 12257 20361 12291
rect 20395 12288 20407 12291
rect 20438 12288 20444 12300
rect 20395 12260 20444 12288
rect 20395 12257 20407 12260
rect 20349 12251 20407 12257
rect 20438 12248 20444 12260
rect 20496 12248 20502 12300
rect 21266 12220 21272 12232
rect 19996 12192 21272 12220
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 15930 12152 15936 12164
rect 12667 12124 13584 12152
rect 13648 12124 15936 12152
rect 12667 12121 12679 12124
rect 12621 12115 12679 12121
rect 10042 12084 10048 12096
rect 8956 12056 10048 12084
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 11054 12044 11060 12096
rect 11112 12084 11118 12096
rect 11517 12087 11575 12093
rect 11517 12084 11529 12087
rect 11112 12056 11529 12084
rect 11112 12044 11118 12056
rect 11517 12053 11529 12056
rect 11563 12053 11575 12087
rect 11974 12084 11980 12096
rect 11935 12056 11980 12084
rect 11517 12047 11575 12053
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 13354 12084 13360 12096
rect 13315 12056 13360 12084
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 13556 12084 13584 12124
rect 15930 12112 15936 12124
rect 15988 12112 15994 12164
rect 17218 12112 17224 12164
rect 17276 12152 17282 12164
rect 17650 12155 17708 12161
rect 17650 12152 17662 12155
rect 17276 12124 17662 12152
rect 17276 12112 17282 12124
rect 17650 12121 17662 12124
rect 17696 12121 17708 12155
rect 17650 12115 17708 12121
rect 17862 12112 17868 12164
rect 17920 12112 17926 12164
rect 20073 12155 20131 12161
rect 20073 12152 20085 12155
rect 17972 12124 20085 12152
rect 16022 12084 16028 12096
rect 13556 12056 16028 12084
rect 16022 12044 16028 12056
rect 16080 12044 16086 12096
rect 17034 12084 17040 12096
rect 16995 12056 17040 12084
rect 17034 12044 17040 12056
rect 17092 12084 17098 12096
rect 17972 12084 18000 12124
rect 20073 12121 20085 12124
rect 20119 12121 20131 12155
rect 20073 12115 20131 12121
rect 17092 12056 18000 12084
rect 17092 12044 17098 12056
rect 20162 12044 20168 12096
rect 20220 12084 20226 12096
rect 20220 12056 20265 12084
rect 20220 12044 20226 12056
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 1854 11840 1860 11892
rect 1912 11880 1918 11892
rect 2501 11883 2559 11889
rect 2501 11880 2513 11883
rect 1912 11852 2513 11880
rect 1912 11840 1918 11852
rect 2501 11849 2513 11852
rect 2547 11849 2559 11883
rect 2501 11843 2559 11849
rect 2961 11883 3019 11889
rect 2961 11849 2973 11883
rect 3007 11880 3019 11883
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3007 11852 3801 11880
rect 3007 11849 3019 11852
rect 2961 11843 3019 11849
rect 3789 11849 3801 11852
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 4249 11883 4307 11889
rect 4249 11880 4261 11883
rect 4120 11852 4261 11880
rect 4120 11840 4126 11852
rect 4249 11849 4261 11852
rect 4295 11849 4307 11883
rect 4249 11843 4307 11849
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 5074 11880 5080 11892
rect 4488 11852 5080 11880
rect 4488 11840 4494 11852
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 6914 11880 6920 11892
rect 6875 11852 6920 11880
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 9493 11883 9551 11889
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 9766 11880 9772 11892
rect 9539 11852 9772 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 12069 11883 12127 11889
rect 12069 11849 12081 11883
rect 12115 11849 12127 11883
rect 12069 11843 12127 11849
rect 12529 11883 12587 11889
rect 12529 11849 12541 11883
rect 12575 11880 12587 11883
rect 17310 11880 17316 11892
rect 12575 11852 17316 11880
rect 12575 11849 12587 11852
rect 12529 11843 12587 11849
rect 2314 11812 2320 11824
rect 1964 11784 2320 11812
rect 1964 11685 1992 11784
rect 2314 11772 2320 11784
rect 2372 11772 2378 11824
rect 2869 11815 2927 11821
rect 2869 11781 2881 11815
rect 2915 11812 2927 11815
rect 3234 11812 3240 11824
rect 2915 11784 3240 11812
rect 2915 11781 2927 11784
rect 2869 11775 2927 11781
rect 3234 11772 3240 11784
rect 3292 11772 3298 11824
rect 4614 11812 4620 11824
rect 3436 11784 4620 11812
rect 3436 11744 3464 11784
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 4985 11815 5043 11821
rect 4985 11781 4997 11815
rect 5031 11812 5043 11815
rect 5350 11812 5356 11824
rect 5031 11784 5356 11812
rect 5031 11781 5043 11784
rect 4985 11775 5043 11781
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 5534 11772 5540 11824
rect 5592 11812 5598 11824
rect 10606 11815 10664 11821
rect 10606 11812 10618 11815
rect 5592 11784 10618 11812
rect 5592 11772 5598 11784
rect 10606 11781 10618 11784
rect 10652 11812 10664 11815
rect 10652 11784 10732 11812
rect 10652 11781 10664 11784
rect 10606 11775 10664 11781
rect 2792 11716 3464 11744
rect 4157 11747 4215 11753
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11645 2007 11679
rect 1949 11639 2007 11645
rect 2222 11636 2228 11688
rect 2280 11676 2286 11688
rect 2792 11676 2820 11716
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 5074 11744 5080 11756
rect 4203 11716 5080 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 5074 11704 5080 11716
rect 5132 11704 5138 11756
rect 7285 11747 7343 11753
rect 5184 11716 6868 11744
rect 2280 11648 2820 11676
rect 2280 11636 2286 11648
rect 2866 11636 2872 11688
rect 2924 11676 2930 11688
rect 3053 11679 3111 11685
rect 3053 11676 3065 11679
rect 2924 11648 3065 11676
rect 2924 11636 2930 11648
rect 3053 11645 3065 11648
rect 3099 11645 3111 11679
rect 3053 11639 3111 11645
rect 4433 11679 4491 11685
rect 4433 11645 4445 11679
rect 4479 11645 4491 11679
rect 4433 11639 4491 11645
rect 2406 11568 2412 11620
rect 2464 11608 2470 11620
rect 3878 11608 3884 11620
rect 2464 11580 3884 11608
rect 2464 11568 2470 11580
rect 3878 11568 3884 11580
rect 3936 11608 3942 11620
rect 4448 11608 4476 11639
rect 4614 11636 4620 11688
rect 4672 11676 4678 11688
rect 5184 11676 5212 11716
rect 4672 11648 5212 11676
rect 5353 11679 5411 11685
rect 4672 11636 4678 11648
rect 5353 11645 5365 11679
rect 5399 11676 5411 11679
rect 5442 11676 5448 11688
rect 5399 11648 5448 11676
rect 5399 11645 5411 11648
rect 5353 11639 5411 11645
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 6730 11676 6736 11688
rect 5767 11648 6736 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 5736 11608 5764 11639
rect 6730 11636 6736 11648
rect 6788 11636 6794 11688
rect 3936 11580 5764 11608
rect 6840 11608 6868 11716
rect 7285 11713 7297 11747
rect 7331 11744 7343 11747
rect 7834 11744 7840 11756
rect 7331 11716 7840 11744
rect 7331 11713 7343 11716
rect 7285 11707 7343 11713
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 10704 11744 10732 11784
rect 10870 11772 10876 11824
rect 10928 11812 10934 11824
rect 11609 11815 11667 11821
rect 11609 11812 11621 11815
rect 10928 11784 11621 11812
rect 10928 11772 10934 11784
rect 11609 11781 11621 11784
rect 11655 11812 11667 11815
rect 12084 11812 12112 11843
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 18046 11880 18052 11892
rect 18007 11852 18052 11880
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 18966 11840 18972 11892
rect 19024 11880 19030 11892
rect 19153 11883 19211 11889
rect 19153 11880 19165 11883
rect 19024 11852 19165 11880
rect 19024 11840 19030 11852
rect 19153 11849 19165 11852
rect 19199 11849 19211 11883
rect 19794 11880 19800 11892
rect 19755 11852 19800 11880
rect 19153 11843 19211 11849
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 20162 11880 20168 11892
rect 20123 11852 20168 11880
rect 20162 11840 20168 11852
rect 20220 11840 20226 11892
rect 20441 11883 20499 11889
rect 20441 11849 20453 11883
rect 20487 11880 20499 11883
rect 20806 11880 20812 11892
rect 20487 11852 20812 11880
rect 20487 11849 20499 11852
rect 20441 11843 20499 11849
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 11655 11784 12112 11812
rect 11655 11781 11667 11784
rect 11609 11775 11667 11781
rect 12158 11772 12164 11824
rect 12216 11812 12222 11824
rect 14378 11815 14436 11821
rect 14378 11812 14390 11815
rect 12216 11784 14390 11812
rect 12216 11772 12222 11784
rect 14378 11781 14390 11784
rect 14424 11781 14436 11815
rect 14378 11775 14436 11781
rect 15188 11815 15246 11821
rect 15188 11781 15200 11815
rect 15234 11812 15246 11815
rect 15838 11812 15844 11824
rect 15234 11784 15844 11812
rect 15234 11781 15246 11784
rect 15188 11775 15246 11781
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 17770 11812 17776 11824
rect 16684 11784 17776 11812
rect 16574 11744 16580 11756
rect 10704 11716 16580 11744
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16684 11753 16712 11784
rect 17770 11772 17776 11784
rect 17828 11772 17834 11824
rect 18230 11812 18236 11824
rect 17880 11784 18236 11812
rect 16669 11747 16727 11753
rect 16669 11713 16681 11747
rect 16715 11713 16727 11747
rect 16925 11747 16983 11753
rect 16925 11744 16937 11747
rect 16669 11707 16727 11713
rect 16776 11716 16937 11744
rect 7374 11676 7380 11688
rect 7335 11648 7380 11676
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 7561 11679 7619 11685
rect 7561 11676 7573 11679
rect 7524 11648 7573 11676
rect 7524 11636 7530 11648
rect 7561 11645 7573 11648
rect 7607 11676 7619 11679
rect 9030 11676 9036 11688
rect 7607 11648 9036 11676
rect 7607 11645 7619 11648
rect 7561 11639 7619 11645
rect 9030 11636 9036 11648
rect 9088 11636 9094 11688
rect 10870 11685 10876 11688
rect 10866 11639 10876 11685
rect 10928 11676 10934 11688
rect 12897 11679 12955 11685
rect 10928 11648 10966 11676
rect 10870 11636 10876 11639
rect 10928 11636 10934 11648
rect 12897 11645 12909 11679
rect 12943 11676 12955 11679
rect 13630 11676 13636 11688
rect 12943 11648 13636 11676
rect 12943 11645 12955 11648
rect 12897 11639 12955 11645
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 14645 11679 14703 11685
rect 14645 11645 14657 11679
rect 14691 11676 14703 11679
rect 14918 11676 14924 11688
rect 14691 11648 14924 11676
rect 14691 11645 14703 11648
rect 14645 11639 14703 11645
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 16776 11676 16804 11716
rect 16925 11713 16937 11716
rect 16971 11744 16983 11747
rect 17880 11744 17908 11784
rect 18230 11772 18236 11784
rect 18288 11812 18294 11824
rect 19705 11815 19763 11821
rect 18288 11784 19656 11812
rect 18288 11772 18294 11784
rect 16971 11716 17908 11744
rect 16971 11713 16983 11716
rect 16925 11707 16983 11713
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18969 11747 19027 11753
rect 18969 11744 18981 11747
rect 18012 11716 18981 11744
rect 18012 11704 18018 11716
rect 18969 11713 18981 11716
rect 19015 11713 19027 11747
rect 19628 11744 19656 11784
rect 19705 11781 19717 11815
rect 19751 11812 19763 11815
rect 20254 11812 20260 11824
rect 19751 11784 20260 11812
rect 19751 11781 19763 11784
rect 19705 11775 19763 11781
rect 20254 11772 20260 11784
rect 20312 11812 20318 11824
rect 20622 11812 20628 11824
rect 20312 11784 20628 11812
rect 20312 11772 20318 11784
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 20809 11747 20867 11753
rect 19628 11716 19748 11744
rect 18969 11707 19027 11713
rect 16684 11648 16804 11676
rect 19613 11679 19671 11685
rect 7929 11611 7987 11617
rect 7929 11608 7941 11611
rect 6840 11580 7941 11608
rect 3936 11568 3942 11580
rect 7929 11577 7941 11580
rect 7975 11577 7987 11611
rect 7929 11571 7987 11577
rect 8757 11611 8815 11617
rect 8757 11577 8769 11611
rect 8803 11608 8815 11611
rect 9858 11608 9864 11620
rect 8803 11580 9864 11608
rect 8803 11577 8815 11580
rect 8757 11571 8815 11577
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 13078 11608 13084 11620
rect 12406 11580 13084 11608
rect 6457 11543 6515 11549
rect 6457 11509 6469 11543
rect 6503 11540 6515 11543
rect 6822 11540 6828 11552
rect 6503 11512 6828 11540
rect 6503 11509 6515 11512
rect 6457 11503 6515 11509
rect 6822 11500 6828 11512
rect 6880 11540 6886 11552
rect 8110 11540 8116 11552
rect 6880 11512 8116 11540
rect 6880 11500 6886 11512
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 8294 11540 8300 11552
rect 8255 11512 8300 11540
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 9125 11543 9183 11549
rect 9125 11509 9137 11543
rect 9171 11540 9183 11543
rect 9490 11540 9496 11552
rect 9171 11512 9496 11540
rect 9171 11509 9183 11512
rect 9125 11503 9183 11509
rect 9490 11500 9496 11512
rect 9548 11540 9554 11552
rect 12406 11540 12434 11580
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 13262 11608 13268 11620
rect 13223 11580 13268 11608
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 16684 11608 16712 11648
rect 19613 11645 19625 11679
rect 19659 11645 19671 11679
rect 19720 11676 19748 11716
rect 20809 11713 20821 11747
rect 20855 11744 20867 11747
rect 21542 11744 21548 11756
rect 20855 11716 21548 11744
rect 20855 11713 20867 11716
rect 20809 11707 20867 11713
rect 21542 11704 21548 11716
rect 21600 11704 21606 11756
rect 20438 11676 20444 11688
rect 19720 11648 20444 11676
rect 19613 11639 19671 11645
rect 16132 11580 16712 11608
rect 9548 11512 12434 11540
rect 9548 11500 9554 11512
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 14826 11540 14832 11552
rect 14700 11512 14832 11540
rect 14700 11500 14706 11512
rect 14826 11500 14832 11512
rect 14884 11540 14890 11552
rect 16132 11540 16160 11580
rect 14884 11512 16160 11540
rect 14884 11500 14890 11512
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16301 11543 16359 11549
rect 16301 11540 16313 11543
rect 16264 11512 16313 11540
rect 16264 11500 16270 11512
rect 16301 11509 16313 11512
rect 16347 11509 16359 11543
rect 16301 11503 16359 11509
rect 16574 11500 16580 11552
rect 16632 11540 16638 11552
rect 17402 11540 17408 11552
rect 16632 11512 17408 11540
rect 16632 11500 16638 11512
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 17862 11500 17868 11552
rect 17920 11540 17926 11552
rect 18417 11543 18475 11549
rect 18417 11540 18429 11543
rect 17920 11512 18429 11540
rect 17920 11500 17926 11512
rect 18417 11509 18429 11512
rect 18463 11540 18475 11543
rect 19058 11540 19064 11552
rect 18463 11512 19064 11540
rect 18463 11509 18475 11512
rect 18417 11503 18475 11509
rect 19058 11500 19064 11512
rect 19116 11500 19122 11552
rect 19628 11540 19656 11639
rect 20438 11636 20444 11648
rect 20496 11636 20502 11688
rect 20714 11636 20720 11688
rect 20772 11676 20778 11688
rect 20898 11676 20904 11688
rect 20772 11648 20904 11676
rect 20772 11636 20778 11648
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 20993 11679 21051 11685
rect 20993 11645 21005 11679
rect 21039 11645 21051 11679
rect 20993 11639 21051 11645
rect 20530 11568 20536 11620
rect 20588 11608 20594 11620
rect 21008 11608 21036 11639
rect 20588 11580 21036 11608
rect 20588 11568 20594 11580
rect 21174 11540 21180 11552
rect 19628 11512 21180 11540
rect 21174 11500 21180 11512
rect 21232 11500 21238 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 1946 11336 1952 11348
rect 1627 11308 1952 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1946 11296 1952 11308
rect 2004 11296 2010 11348
rect 3326 11336 3332 11348
rect 3287 11308 3332 11336
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 3970 11336 3976 11348
rect 3931 11308 3976 11336
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4212 11308 4537 11336
rect 4212 11296 4218 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 6822 11336 6828 11348
rect 4525 11299 4583 11305
rect 4632 11308 6828 11336
rect 4632 11268 4660 11308
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 8478 11336 8484 11348
rect 7668 11308 8484 11336
rect 2792 11240 4660 11268
rect 5092 11240 5672 11268
rect 2792 11209 2820 11240
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11169 2283 11203
rect 2225 11163 2283 11169
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11169 2835 11203
rect 2777 11163 2835 11169
rect 1670 11092 1676 11144
rect 1728 11132 1734 11144
rect 2240 11132 2268 11163
rect 2866 11160 2872 11212
rect 2924 11160 2930 11212
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 5092 11200 5120 11240
rect 4396 11172 5120 11200
rect 5169 11203 5227 11209
rect 4396 11160 4402 11172
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 5258 11200 5264 11212
rect 5215 11172 5264 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 5644 11200 5672 11240
rect 5718 11228 5724 11280
rect 5776 11268 5782 11280
rect 7101 11271 7159 11277
rect 7101 11268 7113 11271
rect 5776 11240 7113 11268
rect 5776 11228 5782 11240
rect 7101 11237 7113 11240
rect 7147 11237 7159 11271
rect 7101 11231 7159 11237
rect 7668 11209 7696 11308
rect 8478 11296 8484 11308
rect 8536 11336 8542 11348
rect 10410 11336 10416 11348
rect 8536 11308 10416 11336
rect 8536 11296 8542 11308
rect 10410 11296 10416 11308
rect 10468 11296 10474 11348
rect 10870 11336 10876 11348
rect 10831 11308 10876 11336
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 11241 11339 11299 11345
rect 11241 11305 11253 11339
rect 11287 11336 11299 11339
rect 11882 11336 11888 11348
rect 11287 11308 11888 11336
rect 11287 11305 11299 11308
rect 11241 11299 11299 11305
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 17034 11336 17040 11348
rect 12124 11308 17040 11336
rect 12124 11296 12130 11308
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 17586 11336 17592 11348
rect 17547 11308 17592 11336
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 18782 11336 18788 11348
rect 17788 11308 18788 11336
rect 10505 11271 10563 11277
rect 10505 11237 10517 11271
rect 10551 11237 10563 11271
rect 10505 11231 10563 11237
rect 13081 11271 13139 11277
rect 13081 11237 13093 11271
rect 13127 11268 13139 11271
rect 13814 11268 13820 11280
rect 13127 11240 13820 11268
rect 13127 11237 13139 11240
rect 13081 11231 13139 11237
rect 6181 11203 6239 11209
rect 6181 11200 6193 11203
rect 5644 11172 6193 11200
rect 6181 11169 6193 11172
rect 6227 11200 6239 11203
rect 7653 11203 7711 11209
rect 7653 11200 7665 11203
rect 6227 11172 7665 11200
rect 6227 11169 6239 11172
rect 6181 11163 6239 11169
rect 7653 11169 7665 11172
rect 7699 11169 7711 11203
rect 9122 11200 9128 11212
rect 9083 11172 9128 11200
rect 7653 11163 7711 11169
rect 9122 11160 9128 11172
rect 9180 11160 9186 11212
rect 2884 11132 2912 11160
rect 1728 11104 2176 11132
rect 2240 11104 2912 11132
rect 1728 11092 1734 11104
rect 2038 11064 2044 11076
rect 1999 11036 2044 11064
rect 2038 11024 2044 11036
rect 2096 11024 2102 11076
rect 2148 11064 2176 11104
rect 3326 11092 3332 11144
rect 3384 11132 3390 11144
rect 6089 11135 6147 11141
rect 6089 11132 6101 11135
rect 3384 11104 6101 11132
rect 3384 11092 3390 11104
rect 6089 11101 6101 11104
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7524 11104 7573 11132
rect 7524 11092 7530 11104
rect 7561 11101 7573 11104
rect 7607 11132 7619 11135
rect 8202 11132 8208 11144
rect 7607 11104 8208 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9381 11135 9439 11141
rect 9381 11132 9393 11135
rect 9272 11104 9393 11132
rect 9272 11092 9278 11104
rect 9381 11101 9393 11104
rect 9427 11101 9439 11135
rect 10520 11132 10548 11231
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 16117 11271 16175 11277
rect 16117 11237 16129 11271
rect 16163 11268 16175 11271
rect 17788 11268 17816 11308
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 19337 11339 19395 11345
rect 19337 11305 19349 11339
rect 19383 11336 19395 11339
rect 19978 11336 19984 11348
rect 19383 11308 19984 11336
rect 19383 11305 19395 11308
rect 19337 11299 19395 11305
rect 19978 11296 19984 11308
rect 20036 11296 20042 11348
rect 21177 11339 21235 11345
rect 21177 11305 21189 11339
rect 21223 11336 21235 11339
rect 22094 11336 22100 11348
rect 21223 11308 22100 11336
rect 21223 11305 21235 11308
rect 21177 11299 21235 11305
rect 22094 11296 22100 11308
rect 22152 11296 22158 11348
rect 17954 11268 17960 11280
rect 16163 11240 17816 11268
rect 17915 11240 17960 11268
rect 16163 11237 16175 11240
rect 16117 11231 16175 11237
rect 17954 11228 17960 11240
rect 18012 11228 18018 11280
rect 18230 11228 18236 11280
rect 18288 11268 18294 11280
rect 18325 11271 18383 11277
rect 18325 11268 18337 11271
rect 18288 11240 18337 11268
rect 18288 11228 18294 11240
rect 18325 11237 18337 11240
rect 18371 11237 18383 11271
rect 18325 11231 18383 11237
rect 18877 11271 18935 11277
rect 18877 11237 18889 11271
rect 18923 11268 18935 11271
rect 19518 11268 19524 11280
rect 18923 11240 19524 11268
rect 18923 11237 18935 11240
rect 18877 11231 18935 11237
rect 19518 11228 19524 11240
rect 19576 11228 19582 11280
rect 10870 11160 10876 11212
rect 10928 11200 10934 11212
rect 11701 11203 11759 11209
rect 11701 11200 11713 11203
rect 10928 11172 11713 11200
rect 10928 11160 10934 11172
rect 11701 11169 11713 11172
rect 11747 11169 11759 11203
rect 11701 11163 11759 11169
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11200 14519 11203
rect 19242 11200 19248 11212
rect 14507 11172 19248 11200
rect 14507 11169 14519 11172
rect 14461 11163 14519 11169
rect 11238 11132 11244 11144
rect 10520 11104 11244 11132
rect 9381 11095 9439 11101
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 11716 11132 11744 11163
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 20717 11203 20775 11209
rect 20717 11169 20729 11203
rect 20763 11200 20775 11203
rect 20990 11200 20996 11212
rect 20763 11172 20996 11200
rect 20763 11169 20775 11172
rect 20717 11163 20775 11169
rect 13357 11135 13415 11141
rect 13357 11132 13369 11135
rect 11716 11104 13369 11132
rect 13357 11101 13369 11104
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 16945 11135 17003 11141
rect 16945 11101 16957 11135
rect 16991 11132 17003 11135
rect 18690 11132 18696 11144
rect 16991 11104 18696 11132
rect 16991 11101 17003 11104
rect 16945 11095 17003 11101
rect 18690 11092 18696 11104
rect 18748 11092 18754 11144
rect 19150 11092 19156 11144
rect 19208 11132 19214 11144
rect 20732 11132 20760 11163
rect 20990 11160 20996 11172
rect 21048 11160 21054 11212
rect 19208 11104 20760 11132
rect 19208 11092 19214 11104
rect 2869 11067 2927 11073
rect 2869 11064 2881 11067
rect 2148 11036 2881 11064
rect 2869 11033 2881 11036
rect 2915 11033 2927 11067
rect 3878 11064 3884 11076
rect 3839 11036 3884 11064
rect 2869 11027 2927 11033
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4890 11064 4896 11076
rect 4172 11036 4896 11064
rect 4172 11008 4200 11036
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 4985 11067 5043 11073
rect 4985 11033 4997 11067
rect 5031 11033 5043 11067
rect 4985 11027 5043 11033
rect 5997 11067 6055 11073
rect 5997 11033 6009 11067
rect 6043 11064 6055 11067
rect 6641 11067 6699 11073
rect 6641 11064 6653 11067
rect 6043 11036 6653 11064
rect 6043 11033 6055 11036
rect 5997 11027 6055 11033
rect 6641 11033 6653 11036
rect 6687 11033 6699 11067
rect 6641 11027 6699 11033
rect 1946 10996 1952 11008
rect 1907 10968 1952 10996
rect 1946 10956 1952 10968
rect 2004 10956 2010 11008
rect 2958 10996 2964 11008
rect 2919 10968 2964 10996
rect 2958 10956 2964 10968
rect 3016 10956 3022 11008
rect 4154 10956 4160 11008
rect 4212 10956 4218 11008
rect 4430 10956 4436 11008
rect 4488 10996 4494 11008
rect 5000 10996 5028 11027
rect 6914 11024 6920 11076
rect 6972 11064 6978 11076
rect 8113 11067 8171 11073
rect 8113 11064 8125 11067
rect 6972 11036 8125 11064
rect 6972 11024 6978 11036
rect 8113 11033 8125 11036
rect 8159 11033 8171 11067
rect 8113 11027 8171 11033
rect 9582 11024 9588 11076
rect 9640 11064 9646 11076
rect 20530 11073 20536 11076
rect 11946 11067 12004 11073
rect 11946 11064 11958 11067
rect 9640 11036 11958 11064
rect 9640 11024 9646 11036
rect 11946 11033 11958 11036
rect 11992 11033 12004 11067
rect 11946 11027 12004 11033
rect 15289 11067 15347 11073
rect 15289 11033 15301 11067
rect 15335 11064 15347 11067
rect 20472 11067 20536 11073
rect 15335 11036 20392 11064
rect 15335 11033 15347 11036
rect 15289 11027 15347 11033
rect 5074 10996 5080 11008
rect 4488 10968 5080 10996
rect 4488 10956 4494 10968
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 5626 10996 5632 11008
rect 5587 10968 5632 10996
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 7098 10956 7104 11008
rect 7156 10996 7162 11008
rect 7469 10999 7527 11005
rect 7469 10996 7481 10999
rect 7156 10968 7481 10996
rect 7156 10956 7162 10968
rect 7469 10965 7481 10968
rect 7515 10965 7527 10999
rect 8478 10996 8484 11008
rect 8439 10968 8484 10996
rect 7469 10959 7527 10965
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 12066 10996 12072 11008
rect 10284 10968 12072 10996
rect 10284 10956 10290 10968
rect 12066 10956 12072 10968
rect 12124 10956 12130 11008
rect 14829 10999 14887 11005
rect 14829 10965 14841 10999
rect 14875 10996 14887 10999
rect 14918 10996 14924 11008
rect 14875 10968 14924 10996
rect 14875 10965 14887 10968
rect 14829 10959 14887 10965
rect 14918 10956 14924 10968
rect 14976 10996 14982 11008
rect 15749 10999 15807 11005
rect 15749 10996 15761 10999
rect 14976 10968 15761 10996
rect 14976 10956 14982 10968
rect 15749 10965 15761 10968
rect 15795 10996 15807 10999
rect 16485 10999 16543 11005
rect 16485 10996 16497 10999
rect 15795 10968 16497 10996
rect 15795 10965 15807 10968
rect 15749 10959 15807 10965
rect 16485 10965 16497 10968
rect 16531 10965 16543 10999
rect 16485 10959 16543 10965
rect 17034 10956 17040 11008
rect 17092 10996 17098 11008
rect 17221 10999 17279 11005
rect 17221 10996 17233 10999
rect 17092 10968 17233 10996
rect 17092 10956 17098 10968
rect 17221 10965 17233 10968
rect 17267 10965 17279 10999
rect 20364 10996 20392 11036
rect 20472 11033 20484 11067
rect 20518 11033 20536 11067
rect 20472 11027 20536 11033
rect 20530 11024 20536 11027
rect 20588 11024 20594 11076
rect 21266 11064 21272 11076
rect 20640 11036 21272 11064
rect 20640 10996 20668 11036
rect 21266 11024 21272 11036
rect 21324 11024 21330 11076
rect 20364 10968 20668 10996
rect 17221 10959 17279 10965
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 1394 10752 1400 10804
rect 1452 10792 1458 10804
rect 2869 10795 2927 10801
rect 2869 10792 2881 10795
rect 1452 10764 2881 10792
rect 1452 10752 1458 10764
rect 2869 10761 2881 10764
rect 2915 10792 2927 10795
rect 4062 10792 4068 10804
rect 2915 10764 4068 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4617 10795 4675 10801
rect 4617 10761 4629 10795
rect 4663 10792 4675 10795
rect 5442 10792 5448 10804
rect 4663 10764 5448 10792
rect 4663 10761 4675 10764
rect 4617 10755 4675 10761
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5994 10752 6000 10804
rect 6052 10792 6058 10804
rect 6270 10792 6276 10804
rect 6052 10764 6276 10792
rect 6052 10752 6058 10764
rect 6270 10752 6276 10764
rect 6328 10792 6334 10804
rect 7745 10795 7803 10801
rect 7745 10792 7757 10795
rect 6328 10764 7757 10792
rect 6328 10752 6334 10764
rect 7745 10761 7757 10764
rect 7791 10792 7803 10795
rect 10870 10792 10876 10804
rect 7791 10764 10732 10792
rect 10831 10764 10876 10792
rect 7791 10761 7803 10764
rect 7745 10755 7803 10761
rect 3142 10684 3148 10736
rect 3200 10724 3206 10736
rect 3513 10727 3571 10733
rect 3513 10724 3525 10727
rect 3200 10696 3525 10724
rect 3200 10684 3206 10696
rect 3513 10693 3525 10696
rect 3559 10693 3571 10727
rect 3513 10687 3571 10693
rect 3878 10684 3884 10736
rect 3936 10724 3942 10736
rect 6365 10727 6423 10733
rect 6365 10724 6377 10727
rect 3936 10696 6377 10724
rect 3936 10684 3942 10696
rect 6365 10693 6377 10696
rect 6411 10693 6423 10727
rect 6365 10687 6423 10693
rect 6454 10684 6460 10736
rect 6512 10724 6518 10736
rect 6638 10724 6644 10736
rect 6512 10696 6644 10724
rect 6512 10684 6518 10696
rect 6638 10684 6644 10696
rect 6696 10684 6702 10736
rect 7282 10684 7288 10736
rect 7340 10724 7346 10736
rect 7377 10727 7435 10733
rect 7377 10724 7389 10727
rect 7340 10696 7389 10724
rect 7340 10684 7346 10696
rect 7377 10693 7389 10696
rect 7423 10724 7435 10727
rect 7466 10724 7472 10736
rect 7423 10696 7472 10724
rect 7423 10693 7435 10696
rect 7377 10687 7435 10693
rect 7466 10684 7472 10696
rect 7524 10684 7530 10736
rect 8113 10727 8171 10733
rect 8113 10693 8125 10727
rect 8159 10724 8171 10727
rect 8294 10724 8300 10736
rect 8159 10696 8300 10724
rect 8159 10693 8171 10696
rect 8113 10687 8171 10693
rect 8294 10684 8300 10696
rect 8352 10724 8358 10736
rect 10134 10724 10140 10736
rect 8352 10696 10140 10724
rect 8352 10684 8358 10696
rect 10134 10684 10140 10696
rect 10192 10684 10198 10736
rect 10260 10727 10318 10733
rect 10260 10693 10272 10727
rect 10306 10724 10318 10727
rect 10594 10724 10600 10736
rect 10306 10696 10600 10724
rect 10306 10693 10318 10696
rect 10260 10687 10318 10693
rect 10594 10684 10600 10696
rect 10652 10684 10658 10736
rect 10704 10724 10732 10764
rect 10870 10752 10876 10764
rect 10928 10792 10934 10804
rect 11977 10795 12035 10801
rect 11977 10792 11989 10795
rect 10928 10764 11989 10792
rect 10928 10752 10934 10764
rect 11977 10761 11989 10764
rect 12023 10761 12035 10795
rect 14366 10792 14372 10804
rect 11977 10755 12035 10761
rect 14292 10764 14372 10792
rect 11054 10724 11060 10736
rect 10704 10696 11060 10724
rect 11054 10684 11060 10696
rect 11112 10684 11118 10736
rect 13814 10724 13820 10736
rect 12406 10696 13820 10724
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1636 10628 1961 10656
rect 1636 10616 1642 10628
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 5534 10656 5540 10668
rect 1949 10619 2007 10625
rect 4448 10628 5540 10656
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10588 2283 10591
rect 2958 10588 2964 10600
rect 2271 10560 2774 10588
rect 2919 10560 2964 10588
rect 2271 10557 2283 10560
rect 2225 10551 2283 10557
rect 2746 10532 2774 10560
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 4448 10597 4476 10628
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 5813 10659 5871 10665
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 5994 10656 6000 10668
rect 5859 10628 6000 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 8018 10616 8024 10668
rect 8076 10656 8082 10668
rect 8757 10659 8815 10665
rect 8757 10656 8769 10659
rect 8076 10628 8769 10656
rect 8076 10616 8082 10628
rect 8757 10625 8769 10628
rect 8803 10656 8815 10659
rect 9858 10656 9864 10668
rect 8803 10628 9864 10656
rect 8803 10625 8815 10628
rect 8757 10619 8815 10625
rect 9858 10616 9864 10628
rect 9916 10656 9922 10668
rect 10505 10659 10563 10665
rect 9916 10628 10465 10656
rect 9916 10616 9922 10628
rect 4433 10591 4491 10597
rect 3108 10560 3153 10588
rect 3108 10548 3114 10560
rect 4433 10557 4445 10591
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10588 4583 10591
rect 4890 10588 4896 10600
rect 4571 10560 4896 10588
rect 4571 10557 4583 10560
rect 4525 10551 4583 10557
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 5258 10548 5264 10600
rect 5316 10588 5322 10600
rect 5445 10591 5503 10597
rect 5445 10588 5457 10591
rect 5316 10560 5457 10588
rect 5316 10548 5322 10560
rect 5445 10557 5457 10560
rect 5491 10588 5503 10591
rect 10437 10588 10465 10628
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 10870 10656 10876 10668
rect 10551 10628 10876 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 10870 10616 10876 10628
rect 10928 10616 10934 10668
rect 10778 10588 10784 10600
rect 5491 10560 9260 10588
rect 10437 10560 10784 10588
rect 5491 10557 5503 10560
rect 5445 10551 5503 10557
rect 2746 10492 2780 10532
rect 2774 10480 2780 10492
rect 2832 10520 2838 10532
rect 8478 10520 8484 10532
rect 2832 10492 8484 10520
rect 2832 10480 2838 10492
rect 8478 10480 8484 10492
rect 8536 10480 8542 10532
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 2501 10455 2559 10461
rect 2501 10452 2513 10455
rect 2188 10424 2513 10452
rect 2188 10412 2194 10424
rect 2501 10421 2513 10424
rect 2547 10421 2559 10455
rect 2501 10415 2559 10421
rect 4985 10455 5043 10461
rect 4985 10421 4997 10455
rect 5031 10452 5043 10455
rect 5166 10452 5172 10464
rect 5031 10424 5172 10452
rect 5031 10421 5043 10424
rect 4985 10415 5043 10421
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 7009 10455 7067 10461
rect 7009 10421 7021 10455
rect 7055 10452 7067 10455
rect 7098 10452 7104 10464
rect 7055 10424 7104 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 9122 10452 9128 10464
rect 9083 10424 9128 10452
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9232 10452 9260 10560
rect 10778 10548 10784 10560
rect 10836 10588 10842 10600
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 10836 10560 11621 10588
rect 10836 10548 10842 10560
rect 11609 10557 11621 10560
rect 11655 10557 11667 10591
rect 11609 10551 11667 10557
rect 12406 10520 12434 10696
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 14292 10733 14320 10764
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 17402 10792 17408 10804
rect 17363 10764 17408 10792
rect 17402 10752 17408 10764
rect 17460 10752 17466 10804
rect 18598 10752 18604 10804
rect 18656 10792 18662 10804
rect 20530 10792 20536 10804
rect 18656 10764 19748 10792
rect 20491 10764 20536 10792
rect 18656 10752 18662 10764
rect 14286 10727 14344 10733
rect 14286 10693 14298 10727
rect 14332 10693 14344 10727
rect 14286 10687 14344 10693
rect 14550 10684 14556 10736
rect 14608 10724 14614 10736
rect 15010 10724 15016 10736
rect 14608 10696 15016 10724
rect 14608 10684 14614 10696
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 17034 10684 17040 10736
rect 17092 10724 17098 10736
rect 18518 10727 18576 10733
rect 18518 10724 18530 10727
rect 17092 10696 18530 10724
rect 17092 10684 17098 10696
rect 18518 10693 18530 10696
rect 18564 10693 18576 10727
rect 18518 10687 18576 10693
rect 19420 10727 19478 10733
rect 19420 10693 19432 10727
rect 19466 10724 19478 10727
rect 19610 10724 19616 10736
rect 19466 10696 19616 10724
rect 19466 10693 19478 10696
rect 19420 10687 19478 10693
rect 19610 10684 19616 10696
rect 19668 10684 19674 10736
rect 19720 10724 19748 10764
rect 20530 10752 20536 10764
rect 20588 10752 20594 10804
rect 21085 10727 21143 10733
rect 21085 10724 21097 10727
rect 19720 10696 21097 10724
rect 21085 10693 21097 10696
rect 21131 10693 21143 10727
rect 21085 10687 21143 10693
rect 12805 10659 12863 10665
rect 12805 10625 12817 10659
rect 12851 10656 12863 10659
rect 18230 10656 18236 10668
rect 12851 10628 18236 10656
rect 12851 10625 12863 10628
rect 12805 10619 12863 10625
rect 18230 10616 18236 10628
rect 18288 10616 18294 10668
rect 18785 10659 18843 10665
rect 18785 10625 18797 10659
rect 18831 10656 18843 10659
rect 19150 10656 19156 10668
rect 18831 10628 19156 10656
rect 18831 10625 18843 10628
rect 18785 10619 18843 10625
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 19242 10616 19248 10668
rect 19300 10656 19306 10668
rect 21266 10656 21272 10668
rect 19300 10628 21272 10656
rect 19300 10616 19306 10628
rect 21266 10616 21272 10628
rect 21324 10616 21330 10668
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10588 14611 10591
rect 14599 10560 14964 10588
rect 14599 10557 14611 10560
rect 14553 10551 14611 10557
rect 13170 10520 13176 10532
rect 10520 10492 12434 10520
rect 13131 10492 13176 10520
rect 10520 10452 10548 10492
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 14936 10464 14964 10560
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 16298 10588 16304 10600
rect 15896 10560 16304 10588
rect 15896 10548 15902 10560
rect 16298 10548 16304 10560
rect 16356 10588 16362 10600
rect 17037 10591 17095 10597
rect 17037 10588 17049 10591
rect 16356 10560 17049 10588
rect 16356 10548 16362 10560
rect 17037 10557 17049 10560
rect 17083 10557 17095 10591
rect 17037 10551 17095 10557
rect 9232 10424 10548 10452
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 14918 10452 14924 10464
rect 12492 10424 12537 10452
rect 14879 10424 14924 10452
rect 12492 10412 12498 10424
rect 14918 10412 14924 10424
rect 14976 10452 14982 10464
rect 15473 10455 15531 10461
rect 15473 10452 15485 10455
rect 14976 10424 15485 10452
rect 14976 10412 14982 10424
rect 15473 10421 15485 10424
rect 15519 10452 15531 10455
rect 15841 10455 15899 10461
rect 15841 10452 15853 10455
rect 15519 10424 15853 10452
rect 15519 10421 15531 10424
rect 15473 10415 15531 10421
rect 15841 10421 15853 10424
rect 15887 10452 15899 10455
rect 16209 10455 16267 10461
rect 16209 10452 16221 10455
rect 15887 10424 16221 10452
rect 15887 10421 15899 10424
rect 15841 10415 15899 10421
rect 16209 10421 16221 10424
rect 16255 10452 16267 10455
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 16255 10424 16681 10452
rect 16255 10421 16267 10424
rect 16209 10415 16267 10421
rect 16669 10421 16681 10424
rect 16715 10421 16727 10455
rect 16669 10415 16727 10421
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1673 10251 1731 10257
rect 1673 10217 1685 10251
rect 1719 10248 1731 10251
rect 1946 10248 1952 10260
rect 1719 10220 1952 10248
rect 1719 10217 1731 10220
rect 1673 10211 1731 10217
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 3418 10248 3424 10260
rect 3379 10220 3424 10248
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 4890 10248 4896 10260
rect 4851 10220 4896 10248
rect 4890 10208 4896 10220
rect 4948 10208 4954 10260
rect 6273 10251 6331 10257
rect 6273 10217 6285 10251
rect 6319 10248 6331 10251
rect 6546 10248 6552 10260
rect 6319 10220 6552 10248
rect 6319 10217 6331 10220
rect 6273 10211 6331 10217
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 6730 10208 6736 10260
rect 6788 10248 6794 10260
rect 7282 10248 7288 10260
rect 6788 10220 7288 10248
rect 6788 10208 6794 10220
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 8941 10251 8999 10257
rect 8941 10217 8953 10251
rect 8987 10248 8999 10251
rect 9214 10248 9220 10260
rect 8987 10220 9220 10248
rect 8987 10217 8999 10220
rect 8941 10211 8999 10217
rect 9214 10208 9220 10220
rect 9272 10208 9278 10260
rect 10689 10251 10747 10257
rect 10689 10217 10701 10251
rect 10735 10248 10747 10251
rect 10870 10248 10876 10260
rect 10735 10220 10876 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 1578 10140 1584 10192
rect 1636 10180 1642 10192
rect 2961 10183 3019 10189
rect 1636 10152 2360 10180
rect 1636 10140 1642 10152
rect 2130 10112 2136 10124
rect 2091 10084 2136 10112
rect 2130 10072 2136 10084
rect 2188 10072 2194 10124
rect 2332 10121 2360 10152
rect 2961 10149 2973 10183
rect 3007 10180 3019 10183
rect 5350 10180 5356 10192
rect 3007 10152 5356 10180
rect 3007 10149 3019 10152
rect 2961 10143 3019 10149
rect 5350 10140 5356 10152
rect 5408 10140 5414 10192
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 5592 10152 5948 10180
rect 5592 10140 5598 10152
rect 2317 10115 2375 10121
rect 2317 10081 2329 10115
rect 2363 10112 2375 10115
rect 2406 10112 2412 10124
rect 2363 10084 2412 10112
rect 2363 10081 2375 10084
rect 2317 10075 2375 10081
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 3418 10072 3424 10124
rect 3476 10112 3482 10124
rect 4154 10112 4160 10124
rect 3476 10084 4160 10112
rect 3476 10072 3482 10084
rect 4154 10072 4160 10084
rect 4212 10072 4218 10124
rect 4338 10112 4344 10124
rect 4299 10084 4344 10112
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 5718 10112 5724 10124
rect 5679 10084 5724 10112
rect 5718 10072 5724 10084
rect 5776 10072 5782 10124
rect 5920 10121 5948 10152
rect 7466 10140 7472 10192
rect 7524 10180 7530 10192
rect 8573 10183 8631 10189
rect 7524 10152 8156 10180
rect 7524 10140 7530 10152
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10081 5963 10115
rect 6822 10112 6828 10124
rect 6783 10084 6828 10112
rect 5905 10075 5963 10081
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10044 2099 10047
rect 3142 10044 3148 10056
rect 2087 10016 3148 10044
rect 2087 10013 2099 10016
rect 2041 10007 2099 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3234 10004 3240 10056
rect 3292 10044 3298 10056
rect 3970 10044 3976 10056
rect 3292 10016 3976 10044
rect 3292 10004 3298 10016
rect 3970 10004 3976 10016
rect 4028 10004 4034 10056
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10044 4491 10047
rect 5442 10044 5448 10056
rect 4479 10016 5448 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5626 10044 5632 10056
rect 5587 10016 5632 10044
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 5920 10044 5948 10075
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 8018 10112 8024 10124
rect 7979 10084 8024 10112
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8128 10121 8156 10152
rect 8573 10149 8585 10183
rect 8619 10149 8631 10183
rect 8573 10143 8631 10149
rect 8113 10115 8171 10121
rect 8113 10081 8125 10115
rect 8159 10081 8171 10115
rect 8113 10075 8171 10081
rect 8478 10044 8484 10056
rect 5920 10016 8484 10044
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8588 10044 8616 10143
rect 10321 10115 10379 10121
rect 10321 10081 10333 10115
rect 10367 10112 10379 10115
rect 10704 10112 10732 10211
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 11517 10251 11575 10257
rect 11517 10217 11529 10251
rect 11563 10248 11575 10251
rect 11563 10220 13768 10248
rect 11563 10217 11575 10220
rect 11517 10211 11575 10217
rect 11977 10183 12035 10189
rect 11977 10149 11989 10183
rect 12023 10180 12035 10183
rect 13740 10180 13768 10220
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14274 10248 14280 10260
rect 13872 10220 14280 10248
rect 13872 10208 13878 10220
rect 14274 10208 14280 10220
rect 14332 10248 14338 10260
rect 14826 10248 14832 10260
rect 14332 10220 14832 10248
rect 14332 10208 14338 10220
rect 14826 10208 14832 10220
rect 14884 10208 14890 10260
rect 16853 10251 16911 10257
rect 15212 10220 16528 10248
rect 15212 10180 15240 10220
rect 12023 10152 12664 10180
rect 13740 10152 15240 10180
rect 12023 10149 12035 10152
rect 11977 10143 12035 10149
rect 10367 10084 10732 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 11238 10044 11244 10056
rect 8588 10016 11244 10044
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 11790 10044 11796 10056
rect 11751 10016 11796 10044
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12636 10044 12664 10152
rect 14366 10112 14372 10124
rect 13556 10084 14372 10112
rect 13556 10044 13584 10084
rect 14366 10072 14372 10084
rect 14424 10072 14430 10124
rect 16500 10112 16528 10220
rect 16853 10217 16865 10251
rect 16899 10248 16911 10251
rect 17126 10248 17132 10260
rect 16899 10220 17132 10248
rect 16899 10217 16911 10220
rect 16853 10211 16911 10217
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 17862 10248 17868 10260
rect 17328 10220 17868 10248
rect 16577 10183 16635 10189
rect 16577 10149 16589 10183
rect 16623 10180 16635 10183
rect 16942 10180 16948 10192
rect 16623 10152 16948 10180
rect 16623 10149 16635 10152
rect 16577 10143 16635 10149
rect 16942 10140 16948 10152
rect 17000 10180 17006 10192
rect 17328 10180 17356 10220
rect 17862 10208 17868 10220
rect 17920 10208 17926 10260
rect 18230 10208 18236 10260
rect 18288 10208 18294 10260
rect 18506 10208 18512 10260
rect 18564 10248 18570 10260
rect 18564 10220 20852 10248
rect 18564 10208 18570 10220
rect 17000 10152 17356 10180
rect 18248 10180 18276 10208
rect 18248 10152 20576 10180
rect 17000 10140 17006 10152
rect 20548 10124 20576 10152
rect 17218 10112 17224 10124
rect 16500 10084 17224 10112
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 18233 10115 18291 10121
rect 18233 10081 18245 10115
rect 18279 10112 18291 10115
rect 19058 10112 19064 10124
rect 18279 10084 19064 10112
rect 18279 10081 18291 10084
rect 18233 10075 18291 10081
rect 19058 10072 19064 10084
rect 19116 10072 19122 10124
rect 19978 10112 19984 10124
rect 19939 10084 19984 10112
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 20530 10112 20536 10124
rect 20443 10084 20536 10112
rect 20530 10072 20536 10084
rect 20588 10072 20594 10124
rect 20824 10121 20852 10220
rect 20809 10115 20867 10121
rect 20809 10081 20821 10115
rect 20855 10081 20867 10115
rect 20809 10075 20867 10081
rect 12636 10016 13584 10044
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10044 13691 10047
rect 13814 10044 13820 10056
rect 13679 10016 13820 10044
rect 13679 10013 13691 10016
rect 13633 10007 13691 10013
rect 13814 10004 13820 10016
rect 13872 10044 13878 10056
rect 14918 10044 14924 10056
rect 13872 10016 14924 10044
rect 13872 10004 13878 10016
rect 14918 10004 14924 10016
rect 14976 10044 14982 10056
rect 15197 10047 15255 10053
rect 15197 10044 15209 10047
rect 14976 10016 15209 10044
rect 14976 10004 14982 10016
rect 15197 10013 15209 10016
rect 15243 10013 15255 10047
rect 19705 10047 19763 10053
rect 15197 10007 15255 10013
rect 15396 10016 19012 10044
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 5902 9976 5908 9988
rect 2832 9948 5908 9976
rect 2832 9936 2838 9948
rect 5902 9936 5908 9948
rect 5960 9936 5966 9988
rect 6270 9936 6276 9988
rect 6328 9976 6334 9988
rect 6641 9979 6699 9985
rect 6641 9976 6653 9979
rect 6328 9948 6653 9976
rect 6328 9936 6334 9948
rect 6641 9945 6653 9948
rect 6687 9945 6699 9979
rect 7466 9976 7472 9988
rect 7427 9948 7472 9976
rect 6641 9939 6699 9945
rect 7466 9936 7472 9948
rect 7524 9976 7530 9988
rect 8202 9976 8208 9988
rect 7524 9948 8208 9976
rect 7524 9936 7530 9948
rect 8202 9936 8208 9948
rect 8260 9936 8266 9988
rect 10042 9936 10048 9988
rect 10100 9985 10106 9988
rect 10100 9976 10112 9985
rect 11149 9979 11207 9985
rect 10100 9948 10145 9976
rect 10100 9939 10112 9948
rect 11149 9945 11161 9979
rect 11195 9976 11207 9979
rect 11195 9948 12388 9976
rect 11195 9945 11207 9948
rect 11149 9939 11207 9945
rect 10100 9936 10106 9939
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 2924 9880 3893 9908
rect 2924 9868 2930 9880
rect 3881 9877 3893 9880
rect 3927 9908 3939 9911
rect 4154 9908 4160 9920
rect 3927 9880 4160 9908
rect 3927 9877 3939 9880
rect 3881 9871 3939 9877
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 4246 9868 4252 9920
rect 4304 9908 4310 9920
rect 4525 9911 4583 9917
rect 4525 9908 4537 9911
rect 4304 9880 4537 9908
rect 4304 9868 4310 9880
rect 4525 9877 4537 9880
rect 4571 9908 4583 9911
rect 4890 9908 4896 9920
rect 4571 9880 4896 9908
rect 4571 9877 4583 9880
rect 4525 9871 4583 9877
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 5258 9908 5264 9920
rect 5219 9880 5264 9908
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 6733 9911 6791 9917
rect 6733 9877 6745 9911
rect 6779 9908 6791 9911
rect 8294 9908 8300 9920
rect 6779 9880 8300 9908
rect 6779 9877 6791 9880
rect 6733 9871 6791 9877
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 11698 9868 11704 9920
rect 11756 9908 11762 9920
rect 11974 9908 11980 9920
rect 11756 9880 11980 9908
rect 11756 9868 11762 9880
rect 11974 9868 11980 9880
rect 12032 9908 12038 9920
rect 12253 9911 12311 9917
rect 12253 9908 12265 9911
rect 12032 9880 12265 9908
rect 12032 9868 12038 9880
rect 12253 9877 12265 9880
rect 12299 9877 12311 9911
rect 12360 9908 12388 9948
rect 13262 9936 13268 9988
rect 13320 9976 13326 9988
rect 13366 9979 13424 9985
rect 13366 9976 13378 9979
rect 13320 9948 13378 9976
rect 13320 9936 13326 9948
rect 13366 9945 13378 9948
rect 13412 9945 13424 9979
rect 14458 9976 14464 9988
rect 13366 9939 13424 9945
rect 13740 9948 14464 9976
rect 13740 9908 13768 9948
rect 14458 9936 14464 9948
rect 14516 9936 14522 9988
rect 14553 9979 14611 9985
rect 14553 9945 14565 9979
rect 14599 9976 14611 9979
rect 15396 9976 15424 10016
rect 14599 9948 15424 9976
rect 15464 9979 15522 9985
rect 14599 9945 14611 9948
rect 14553 9939 14611 9945
rect 15464 9945 15476 9979
rect 15510 9945 15522 9979
rect 15464 9939 15522 9945
rect 12360 9880 13768 9908
rect 12253 9871 12311 9877
rect 13814 9868 13820 9920
rect 13872 9908 13878 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13872 9880 14105 9908
rect 13872 9868 13878 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 14093 9871 14151 9877
rect 14826 9868 14832 9920
rect 14884 9908 14890 9920
rect 15488 9908 15516 9939
rect 15838 9936 15844 9988
rect 15896 9976 15902 9988
rect 17966 9979 18024 9985
rect 17966 9976 17978 9979
rect 15896 9948 17978 9976
rect 15896 9936 15902 9948
rect 17966 9945 17978 9948
rect 18012 9945 18024 9979
rect 18984 9976 19012 10016
rect 19705 10013 19717 10047
rect 19751 10044 19763 10047
rect 20070 10044 20076 10056
rect 19751 10016 20076 10044
rect 19751 10013 19763 10016
rect 19705 10007 19763 10013
rect 20070 10004 20076 10016
rect 20128 10004 20134 10056
rect 20162 9976 20168 9988
rect 17966 9939 18024 9945
rect 18064 9948 18920 9976
rect 18984 9948 20168 9976
rect 14884 9880 15516 9908
rect 14884 9868 14890 9880
rect 17310 9868 17316 9920
rect 17368 9908 17374 9920
rect 18064 9908 18092 9948
rect 17368 9880 18092 9908
rect 17368 9868 17374 9880
rect 18138 9868 18144 9920
rect 18196 9908 18202 9920
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 18196 9880 18797 9908
rect 18196 9868 18202 9880
rect 18785 9877 18797 9880
rect 18831 9877 18843 9911
rect 18892 9908 18920 9948
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 19521 9911 19579 9917
rect 19521 9908 19533 9911
rect 18892 9880 19533 9908
rect 18785 9871 18843 9877
rect 19521 9877 19533 9880
rect 19567 9877 19579 9911
rect 19521 9871 19579 9877
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 4154 9704 4160 9716
rect 1872 9676 4160 9704
rect 1489 9639 1547 9645
rect 1489 9605 1501 9639
rect 1535 9636 1547 9639
rect 1872 9636 1900 9676
rect 4154 9664 4160 9676
rect 4212 9704 4218 9716
rect 9490 9704 9496 9716
rect 4212 9676 9496 9704
rect 4212 9664 4218 9676
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 10870 9704 10876 9716
rect 10831 9676 10876 9704
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 11054 9664 11060 9716
rect 11112 9704 11118 9716
rect 11790 9704 11796 9716
rect 11112 9676 11796 9704
rect 11112 9664 11118 9676
rect 11790 9664 11796 9676
rect 11848 9664 11854 9716
rect 12434 9664 12440 9716
rect 12492 9704 12498 9716
rect 12492 9676 19288 9704
rect 12492 9664 12498 9676
rect 1535 9608 1900 9636
rect 1964 9608 2774 9636
rect 1535 9605 1547 9608
rect 1489 9599 1547 9605
rect 1964 9509 1992 9608
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9469 2007 9503
rect 1949 9463 2007 9469
rect 2041 9503 2099 9509
rect 2041 9469 2053 9503
rect 2087 9500 2099 9503
rect 2314 9500 2320 9512
rect 2087 9472 2320 9500
rect 2087 9469 2099 9472
rect 2041 9463 2099 9469
rect 2314 9460 2320 9472
rect 2372 9460 2378 9512
rect 2746 9500 2774 9608
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 3237 9639 3295 9645
rect 3237 9636 3249 9639
rect 3016 9608 3249 9636
rect 3016 9596 3022 9608
rect 3237 9605 3249 9608
rect 3283 9636 3295 9639
rect 4062 9636 4068 9648
rect 3283 9608 4068 9636
rect 3283 9605 3295 9608
rect 3237 9599 3295 9605
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 5074 9636 5080 9648
rect 4172 9608 5080 9636
rect 3142 9568 3148 9580
rect 3103 9540 3148 9568
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3878 9568 3884 9580
rect 3252 9540 3464 9568
rect 3839 9540 3884 9568
rect 3252 9500 3280 9540
rect 2746 9472 3280 9500
rect 3329 9503 3387 9509
rect 3329 9469 3341 9503
rect 3375 9469 3387 9503
rect 3329 9463 3387 9469
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 3344 9432 3372 9463
rect 1912 9404 3372 9432
rect 3436 9432 3464 9540
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 4172 9500 4200 9608
rect 5074 9596 5080 9608
rect 5132 9596 5138 9648
rect 5718 9596 5724 9648
rect 5776 9636 5782 9648
rect 8570 9636 8576 9648
rect 5776 9608 8576 9636
rect 5776 9596 5782 9608
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 9122 9596 9128 9648
rect 9180 9596 9186 9648
rect 9214 9596 9220 9648
rect 9272 9636 9278 9648
rect 9272 9608 9674 9636
rect 9272 9596 9278 9608
rect 4430 9528 4436 9580
rect 4488 9568 4494 9580
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 4488 9540 4537 9568
rect 4488 9528 4494 9540
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5350 9568 5356 9580
rect 5215 9540 5356 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 5994 9568 6000 9580
rect 5500 9540 6000 9568
rect 5500 9528 5506 9540
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 6822 9528 6828 9580
rect 6880 9568 6886 9580
rect 7009 9571 7067 9577
rect 7009 9568 7021 9571
rect 6880 9540 7021 9568
rect 6880 9528 6886 9540
rect 7009 9537 7021 9540
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 8389 9571 8447 9577
rect 8389 9568 8401 9571
rect 7791 9540 8401 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 8389 9537 8401 9540
rect 8435 9537 8447 9571
rect 9140 9568 9168 9596
rect 9473 9571 9531 9577
rect 9473 9568 9485 9571
rect 8389 9531 8447 9537
rect 8588 9540 9485 9568
rect 4890 9500 4896 9512
rect 3752 9472 4200 9500
rect 4264 9472 4896 9500
rect 3752 9460 3758 9472
rect 4264 9432 4292 9472
rect 4890 9460 4896 9472
rect 4948 9460 4954 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5626 9500 5632 9512
rect 5123 9472 5632 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9500 6791 9503
rect 7837 9503 7895 9509
rect 7837 9500 7849 9503
rect 6779 9472 7849 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 7837 9469 7849 9472
rect 7883 9469 7895 9503
rect 7837 9463 7895 9469
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8294 9500 8300 9512
rect 8067 9472 8300 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 3436 9404 4292 9432
rect 4341 9435 4399 9441
rect 1912 9392 1918 9404
rect 4341 9401 4353 9435
rect 4387 9432 4399 9435
rect 4522 9432 4528 9444
rect 4387 9404 4528 9432
rect 4387 9401 4399 9404
rect 4341 9395 4399 9401
rect 4522 9392 4528 9404
rect 4580 9392 4586 9444
rect 6748 9432 6776 9463
rect 4816 9404 6776 9432
rect 7852 9432 7880 9463
rect 8294 9460 8300 9472
rect 8352 9500 8358 9512
rect 8588 9500 8616 9540
rect 9473 9537 9485 9540
rect 9519 9537 9531 9571
rect 9646 9568 9674 9608
rect 10778 9596 10784 9648
rect 10836 9636 10842 9648
rect 10888 9636 10916 9664
rect 16669 9639 16727 9645
rect 16669 9636 16681 9639
rect 10836 9608 10916 9636
rect 14180 9608 16681 9636
rect 10836 9596 10842 9608
rect 9646 9540 11744 9568
rect 9473 9531 9531 9537
rect 8352 9472 8616 9500
rect 8352 9460 8358 9472
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9217 9503 9275 9509
rect 9217 9500 9229 9503
rect 9180 9472 9229 9500
rect 9180 9460 9186 9472
rect 9217 9469 9229 9472
rect 9263 9469 9275 9503
rect 9217 9463 9275 9469
rect 11716 9444 11744 9540
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 12906 9571 12964 9577
rect 12906 9568 12918 9571
rect 12400 9540 12918 9568
rect 12400 9528 12406 9540
rect 12906 9537 12918 9540
rect 12952 9537 12964 9571
rect 12906 9531 12964 9537
rect 13078 9528 13084 9580
rect 13136 9568 13142 9580
rect 14180 9577 14208 9608
rect 16669 9605 16681 9608
rect 16715 9636 16727 9639
rect 17494 9636 17500 9648
rect 16715 9608 17500 9636
rect 16715 9605 16727 9608
rect 16669 9599 16727 9605
rect 17494 9596 17500 9608
rect 17552 9596 17558 9648
rect 19260 9636 19288 9676
rect 20162 9664 20168 9716
rect 20220 9704 20226 9716
rect 20438 9704 20444 9716
rect 20220 9676 20444 9704
rect 20220 9664 20226 9676
rect 20438 9664 20444 9676
rect 20496 9664 20502 9716
rect 19260 9608 20576 9636
rect 20548 9580 20576 9608
rect 14165 9571 14223 9577
rect 14165 9568 14177 9571
rect 13136 9540 14177 9568
rect 13136 9528 13142 9540
rect 14165 9537 14177 9540
rect 14211 9537 14223 9571
rect 14165 9531 14223 9537
rect 16301 9571 16359 9577
rect 16301 9537 16313 9571
rect 16347 9568 16359 9571
rect 17405 9571 17463 9577
rect 17405 9568 17417 9571
rect 16347 9540 17417 9568
rect 16347 9537 16359 9540
rect 16301 9531 16359 9537
rect 17405 9537 17417 9540
rect 17451 9537 17463 9571
rect 17405 9531 17463 9537
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 18230 9568 18236 9580
rect 17920 9540 18236 9568
rect 17920 9528 17926 9540
rect 18230 9528 18236 9540
rect 18288 9568 18294 9580
rect 19438 9571 19496 9577
rect 19438 9568 19450 9571
rect 18288 9540 19450 9568
rect 18288 9528 18294 9540
rect 19438 9537 19450 9540
rect 19484 9537 19496 9571
rect 19438 9531 19496 9537
rect 19610 9528 19616 9580
rect 19668 9568 19674 9580
rect 20257 9571 20315 9577
rect 20257 9568 20269 9571
rect 19668 9540 20269 9568
rect 19668 9528 19674 9540
rect 20257 9537 20269 9540
rect 20303 9537 20315 9571
rect 20530 9568 20536 9580
rect 20443 9540 20536 9568
rect 20257 9531 20315 9537
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 13173 9503 13231 9509
rect 13173 9469 13185 9503
rect 13219 9469 13231 9503
rect 13814 9500 13820 9512
rect 13173 9463 13231 9469
rect 13556 9472 13820 9500
rect 7852 9404 8984 9432
rect 2501 9367 2559 9373
rect 2501 9333 2513 9367
rect 2547 9364 2559 9367
rect 2590 9364 2596 9376
rect 2547 9336 2596 9364
rect 2547 9333 2559 9336
rect 2501 9327 2559 9333
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 2832 9336 2877 9364
rect 2832 9324 2838 9336
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 3510 9364 3516 9376
rect 3016 9336 3516 9364
rect 3016 9324 3022 9336
rect 3510 9324 3516 9336
rect 3568 9324 3574 9376
rect 3973 9367 4031 9373
rect 3973 9333 3985 9367
rect 4019 9364 4031 9367
rect 4816 9364 4844 9404
rect 5534 9364 5540 9376
rect 4019 9336 4844 9364
rect 5495 9336 5540 9364
rect 4019 9333 4031 9336
rect 3973 9327 4031 9333
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5905 9367 5963 9373
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 5994 9364 6000 9376
rect 5951 9336 6000 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 7377 9367 7435 9373
rect 7377 9364 7389 9367
rect 7340 9336 7389 9364
rect 7340 9324 7346 9336
rect 7377 9333 7389 9336
rect 7423 9333 7435 9367
rect 7377 9327 7435 9333
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 7524 9336 8861 9364
rect 7524 9324 7530 9336
rect 8849 9333 8861 9336
rect 8895 9333 8907 9367
rect 8956 9364 8984 9404
rect 11698 9392 11704 9444
rect 11756 9432 11762 9444
rect 12066 9432 12072 9444
rect 11756 9404 12072 9432
rect 11756 9392 11762 9404
rect 12066 9392 12072 9404
rect 12124 9392 12130 9444
rect 13188 9432 13216 9463
rect 13556 9444 13584 9472
rect 13814 9460 13820 9472
rect 13872 9500 13878 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13872 9472 13921 9500
rect 13872 9460 13878 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 17494 9500 17500 9512
rect 17455 9472 17500 9500
rect 13909 9463 13967 9469
rect 17494 9460 17500 9472
rect 17552 9460 17558 9512
rect 17586 9460 17592 9512
rect 17644 9500 17650 9512
rect 19702 9500 19708 9512
rect 17644 9472 17689 9500
rect 19663 9472 19708 9500
rect 17644 9460 17650 9472
rect 19702 9460 19708 9472
rect 19760 9460 19766 9512
rect 20806 9500 20812 9512
rect 20767 9472 20812 9500
rect 20806 9460 20812 9472
rect 20864 9460 20870 9512
rect 13538 9432 13544 9444
rect 13188 9404 13544 9432
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 15470 9392 15476 9444
rect 15528 9432 15534 9444
rect 17037 9435 17095 9441
rect 17037 9432 17049 9435
rect 15528 9404 17049 9432
rect 15528 9392 15534 9404
rect 17037 9401 17049 9404
rect 17083 9401 17095 9435
rect 17037 9395 17095 9401
rect 17678 9392 17684 9444
rect 17736 9432 17742 9444
rect 18325 9435 18383 9441
rect 18325 9432 18337 9435
rect 17736 9404 18337 9432
rect 17736 9392 17742 9404
rect 18325 9401 18337 9404
rect 18371 9401 18383 9435
rect 18325 9395 18383 9401
rect 19886 9392 19892 9444
rect 19944 9432 19950 9444
rect 20073 9435 20131 9441
rect 20073 9432 20085 9435
rect 19944 9404 20085 9432
rect 19944 9392 19950 9404
rect 20073 9401 20085 9404
rect 20119 9401 20131 9435
rect 20073 9395 20131 9401
rect 9398 9364 9404 9376
rect 8956 9336 9404 9364
rect 8849 9327 8907 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 10594 9364 10600 9376
rect 10555 9336 10600 9364
rect 10594 9324 10600 9336
rect 10652 9324 10658 9376
rect 11793 9367 11851 9373
rect 11793 9333 11805 9367
rect 11839 9364 11851 9367
rect 12986 9364 12992 9376
rect 11839 9336 12992 9364
rect 11839 9333 11851 9336
rect 11793 9327 11851 9333
rect 12986 9324 12992 9336
rect 13044 9324 13050 9376
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 13504 9336 15301 9364
rect 13504 9324 13510 9336
rect 15289 9333 15301 9336
rect 15335 9333 15347 9367
rect 15562 9364 15568 9376
rect 15523 9336 15568 9364
rect 15289 9327 15347 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 16206 9324 16212 9376
rect 16264 9364 16270 9376
rect 19978 9364 19984 9376
rect 16264 9336 19984 9364
rect 16264 9324 16270 9336
rect 19978 9324 19984 9336
rect 20036 9364 20042 9376
rect 20622 9364 20628 9376
rect 20036 9336 20628 9364
rect 20036 9324 20042 9336
rect 20622 9324 20628 9336
rect 20680 9324 20686 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 5718 9160 5724 9172
rect 2240 9132 5724 9160
rect 1762 8984 1768 9036
rect 1820 9024 1826 9036
rect 1949 9027 2007 9033
rect 1949 9024 1961 9027
rect 1820 8996 1961 9024
rect 1820 8984 1826 8996
rect 1949 8993 1961 8996
rect 1995 8993 2007 9027
rect 1949 8987 2007 8993
rect 2240 8968 2268 9132
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 7006 9120 7012 9172
rect 7064 9160 7070 9172
rect 7929 9163 7987 9169
rect 7929 9160 7941 9163
rect 7064 9132 7941 9160
rect 7064 9120 7070 9132
rect 7929 9129 7941 9132
rect 7975 9160 7987 9163
rect 8018 9160 8024 9172
rect 7975 9132 8024 9160
rect 7975 9129 7987 9132
rect 7929 9123 7987 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9160 8631 9163
rect 9214 9160 9220 9172
rect 8619 9132 9220 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 9309 9163 9367 9169
rect 9309 9129 9321 9163
rect 9355 9160 9367 9163
rect 9582 9160 9588 9172
rect 9355 9132 9588 9160
rect 9355 9129 9367 9132
rect 9309 9123 9367 9129
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 9692 9132 10732 9160
rect 3050 9092 3056 9104
rect 2516 9064 3056 9092
rect 2222 8956 2228 8968
rect 2183 8928 2228 8956
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 2516 8897 2544 9064
rect 3050 9052 3056 9064
rect 3108 9052 3114 9104
rect 4522 9052 4528 9104
rect 4580 9092 4586 9104
rect 5350 9092 5356 9104
rect 4580 9064 5356 9092
rect 4580 9052 4586 9064
rect 5350 9052 5356 9064
rect 5408 9092 5414 9104
rect 6273 9095 6331 9101
rect 6273 9092 6285 9095
rect 5408 9064 6285 9092
rect 5408 9052 5414 9064
rect 6273 9061 6285 9064
rect 6319 9092 6331 9095
rect 7558 9092 7564 9104
rect 6319 9064 7564 9092
rect 6319 9061 6331 9064
rect 6273 9055 6331 9061
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 7653 9095 7711 9101
rect 7653 9061 7665 9095
rect 7699 9092 7711 9095
rect 8478 9092 8484 9104
rect 7699 9064 8484 9092
rect 7699 9061 7711 9064
rect 7653 9055 7711 9061
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 9030 9052 9036 9104
rect 9088 9092 9094 9104
rect 9692 9092 9720 9132
rect 9088 9064 9720 9092
rect 10704 9092 10732 9132
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 10965 9163 11023 9169
rect 10965 9160 10977 9163
rect 10928 9132 10977 9160
rect 10928 9120 10934 9132
rect 10965 9129 10977 9132
rect 11011 9129 11023 9163
rect 10965 9123 11023 9129
rect 11238 9120 11244 9172
rect 11296 9160 11302 9172
rect 16298 9160 16304 9172
rect 11296 9132 16304 9160
rect 11296 9120 11302 9132
rect 16298 9120 16304 9132
rect 16356 9120 16362 9172
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 19794 9160 19800 9172
rect 17276 9132 19656 9160
rect 19755 9132 19800 9160
rect 17276 9120 17282 9132
rect 11146 9092 11152 9104
rect 10704 9064 11152 9092
rect 9088 9052 9094 9064
rect 11146 9052 11152 9064
rect 11204 9092 11210 9104
rect 11514 9092 11520 9104
rect 11204 9064 11520 9092
rect 11204 9052 11210 9064
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 14185 9095 14243 9101
rect 14185 9061 14197 9095
rect 14231 9092 14243 9095
rect 14274 9092 14280 9104
rect 14231 9064 14280 9092
rect 14231 9061 14243 9064
rect 14185 9055 14243 9061
rect 14274 9052 14280 9064
rect 14332 9052 14338 9104
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 19337 9095 19395 9101
rect 19337 9092 19349 9095
rect 17828 9064 19349 9092
rect 17828 9052 17834 9064
rect 19337 9061 19349 9064
rect 19383 9061 19395 9095
rect 19337 9055 19395 9061
rect 3142 9024 3148 9036
rect 3103 8996 3148 9024
rect 3142 8984 3148 8996
rect 3200 8984 3206 9036
rect 3973 9027 4031 9033
rect 3973 8993 3985 9027
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 3988 8956 4016 8987
rect 4430 8984 4436 9036
rect 4488 9024 4494 9036
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 4488 8996 5457 9024
rect 4488 8984 4494 8996
rect 5445 8993 5457 8996
rect 5491 9024 5503 9027
rect 6822 9024 6828 9036
rect 5491 8996 6828 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7101 9027 7159 9033
rect 7101 8993 7113 9027
rect 7147 9024 7159 9027
rect 10689 9027 10747 9033
rect 7147 8996 9720 9024
rect 7147 8993 7159 8996
rect 7101 8987 7159 8993
rect 4890 8956 4896 8968
rect 3988 8928 4896 8956
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8956 5319 8959
rect 5534 8956 5540 8968
rect 5307 8928 5540 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 7282 8956 7288 8968
rect 7243 8928 7288 8956
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 9692 8956 9720 8996
rect 10689 8993 10701 9027
rect 10735 9024 10747 9027
rect 10870 9024 10876 9036
rect 10735 8996 10876 9024
rect 10735 8993 10747 8996
rect 10689 8987 10747 8993
rect 10870 8984 10876 8996
rect 10928 9024 10934 9036
rect 11885 9027 11943 9033
rect 11885 9024 11897 9027
rect 10928 8996 11897 9024
rect 10928 8984 10934 8996
rect 11885 8993 11897 8996
rect 11931 8993 11943 9027
rect 15562 9024 15568 9036
rect 15523 8996 15568 9024
rect 11885 8987 11943 8993
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 18049 9027 18107 9033
rect 18049 8993 18061 9027
rect 18095 9024 18107 9027
rect 18095 8996 18460 9024
rect 18095 8993 18107 8996
rect 18049 8987 18107 8993
rect 10594 8956 10600 8968
rect 9692 8928 10600 8956
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 12141 8959 12199 8965
rect 12141 8956 12153 8959
rect 11572 8928 12153 8956
rect 11572 8916 11578 8928
rect 12141 8925 12153 8928
rect 12187 8925 12199 8959
rect 13541 8959 13599 8965
rect 13541 8956 13553 8959
rect 12141 8919 12199 8925
rect 12406 8928 13553 8956
rect 12406 8900 12434 8928
rect 13541 8925 13553 8928
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 14550 8916 14556 8968
rect 14608 8956 14614 8968
rect 15654 8956 15660 8968
rect 14608 8928 15660 8956
rect 14608 8916 14614 8928
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 17497 8959 17555 8965
rect 17497 8925 17509 8959
rect 17543 8956 17555 8959
rect 17954 8956 17960 8968
rect 17543 8928 17960 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 17954 8916 17960 8928
rect 18012 8956 18018 8968
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 18012 8928 18337 8956
rect 18012 8916 18018 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 2501 8891 2559 8897
rect 2501 8888 2513 8891
rect 2464 8860 2513 8888
rect 2464 8848 2470 8860
rect 2501 8857 2513 8860
rect 2547 8857 2559 8891
rect 2501 8851 2559 8857
rect 2685 8891 2743 8897
rect 2685 8857 2697 8891
rect 2731 8888 2743 8891
rect 3142 8888 3148 8900
rect 2731 8860 3148 8888
rect 2731 8857 2743 8860
rect 2685 8851 2743 8857
rect 3142 8848 3148 8860
rect 3200 8848 3206 8900
rect 3786 8848 3792 8900
rect 3844 8888 3850 8900
rect 4157 8891 4215 8897
rect 4157 8888 4169 8891
rect 3844 8860 4169 8888
rect 3844 8848 3850 8860
rect 4157 8857 4169 8860
rect 4203 8857 4215 8891
rect 5353 8891 5411 8897
rect 5353 8888 5365 8891
rect 4157 8851 4215 8857
rect 4540 8860 5365 8888
rect 4065 8823 4123 8829
rect 4065 8789 4077 8823
rect 4111 8820 4123 8823
rect 4246 8820 4252 8832
rect 4111 8792 4252 8820
rect 4111 8789 4123 8792
rect 4065 8783 4123 8789
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4540 8829 4568 8860
rect 5353 8857 5365 8860
rect 5399 8857 5411 8891
rect 5353 8851 5411 8857
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 10134 8888 10140 8900
rect 9732 8860 10140 8888
rect 9732 8848 9738 8860
rect 10134 8848 10140 8860
rect 10192 8848 10198 8900
rect 10444 8891 10502 8897
rect 10444 8857 10456 8891
rect 10490 8888 10502 8891
rect 11974 8888 11980 8900
rect 10490 8860 11980 8888
rect 10490 8857 10502 8860
rect 10444 8851 10502 8857
rect 11974 8848 11980 8860
rect 12032 8848 12038 8900
rect 12342 8848 12348 8900
rect 12400 8860 12434 8900
rect 12400 8848 12406 8860
rect 12802 8848 12808 8900
rect 12860 8888 12866 8900
rect 13446 8888 13452 8900
rect 12860 8860 13452 8888
rect 12860 8848 12866 8860
rect 13446 8848 13452 8860
rect 13504 8848 13510 8900
rect 15286 8848 15292 8900
rect 15344 8897 15350 8900
rect 15344 8888 15356 8897
rect 17034 8888 17040 8900
rect 15344 8860 15389 8888
rect 16049 8860 17040 8888
rect 15344 8851 15356 8860
rect 15344 8848 15350 8851
rect 4525 8823 4583 8829
rect 4525 8789 4537 8823
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 4893 8823 4951 8829
rect 4893 8789 4905 8823
rect 4939 8820 4951 8823
rect 5074 8820 5080 8832
rect 4939 8792 5080 8820
rect 4939 8789 4951 8792
rect 4893 8783 4951 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 5905 8823 5963 8829
rect 5905 8820 5917 8823
rect 5776 8792 5917 8820
rect 5776 8780 5782 8792
rect 5905 8789 5917 8792
rect 5951 8789 5963 8823
rect 5905 8783 5963 8789
rect 7193 8823 7251 8829
rect 7193 8789 7205 8823
rect 7239 8820 7251 8823
rect 7282 8820 7288 8832
rect 7239 8792 7288 8820
rect 7239 8789 7251 8792
rect 7193 8783 7251 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 9033 8823 9091 8829
rect 9033 8789 9045 8823
rect 9079 8820 9091 8823
rect 9214 8820 9220 8832
rect 9079 8792 9220 8820
rect 9079 8789 9091 8792
rect 9033 8783 9091 8789
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 9490 8780 9496 8832
rect 9548 8820 9554 8832
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 9548 8792 13277 8820
rect 9548 8780 9554 8792
rect 13265 8789 13277 8792
rect 13311 8820 13323 8823
rect 16049 8820 16077 8860
rect 17034 8848 17040 8860
rect 17092 8848 17098 8900
rect 17218 8888 17224 8900
rect 17276 8897 17282 8900
rect 17188 8860 17224 8888
rect 17218 8848 17224 8860
rect 17276 8851 17288 8897
rect 17865 8891 17923 8897
rect 17865 8888 17877 8891
rect 17328 8860 17877 8888
rect 17276 8848 17282 8851
rect 13311 8792 16077 8820
rect 13311 8789 13323 8792
rect 13265 8783 13323 8789
rect 16114 8780 16120 8832
rect 16172 8820 16178 8832
rect 17328 8820 17356 8860
rect 17865 8857 17877 8860
rect 17911 8857 17923 8891
rect 17865 8851 17923 8857
rect 16172 8792 17356 8820
rect 18340 8820 18368 8919
rect 18432 8888 18460 8996
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 19116 8928 19533 8956
rect 19116 8916 19122 8928
rect 19521 8925 19533 8928
rect 19567 8925 19579 8959
rect 19628 8956 19656 9132
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 20162 8984 20168 9036
rect 20220 9024 20226 9036
rect 20349 9027 20407 9033
rect 20349 9024 20361 9027
rect 20220 8996 20361 9024
rect 20220 8984 20226 8996
rect 20349 8993 20361 8996
rect 20395 8993 20407 9027
rect 20349 8987 20407 8993
rect 21266 8956 21272 8968
rect 19628 8928 21272 8956
rect 19521 8919 19579 8925
rect 21266 8916 21272 8928
rect 21324 8916 21330 8968
rect 19334 8888 19340 8900
rect 18432 8860 19340 8888
rect 19334 8848 19340 8860
rect 19392 8888 19398 8900
rect 21082 8888 21088 8900
rect 19392 8860 20484 8888
rect 21043 8860 21088 8888
rect 19392 8848 19398 8860
rect 18690 8820 18696 8832
rect 18340 8792 18696 8820
rect 16172 8780 16178 8792
rect 18690 8780 18696 8792
rect 18748 8780 18754 8832
rect 20162 8820 20168 8832
rect 20123 8792 20168 8820
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 20254 8780 20260 8832
rect 20312 8820 20318 8832
rect 20456 8820 20484 8860
rect 21082 8848 21088 8860
rect 21140 8848 21146 8900
rect 20530 8820 20536 8832
rect 20312 8792 20357 8820
rect 20443 8792 20536 8820
rect 20312 8780 20318 8792
rect 20530 8780 20536 8792
rect 20588 8820 20594 8832
rect 21358 8820 21364 8832
rect 20588 8792 21364 8820
rect 20588 8780 20594 8792
rect 21358 8780 21364 8792
rect 21416 8780 21422 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 3513 8619 3571 8625
rect 3513 8616 3525 8619
rect 2188 8588 3525 8616
rect 2188 8576 2194 8588
rect 3513 8585 3525 8588
rect 3559 8585 3571 8619
rect 3513 8579 3571 8585
rect 3970 8576 3976 8628
rect 4028 8616 4034 8628
rect 5813 8619 5871 8625
rect 5813 8616 5825 8619
rect 4028 8588 5825 8616
rect 4028 8576 4034 8588
rect 5813 8585 5825 8588
rect 5859 8585 5871 8619
rect 5813 8579 5871 8585
rect 6457 8619 6515 8625
rect 6457 8585 6469 8619
rect 6503 8616 6515 8619
rect 6638 8616 6644 8628
rect 6503 8588 6644 8616
rect 6503 8585 6515 8588
rect 6457 8579 6515 8585
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 8754 8616 8760 8628
rect 8715 8588 8760 8616
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9122 8616 9128 8628
rect 9048 8588 9128 8616
rect 2961 8551 3019 8557
rect 2961 8517 2973 8551
rect 3007 8548 3019 8551
rect 5350 8548 5356 8560
rect 3007 8520 5356 8548
rect 3007 8517 3019 8520
rect 2961 8511 3019 8517
rect 5350 8508 5356 8520
rect 5408 8508 5414 8560
rect 7190 8508 7196 8560
rect 7248 8548 7254 8560
rect 7561 8551 7619 8557
rect 7561 8548 7573 8551
rect 7248 8520 7573 8548
rect 7248 8508 7254 8520
rect 7561 8517 7573 8520
rect 7607 8548 7619 8551
rect 8202 8548 8208 8560
rect 7607 8520 8208 8548
rect 7607 8517 7619 8520
rect 7561 8511 7619 8517
rect 8202 8508 8208 8520
rect 8260 8508 8266 8560
rect 1486 8440 1492 8492
rect 1544 8480 1550 8492
rect 1949 8483 2007 8489
rect 1949 8480 1961 8483
rect 1544 8452 1961 8480
rect 1544 8440 1550 8452
rect 1949 8449 1961 8452
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 2869 8483 2927 8489
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 4706 8480 4712 8492
rect 2915 8452 4712 8480
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 4706 8440 4712 8452
rect 4764 8480 4770 8492
rect 5077 8483 5135 8489
rect 4764 8452 4936 8480
rect 4764 8440 4770 8452
rect 2222 8412 2228 8424
rect 2183 8384 2228 8412
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 3142 8412 3148 8424
rect 3103 8384 3148 8412
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 4065 8415 4123 8421
rect 4065 8381 4077 8415
rect 4111 8412 4123 8415
rect 4154 8412 4160 8424
rect 4111 8384 4160 8412
rect 4111 8381 4123 8384
rect 4065 8375 4123 8381
rect 4154 8372 4160 8384
rect 4212 8372 4218 8424
rect 4246 8372 4252 8424
rect 4304 8412 4310 8424
rect 4433 8415 4491 8421
rect 4433 8412 4445 8415
rect 4304 8384 4445 8412
rect 4304 8372 4310 8384
rect 4433 8381 4445 8384
rect 4479 8381 4491 8415
rect 4908 8412 4936 8452
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5442 8480 5448 8492
rect 5123 8452 5448 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 7469 8483 7527 8489
rect 7469 8480 7481 8483
rect 5684 8452 7481 8480
rect 5684 8440 5690 8452
rect 7469 8449 7481 8452
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 5534 8412 5540 8424
rect 4908 8384 5540 8412
rect 4433 8375 4491 8381
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 8294 8412 8300 8424
rect 7791 8384 8300 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 2501 8347 2559 8353
rect 2501 8313 2513 8347
rect 2547 8344 2559 8347
rect 2682 8344 2688 8356
rect 2547 8316 2688 8344
rect 2547 8313 2559 8316
rect 2501 8307 2559 8313
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 3786 8304 3792 8356
rect 3844 8344 3850 8356
rect 3970 8344 3976 8356
rect 3844 8316 3976 8344
rect 3844 8304 3850 8316
rect 3970 8304 3976 8316
rect 4028 8344 4034 8356
rect 6638 8344 6644 8356
rect 4028 8316 6644 8344
rect 4028 8304 4034 8316
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 7101 8347 7159 8353
rect 7101 8313 7113 8347
rect 7147 8344 7159 8347
rect 7282 8344 7288 8356
rect 7147 8316 7288 8344
rect 7147 8313 7159 8316
rect 7101 8307 7159 8313
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 9048 8344 9076 8588
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 9548 8588 9996 8616
rect 9548 8576 9554 8588
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 9364 8520 9628 8548
rect 9364 8508 9370 8520
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 9600 8480 9628 8520
rect 9766 8508 9772 8560
rect 9824 8508 9830 8560
rect 9968 8548 9996 8588
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 10100 8588 10793 8616
rect 10100 8576 10106 8588
rect 10781 8585 10793 8588
rect 10827 8585 10839 8619
rect 10781 8579 10839 8585
rect 11701 8619 11759 8625
rect 11701 8585 11713 8619
rect 11747 8616 11759 8619
rect 12250 8616 12256 8628
rect 11747 8588 12256 8616
rect 11747 8585 11759 8588
rect 11701 8579 11759 8585
rect 12250 8576 12256 8588
rect 12308 8576 12314 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 16114 8616 16120 8628
rect 13412 8588 16120 8616
rect 13412 8576 13418 8588
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 16356 8588 16681 8616
rect 16356 8576 16362 8588
rect 16669 8585 16681 8588
rect 16715 8585 16727 8619
rect 16669 8579 16727 8585
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 20073 8619 20131 8625
rect 20073 8616 20085 8619
rect 17552 8588 20085 8616
rect 17552 8576 17558 8588
rect 20073 8585 20085 8588
rect 20119 8585 20131 8619
rect 20438 8616 20444 8628
rect 20399 8588 20444 8616
rect 20073 8579 20131 8585
rect 20438 8576 20444 8588
rect 20496 8576 20502 8628
rect 15194 8548 15200 8560
rect 9968 8520 15200 8548
rect 15194 8508 15200 8520
rect 15252 8508 15258 8560
rect 15286 8508 15292 8560
rect 15344 8548 15350 8560
rect 16025 8551 16083 8557
rect 16025 8548 16037 8551
rect 15344 8520 16037 8548
rect 15344 8508 15350 8520
rect 16025 8517 16037 8520
rect 16071 8517 16083 8551
rect 16025 8511 16083 8517
rect 17218 8508 17224 8560
rect 17276 8548 17282 8560
rect 17402 8548 17408 8560
rect 17276 8520 17408 8548
rect 17276 8508 17282 8520
rect 17402 8508 17408 8520
rect 17460 8508 17466 8560
rect 17678 8508 17684 8560
rect 17736 8548 17742 8560
rect 17782 8551 17840 8557
rect 17782 8548 17794 8551
rect 17736 8520 17794 8548
rect 17736 8508 17742 8520
rect 17782 8517 17794 8520
rect 17828 8548 17840 8551
rect 18230 8548 18236 8560
rect 17828 8520 18236 8548
rect 17828 8517 17840 8520
rect 17782 8511 17840 8517
rect 18230 8508 18236 8520
rect 18288 8508 18294 8560
rect 18322 8508 18328 8560
rect 18380 8548 18386 8560
rect 18690 8548 18696 8560
rect 18380 8520 18425 8548
rect 18651 8520 18696 8548
rect 18380 8508 18386 8520
rect 18690 8508 18696 8520
rect 18748 8508 18754 8560
rect 19334 8508 19340 8560
rect 19392 8508 19398 8560
rect 19518 8508 19524 8560
rect 19576 8548 19582 8560
rect 20533 8551 20591 8557
rect 20533 8548 20545 8551
rect 19576 8520 20545 8548
rect 19576 8508 19582 8520
rect 20533 8517 20545 8520
rect 20579 8517 20591 8551
rect 20533 8511 20591 8517
rect 21269 8551 21327 8557
rect 21269 8517 21281 8551
rect 21315 8548 21327 8551
rect 21358 8548 21364 8560
rect 21315 8520 21364 8548
rect 21315 8517 21327 8520
rect 21269 8511 21327 8517
rect 21358 8508 21364 8520
rect 21416 8508 21422 8560
rect 9657 8483 9715 8489
rect 9657 8480 9669 8483
rect 9456 8452 9501 8480
rect 9600 8452 9669 8480
rect 9456 8440 9462 8452
rect 9657 8449 9669 8452
rect 9703 8449 9715 8483
rect 9784 8480 9812 8508
rect 13101 8483 13159 8489
rect 9784 8452 12020 8480
rect 9657 8443 9715 8449
rect 9398 8344 9404 8356
rect 9048 8316 9404 8344
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 11992 8353 12020 8452
rect 13101 8449 13113 8483
rect 13147 8480 13159 8483
rect 13262 8480 13268 8492
rect 13147 8452 13268 8480
rect 13147 8449 13159 8452
rect 13101 8443 13159 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 14642 8480 14648 8492
rect 14603 8452 14648 8480
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 15013 8483 15071 8489
rect 15013 8449 15025 8483
rect 15059 8480 15071 8483
rect 19058 8480 19064 8492
rect 15059 8452 19064 8480
rect 15059 8449 15071 8452
rect 15013 8443 15071 8449
rect 19058 8440 19064 8452
rect 19116 8440 19122 8492
rect 19352 8480 19380 8508
rect 19260 8452 19380 8480
rect 19429 8483 19487 8489
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8412 13415 8415
rect 13538 8412 13544 8424
rect 13403 8384 13544 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 13538 8372 13544 8384
rect 13596 8412 13602 8424
rect 18049 8415 18107 8421
rect 13596 8384 13768 8412
rect 13596 8372 13602 8384
rect 11977 8347 12035 8353
rect 11977 8313 11989 8347
rect 12023 8313 12035 8347
rect 11977 8307 12035 8313
rect 6546 8236 6552 8288
rect 6604 8276 6610 8288
rect 6825 8279 6883 8285
rect 6825 8276 6837 8279
rect 6604 8248 6837 8276
rect 6604 8236 6610 8248
rect 6825 8245 6837 8248
rect 6871 8276 6883 8279
rect 9122 8276 9128 8288
rect 6871 8248 9128 8276
rect 6871 8245 6883 8248
rect 6825 8239 6883 8245
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 9416 8276 9444 8304
rect 10778 8276 10784 8288
rect 9416 8248 10784 8276
rect 10778 8236 10784 8248
rect 10836 8276 10842 8288
rect 11146 8276 11152 8288
rect 10836 8248 11152 8276
rect 10836 8236 10842 8248
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 13740 8285 13768 8384
rect 18049 8381 18061 8415
rect 18095 8412 18107 8415
rect 18690 8412 18696 8424
rect 18095 8384 18696 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 19260 8421 19288 8452
rect 19429 8449 19441 8483
rect 19475 8480 19487 8483
rect 19886 8480 19892 8492
rect 19475 8452 19892 8480
rect 19475 8449 19487 8452
rect 19429 8443 19487 8449
rect 19886 8440 19892 8452
rect 19944 8440 19950 8492
rect 20714 8480 20720 8492
rect 20548 8452 20720 8480
rect 19245 8415 19303 8421
rect 19245 8381 19257 8415
rect 19291 8381 19303 8415
rect 19245 8375 19303 8381
rect 19337 8415 19395 8421
rect 19337 8381 19349 8415
rect 19383 8412 19395 8415
rect 20548 8412 20576 8452
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 19383 8384 20576 8412
rect 19383 8381 19395 8384
rect 19337 8375 19395 8381
rect 20622 8372 20628 8424
rect 20680 8412 20686 8424
rect 20680 8384 20725 8412
rect 20680 8372 20686 8384
rect 15378 8344 15384 8356
rect 15339 8316 15384 8344
rect 15378 8304 15384 8316
rect 15436 8304 15442 8356
rect 18708 8344 18736 8372
rect 21082 8344 21088 8356
rect 18708 8316 20668 8344
rect 21043 8316 21088 8344
rect 19720 8288 19748 8316
rect 20640 8288 20668 8316
rect 21082 8304 21088 8316
rect 21140 8304 21146 8356
rect 13725 8279 13783 8285
rect 13725 8245 13737 8279
rect 13771 8276 13783 8279
rect 14093 8279 14151 8285
rect 14093 8276 14105 8279
rect 13771 8248 14105 8276
rect 13771 8245 13783 8248
rect 13725 8239 13783 8245
rect 14093 8245 14105 8248
rect 14139 8276 14151 8279
rect 15749 8279 15807 8285
rect 15749 8276 15761 8279
rect 14139 8248 15761 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 15749 8245 15761 8248
rect 15795 8276 15807 8279
rect 16114 8276 16120 8288
rect 15795 8248 16120 8276
rect 15795 8245 15807 8248
rect 15749 8239 15807 8245
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 17034 8236 17040 8288
rect 17092 8276 17098 8288
rect 19058 8276 19064 8288
rect 17092 8248 19064 8276
rect 17092 8236 17098 8248
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 19702 8236 19708 8288
rect 19760 8236 19766 8288
rect 19797 8279 19855 8285
rect 19797 8245 19809 8279
rect 19843 8276 19855 8279
rect 20438 8276 20444 8288
rect 19843 8248 20444 8276
rect 19843 8245 19855 8248
rect 19797 8239 19855 8245
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 20622 8236 20628 8288
rect 20680 8236 20686 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 2372 8044 3801 8072
rect 2372 8032 2378 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 3878 8032 3884 8084
rect 3936 8072 3942 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 3936 8044 4261 8072
rect 3936 8032 3942 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 5902 8072 5908 8084
rect 5863 8044 5908 8072
rect 4249 8035 4307 8041
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 6822 8032 6828 8084
rect 6880 8072 6886 8084
rect 8662 8072 8668 8084
rect 6880 8044 8668 8072
rect 6880 8032 6886 8044
rect 8662 8032 8668 8044
rect 8720 8072 8726 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8720 8044 8953 8072
rect 8720 8032 8726 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 9401 8075 9459 8081
rect 9401 8041 9413 8075
rect 9447 8072 9459 8075
rect 9674 8072 9680 8084
rect 9447 8044 9680 8072
rect 9447 8041 9459 8044
rect 9401 8035 9459 8041
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 12161 8075 12219 8081
rect 12161 8041 12173 8075
rect 12207 8072 12219 8075
rect 18690 8072 18696 8084
rect 12207 8044 18696 8072
rect 12207 8041 12219 8044
rect 12161 8035 12219 8041
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 18877 8075 18935 8081
rect 18877 8041 18889 8075
rect 18923 8072 18935 8075
rect 20990 8072 20996 8084
rect 18923 8044 20996 8072
rect 18923 8041 18935 8044
rect 18877 8035 18935 8041
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 21177 8075 21235 8081
rect 21177 8041 21189 8075
rect 21223 8072 21235 8075
rect 21450 8072 21456 8084
rect 21223 8044 21456 8072
rect 21223 8041 21235 8044
rect 21177 8035 21235 8041
rect 21450 8032 21456 8044
rect 21508 8032 21514 8084
rect 2869 8007 2927 8013
rect 2869 7973 2881 8007
rect 2915 8004 2927 8007
rect 2958 8004 2964 8016
rect 2915 7976 2964 8004
rect 2915 7973 2927 7976
rect 2869 7967 2927 7973
rect 2958 7964 2964 7976
rect 3016 7964 3022 8016
rect 3326 8004 3332 8016
rect 3287 7976 3332 8004
rect 3326 7964 3332 7976
rect 3384 7964 3390 8016
rect 8573 8007 8631 8013
rect 8573 8004 8585 8007
rect 7576 7976 8585 8004
rect 1670 7896 1676 7948
rect 1728 7936 1734 7948
rect 2041 7939 2099 7945
rect 2041 7936 2053 7939
rect 1728 7908 2053 7936
rect 1728 7896 1734 7908
rect 2041 7905 2053 7908
rect 2087 7905 2099 7939
rect 2041 7899 2099 7905
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2406 7936 2412 7948
rect 2271 7908 2412 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 4985 7939 5043 7945
rect 4985 7905 4997 7939
rect 5031 7905 5043 7939
rect 5166 7936 5172 7948
rect 5127 7908 5172 7936
rect 4985 7899 5043 7905
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 2866 7868 2872 7880
rect 2731 7840 2872 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 2866 7828 2872 7840
rect 2924 7828 2930 7880
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7868 3203 7871
rect 3234 7868 3240 7880
rect 3191 7840 3240 7868
rect 3191 7837 3203 7840
rect 3145 7831 3203 7837
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 3970 7868 3976 7880
rect 3883 7840 3976 7868
rect 3970 7828 3976 7840
rect 4028 7868 4034 7880
rect 4614 7868 4620 7880
rect 4028 7840 4620 7868
rect 4028 7828 4034 7840
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 5000 7800 5028 7899
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 5776 7908 6929 7936
rect 5776 7896 5782 7908
rect 6917 7905 6929 7908
rect 6963 7936 6975 7939
rect 7006 7936 7012 7948
rect 6963 7908 7012 7936
rect 6963 7905 6975 7908
rect 6917 7899 6975 7905
rect 7006 7896 7012 7908
rect 7064 7896 7070 7948
rect 7101 7939 7159 7945
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 7282 7936 7288 7948
rect 7147 7908 7288 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 7576 7945 7604 7976
rect 8573 7973 8585 7976
rect 8619 8004 8631 8007
rect 9766 8004 9772 8016
rect 8619 7976 9772 8004
rect 8619 7973 8631 7976
rect 8573 7967 8631 7973
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 13173 8007 13231 8013
rect 13173 7973 13185 8007
rect 13219 8004 13231 8007
rect 15102 8004 15108 8016
rect 13219 7976 15108 8004
rect 13219 7973 13231 7976
rect 13173 7967 13231 7973
rect 15102 7964 15108 7976
rect 15160 7964 15166 8016
rect 18782 7964 18788 8016
rect 18840 8004 18846 8016
rect 19518 8004 19524 8016
rect 18840 7976 19524 8004
rect 18840 7964 18846 7976
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7905 7619 7939
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7561 7899 7619 7905
rect 7668 7908 7757 7936
rect 5258 7868 5264 7880
rect 5219 7840 5264 7868
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 7374 7868 7380 7880
rect 6052 7840 7380 7868
rect 6052 7828 6058 7840
rect 7374 7828 7380 7840
rect 7432 7868 7438 7880
rect 7668 7868 7696 7908
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 7745 7899 7803 7905
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7905 12587 7939
rect 12710 7936 12716 7948
rect 12671 7908 12716 7936
rect 12529 7899 12587 7905
rect 7834 7868 7840 7880
rect 7432 7840 7696 7868
rect 7795 7840 7840 7868
rect 7432 7828 7438 7840
rect 7834 7828 7840 7840
rect 7892 7868 7898 7880
rect 8294 7868 8300 7880
rect 7892 7840 8300 7868
rect 7892 7828 7898 7840
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 10042 7828 10048 7880
rect 10100 7868 10106 7880
rect 10686 7868 10692 7880
rect 10100 7840 10692 7868
rect 10100 7828 10106 7840
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 10781 7871 10839 7877
rect 10781 7837 10793 7871
rect 10827 7868 10839 7871
rect 11146 7868 11152 7880
rect 10827 7840 11152 7868
rect 10827 7837 10839 7840
rect 10781 7831 10839 7837
rect 11146 7828 11152 7840
rect 11204 7828 11210 7880
rect 7558 7800 7564 7812
rect 5000 7772 7564 7800
rect 7558 7760 7564 7772
rect 7616 7800 7622 7812
rect 10514 7803 10572 7809
rect 10514 7800 10526 7803
rect 7616 7772 10526 7800
rect 7616 7760 7622 7772
rect 10514 7769 10526 7772
rect 10560 7769 10572 7803
rect 12544 7800 12572 7899
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 12802 7868 12808 7880
rect 12763 7840 12808 7868
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 17126 7877 17132 7880
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7868 14703 7871
rect 16853 7871 16911 7877
rect 14691 7840 16160 7868
rect 14691 7837 14703 7840
rect 14645 7831 14703 7837
rect 14274 7800 14280 7812
rect 10514 7763 10572 7769
rect 10612 7772 11275 7800
rect 12544 7772 14280 7800
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 1854 7732 1860 7744
rect 1627 7704 1860 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 1949 7735 2007 7741
rect 1949 7701 1961 7735
rect 1995 7732 2007 7735
rect 2130 7732 2136 7744
rect 1995 7704 2136 7732
rect 1995 7701 2007 7704
rect 1949 7695 2007 7701
rect 2130 7692 2136 7704
rect 2188 7732 2194 7744
rect 4338 7732 4344 7744
rect 2188 7704 4344 7732
rect 2188 7692 2194 7704
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 5629 7735 5687 7741
rect 5629 7701 5641 7735
rect 5675 7732 5687 7735
rect 5810 7732 5816 7744
rect 5675 7704 5816 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 6457 7735 6515 7741
rect 6457 7701 6469 7735
rect 6503 7732 6515 7735
rect 6730 7732 6736 7744
rect 6503 7704 6736 7732
rect 6503 7701 6515 7704
rect 6457 7695 6515 7701
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 6822 7692 6828 7744
rect 6880 7732 6886 7744
rect 8202 7732 8208 7744
rect 6880 7704 6925 7732
rect 8163 7704 8208 7732
rect 6880 7692 6886 7704
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 9674 7692 9680 7744
rect 9732 7732 9738 7744
rect 10612 7732 10640 7772
rect 11146 7732 11152 7744
rect 9732 7704 10640 7732
rect 11107 7704 11152 7732
rect 9732 7692 9738 7704
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11247 7732 11275 7772
rect 14274 7760 14280 7772
rect 14332 7760 14338 7812
rect 14369 7803 14427 7809
rect 14369 7769 14381 7803
rect 14415 7800 14427 7803
rect 14660 7800 14688 7831
rect 16132 7812 16160 7840
rect 16853 7837 16865 7871
rect 16899 7868 16911 7871
rect 17120 7868 17132 7877
rect 16899 7840 16933 7868
rect 17087 7840 17132 7868
rect 16899 7837 16911 7840
rect 16853 7831 16911 7837
rect 17120 7831 17132 7840
rect 16114 7800 16120 7812
rect 14415 7772 14688 7800
rect 16027 7772 16120 7800
rect 14415 7769 14427 7772
rect 14369 7763 14427 7769
rect 11793 7735 11851 7741
rect 11793 7732 11805 7735
rect 11247 7704 11805 7732
rect 11793 7701 11805 7704
rect 11839 7732 11851 7735
rect 13630 7732 13636 7744
rect 11839 7704 13636 7732
rect 11839 7701 11851 7704
rect 11793 7695 11851 7701
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 13725 7735 13783 7741
rect 13725 7701 13737 7735
rect 13771 7732 13783 7735
rect 14384 7732 14412 7763
rect 16114 7760 16120 7772
rect 16172 7800 16178 7812
rect 16485 7803 16543 7809
rect 16485 7800 16497 7803
rect 16172 7772 16497 7800
rect 16172 7760 16178 7772
rect 16485 7769 16497 7772
rect 16531 7800 16543 7803
rect 16868 7800 16896 7831
rect 17126 7828 17132 7831
rect 17184 7828 17190 7880
rect 18690 7868 18696 7880
rect 18651 7840 18696 7868
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 20622 7828 20628 7880
rect 20680 7868 20686 7880
rect 20717 7871 20775 7877
rect 20717 7868 20729 7871
rect 20680 7840 20729 7868
rect 20680 7828 20686 7840
rect 20717 7837 20729 7840
rect 20763 7837 20775 7871
rect 20717 7831 20775 7837
rect 17034 7800 17040 7812
rect 16531 7772 17040 7800
rect 16531 7769 16543 7772
rect 16485 7763 16543 7769
rect 17034 7760 17040 7772
rect 17092 7760 17098 7812
rect 17862 7760 17868 7812
rect 17920 7800 17926 7812
rect 20530 7809 20536 7812
rect 20472 7803 20536 7809
rect 17920 7772 20392 7800
rect 17920 7760 17926 7772
rect 13771 7704 14412 7732
rect 13771 7701 13783 7704
rect 13725 7695 13783 7701
rect 14918 7692 14924 7744
rect 14976 7732 14982 7744
rect 15013 7735 15071 7741
rect 15013 7732 15025 7735
rect 14976 7704 15025 7732
rect 14976 7692 14982 7704
rect 15013 7701 15025 7704
rect 15059 7701 15071 7735
rect 15013 7695 15071 7701
rect 15749 7735 15807 7741
rect 15749 7701 15761 7735
rect 15795 7732 15807 7735
rect 15838 7732 15844 7744
rect 15795 7704 15844 7732
rect 15795 7701 15807 7704
rect 15749 7695 15807 7701
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 17954 7732 17960 7744
rect 16080 7704 17960 7732
rect 16080 7692 16086 7704
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18233 7735 18291 7741
rect 18233 7701 18245 7735
rect 18279 7732 18291 7735
rect 18322 7732 18328 7744
rect 18279 7704 18328 7732
rect 18279 7701 18291 7704
rect 18233 7695 18291 7701
rect 18322 7692 18328 7704
rect 18380 7692 18386 7744
rect 19337 7735 19395 7741
rect 19337 7701 19349 7735
rect 19383 7732 19395 7735
rect 19518 7732 19524 7744
rect 19383 7704 19524 7732
rect 19383 7701 19395 7704
rect 19337 7695 19395 7701
rect 19518 7692 19524 7704
rect 19576 7692 19582 7744
rect 20364 7732 20392 7772
rect 20472 7769 20484 7803
rect 20518 7769 20536 7803
rect 20472 7763 20536 7769
rect 20530 7760 20536 7763
rect 20588 7760 20594 7812
rect 21266 7800 21272 7812
rect 21179 7772 21272 7800
rect 21266 7760 21272 7772
rect 21324 7760 21330 7812
rect 21284 7732 21312 7760
rect 20364 7704 21312 7732
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 658 7488 664 7540
rect 716 7528 722 7540
rect 1118 7528 1124 7540
rect 716 7500 1124 7528
rect 716 7488 722 7500
rect 1118 7488 1124 7500
rect 1176 7488 1182 7540
rect 1854 7528 1860 7540
rect 1815 7500 1860 7528
rect 1854 7488 1860 7500
rect 1912 7488 1918 7540
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2317 7531 2375 7537
rect 2317 7528 2329 7531
rect 2096 7500 2329 7528
rect 2096 7488 2102 7500
rect 2317 7497 2329 7500
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 2648 7500 3985 7528
rect 2648 7488 2654 7500
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 3973 7491 4031 7497
rect 4341 7531 4399 7537
rect 4341 7497 4353 7531
rect 4387 7528 4399 7531
rect 4985 7531 5043 7537
rect 4985 7528 4997 7531
rect 4387 7500 4997 7528
rect 4387 7497 4399 7500
rect 4341 7491 4399 7497
rect 4985 7497 4997 7500
rect 5031 7497 5043 7531
rect 4985 7491 5043 7497
rect 5074 7488 5080 7540
rect 5132 7528 5138 7540
rect 5132 7500 5177 7528
rect 5132 7488 5138 7500
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 6546 7528 6552 7540
rect 5408 7500 6552 7528
rect 5408 7488 5414 7500
rect 6546 7488 6552 7500
rect 6604 7528 6610 7540
rect 6733 7531 6791 7537
rect 6733 7528 6745 7531
rect 6604 7500 6745 7528
rect 6604 7488 6610 7500
rect 6733 7497 6745 7500
rect 6779 7497 6791 7531
rect 9306 7528 9312 7540
rect 9267 7500 9312 7528
rect 6733 7491 6791 7497
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 9398 7488 9404 7540
rect 9456 7528 9462 7540
rect 12158 7528 12164 7540
rect 9456 7500 12164 7528
rect 9456 7488 9462 7500
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 14369 7531 14427 7537
rect 14369 7497 14381 7531
rect 14415 7528 14427 7531
rect 14642 7528 14648 7540
rect 14415 7500 14648 7528
rect 14415 7497 14427 7500
rect 14369 7491 14427 7497
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 17497 7531 17555 7537
rect 17497 7497 17509 7531
rect 17543 7528 17555 7531
rect 17543 7500 18276 7528
rect 17543 7497 17555 7500
rect 17497 7491 17555 7497
rect 2869 7463 2927 7469
rect 2869 7429 2881 7463
rect 2915 7460 2927 7463
rect 7834 7460 7840 7472
rect 2915 7432 5028 7460
rect 2915 7429 2927 7432
rect 2869 7423 2927 7429
rect 5000 7404 5028 7432
rect 5276 7432 7840 7460
rect 934 7352 940 7404
rect 992 7392 998 7404
rect 1118 7392 1124 7404
rect 992 7364 1124 7392
rect 992 7352 998 7364
rect 1118 7352 1124 7364
rect 1176 7352 1182 7404
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 2682 7392 2688 7404
rect 2643 7364 2688 7392
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 3326 7392 3332 7404
rect 3287 7364 3332 7392
rect 3326 7352 3332 7364
rect 3384 7352 3390 7404
rect 4430 7392 4436 7404
rect 3712 7364 4436 7392
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1636 7296 1685 7324
rect 1636 7284 1642 7296
rect 1673 7293 1685 7296
rect 1719 7293 1731 7327
rect 1673 7287 1731 7293
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 3344 7324 3372 7352
rect 3712 7333 3740 7364
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 2924 7296 3372 7324
rect 3697 7327 3755 7333
rect 2924 7284 2930 7296
rect 3697 7293 3709 7327
rect 3743 7293 3755 7327
rect 3878 7324 3884 7336
rect 3839 7296 3884 7324
rect 3697 7287 3755 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 5276 7333 5304 7432
rect 7834 7420 7840 7432
rect 7892 7420 7898 7472
rect 8665 7463 8723 7469
rect 8665 7429 8677 7463
rect 8711 7460 8723 7463
rect 12342 7460 12348 7472
rect 8711 7432 12348 7460
rect 8711 7429 8723 7432
rect 8665 7423 8723 7429
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 14660 7460 14688 7488
rect 14890 7463 14948 7469
rect 14890 7460 14902 7463
rect 14660 7432 14902 7460
rect 14890 7429 14902 7432
rect 14936 7429 14948 7463
rect 14890 7423 14948 7429
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7392 6883 7395
rect 7377 7395 7435 7401
rect 6871 7364 7144 7392
rect 6871 7361 6883 7364
rect 6825 7355 6883 7361
rect 5261 7327 5319 7333
rect 5261 7293 5273 7327
rect 5307 7293 5319 7327
rect 5261 7287 5319 7293
rect 6638 7284 6644 7336
rect 6696 7324 6702 7336
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6696 7296 6929 7324
rect 6696 7284 6702 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 7116 7324 7144 7364
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 8386 7392 8392 7404
rect 7423 7364 8392 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 10433 7395 10491 7401
rect 10433 7361 10445 7395
rect 10479 7392 10491 7395
rect 10594 7392 10600 7404
rect 10479 7364 10600 7392
rect 10479 7361 10491 7364
rect 10433 7355 10491 7361
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 11974 7352 11980 7404
rect 12032 7392 12038 7404
rect 12805 7395 12863 7401
rect 12805 7392 12817 7395
rect 12032 7364 12817 7392
rect 12032 7352 12038 7364
rect 12805 7361 12817 7364
rect 12851 7361 12863 7395
rect 13630 7392 13636 7404
rect 13591 7364 13636 7392
rect 12805 7355 12863 7361
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 14642 7392 14648 7404
rect 14603 7364 14648 7392
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 15746 7392 15752 7404
rect 14752 7364 15752 7392
rect 8297 7327 8355 7333
rect 8297 7324 8309 7327
rect 7116 7296 8309 7324
rect 6917 7287 6975 7293
rect 8297 7293 8309 7296
rect 8343 7324 8355 7327
rect 8570 7324 8576 7336
rect 8343 7296 8576 7324
rect 8343 7293 8355 7296
rect 8297 7287 8355 7293
rect 8570 7284 8576 7296
rect 8628 7324 8634 7336
rect 9306 7324 9312 7336
rect 8628 7296 9312 7324
rect 8628 7284 8634 7296
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 11146 7324 11152 7336
rect 10744 7296 11152 7324
rect 10744 7284 10750 7296
rect 11146 7284 11152 7296
rect 11204 7284 11210 7336
rect 12345 7327 12403 7333
rect 12345 7293 12357 7327
rect 12391 7324 12403 7327
rect 14752 7324 14780 7364
rect 15746 7352 15752 7364
rect 15804 7352 15810 7404
rect 16761 7395 16819 7401
rect 16761 7361 16773 7395
rect 16807 7392 16819 7395
rect 17034 7392 17040 7404
rect 16807 7364 17040 7392
rect 16807 7361 16819 7364
rect 16761 7355 16819 7361
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 17126 7352 17132 7404
rect 17184 7392 17190 7404
rect 18248 7401 18276 7500
rect 20254 7488 20260 7540
rect 20312 7528 20318 7540
rect 20625 7531 20683 7537
rect 20625 7528 20637 7531
rect 20312 7500 20637 7528
rect 20312 7488 20318 7500
rect 20625 7497 20637 7500
rect 20671 7497 20683 7531
rect 20625 7491 20683 7497
rect 20714 7488 20720 7540
rect 20772 7528 20778 7540
rect 21085 7531 21143 7537
rect 21085 7528 21097 7531
rect 20772 7500 21097 7528
rect 20772 7488 20778 7500
rect 21085 7497 21097 7500
rect 21131 7497 21143 7531
rect 21085 7491 21143 7497
rect 18874 7420 18880 7472
rect 18932 7460 18938 7472
rect 20082 7463 20140 7469
rect 20082 7460 20094 7463
rect 18932 7432 20094 7460
rect 18932 7420 18938 7432
rect 20082 7429 20094 7432
rect 20128 7429 20140 7463
rect 20082 7423 20140 7429
rect 20993 7463 21051 7469
rect 20993 7429 21005 7463
rect 21039 7460 21051 7463
rect 21174 7460 21180 7472
rect 21039 7432 21180 7460
rect 21039 7429 21051 7432
rect 20993 7423 21051 7429
rect 17313 7395 17371 7401
rect 17313 7392 17325 7395
rect 17184 7364 17325 7392
rect 17184 7352 17190 7364
rect 17313 7361 17325 7364
rect 17359 7361 17371 7395
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 17313 7355 17371 7361
rect 17889 7364 18153 7392
rect 17144 7324 17172 7352
rect 12391 7296 14780 7324
rect 16049 7296 17172 7324
rect 12391 7293 12403 7296
rect 12345 7287 12403 7293
rect 2590 7216 2596 7268
rect 2648 7256 2654 7268
rect 4617 7259 4675 7265
rect 4617 7256 4629 7259
rect 2648 7228 4629 7256
rect 2648 7216 2654 7228
rect 4617 7225 4629 7228
rect 4663 7225 4675 7259
rect 4617 7219 4675 7225
rect 5997 7259 6055 7265
rect 5997 7225 6009 7259
rect 6043 7256 6055 7259
rect 7190 7256 7196 7268
rect 6043 7228 7196 7256
rect 6043 7225 6055 7228
rect 5997 7219 6055 7225
rect 7190 7216 7196 7228
rect 7248 7216 7254 7268
rect 7561 7259 7619 7265
rect 7561 7225 7573 7259
rect 7607 7256 7619 7259
rect 8386 7256 8392 7268
rect 7607 7228 8392 7256
rect 7607 7225 7619 7228
rect 7561 7219 7619 7225
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 9490 7256 9496 7268
rect 8956 7228 9496 7256
rect 3145 7191 3203 7197
rect 3145 7157 3157 7191
rect 3191 7188 3203 7191
rect 3418 7188 3424 7200
rect 3191 7160 3424 7188
rect 3191 7157 3203 7160
rect 3145 7151 3203 7157
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 6362 7188 6368 7200
rect 6323 7160 6368 7188
rect 6362 7148 6368 7160
rect 6420 7148 6426 7200
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 7929 7191 7987 7197
rect 7929 7188 7941 7191
rect 7064 7160 7941 7188
rect 7064 7148 7070 7160
rect 7929 7157 7941 7160
rect 7975 7188 7987 7191
rect 8956 7188 8984 7228
rect 9490 7216 9496 7228
rect 9548 7216 9554 7268
rect 11057 7259 11115 7265
rect 11057 7225 11069 7259
rect 11103 7256 11115 7259
rect 11164 7256 11192 7284
rect 12618 7256 12624 7268
rect 11103 7228 12020 7256
rect 12579 7228 12624 7256
rect 11103 7225 11115 7228
rect 11057 7219 11115 7225
rect 7975 7160 8984 7188
rect 9033 7191 9091 7197
rect 7975 7157 7987 7160
rect 7929 7151 7987 7157
rect 9033 7157 9045 7191
rect 9079 7188 9091 7191
rect 10778 7188 10784 7200
rect 9079 7160 10784 7188
rect 9079 7157 9091 7160
rect 9033 7151 9091 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11992 7197 12020 7228
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 16049 7256 16077 7296
rect 17218 7284 17224 7336
rect 17276 7324 17282 7336
rect 17889 7324 17917 7364
rect 18141 7361 18153 7364
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7392 18291 7395
rect 21008 7392 21036 7423
rect 21174 7420 21180 7432
rect 21232 7420 21238 7472
rect 18279 7364 21036 7392
rect 18279 7361 18291 7364
rect 18233 7355 18291 7361
rect 18414 7324 18420 7336
rect 17276 7296 17917 7324
rect 18327 7296 18420 7324
rect 17276 7284 17282 7296
rect 18414 7284 18420 7296
rect 18472 7324 18478 7336
rect 18966 7324 18972 7336
rect 18472 7296 18972 7324
rect 18472 7284 18478 7296
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 20349 7327 20407 7333
rect 20349 7293 20361 7327
rect 20395 7324 20407 7327
rect 20622 7324 20628 7336
rect 20395 7296 20628 7324
rect 20395 7293 20407 7296
rect 20349 7287 20407 7293
rect 20622 7284 20628 7296
rect 20680 7284 20686 7336
rect 21266 7324 21272 7336
rect 21227 7296 21272 7324
rect 21266 7284 21272 7296
rect 21324 7284 21330 7336
rect 15948 7228 16077 7256
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 11204 7160 11529 7188
rect 11204 7148 11210 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 11977 7191 12035 7197
rect 11977 7157 11989 7191
rect 12023 7188 12035 7191
rect 12066 7188 12072 7200
rect 12023 7160 12072 7188
rect 12023 7157 12035 7160
rect 11977 7151 12035 7157
rect 12066 7148 12072 7160
rect 12124 7148 12130 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 13173 7191 13231 7197
rect 13173 7188 13185 7191
rect 12492 7160 13185 7188
rect 12492 7148 12498 7160
rect 13173 7157 13185 7160
rect 13219 7188 13231 7191
rect 13446 7188 13452 7200
rect 13219 7160 13452 7188
rect 13219 7157 13231 7160
rect 13173 7151 13231 7157
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 14001 7191 14059 7197
rect 14001 7157 14013 7191
rect 14047 7188 14059 7191
rect 15948 7188 15976 7228
rect 16114 7216 16120 7268
rect 16172 7256 16178 7268
rect 17773 7259 17831 7265
rect 17773 7256 17785 7259
rect 16172 7228 17785 7256
rect 16172 7216 16178 7228
rect 17773 7225 17785 7228
rect 17819 7225 17831 7259
rect 17773 7219 17831 7225
rect 17954 7216 17960 7268
rect 18012 7256 18018 7268
rect 18012 7228 19472 7256
rect 18012 7216 18018 7228
rect 14047 7160 15976 7188
rect 16025 7191 16083 7197
rect 14047 7157 14059 7160
rect 14001 7151 14059 7157
rect 16025 7157 16037 7191
rect 16071 7188 16083 7191
rect 17862 7188 17868 7200
rect 16071 7160 17868 7188
rect 16071 7157 16083 7160
rect 16025 7151 16083 7157
rect 17862 7148 17868 7160
rect 17920 7148 17926 7200
rect 18782 7148 18788 7200
rect 18840 7188 18846 7200
rect 18969 7191 19027 7197
rect 18969 7188 18981 7191
rect 18840 7160 18981 7188
rect 18840 7148 18846 7160
rect 18969 7157 18981 7160
rect 19015 7157 19027 7191
rect 19444 7188 19472 7228
rect 20530 7188 20536 7200
rect 19444 7160 20536 7188
rect 18969 7151 19027 7157
rect 20530 7148 20536 7160
rect 20588 7148 20594 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 1673 6987 1731 6993
rect 1673 6953 1685 6987
rect 1719 6984 1731 6987
rect 1946 6984 1952 6996
rect 1719 6956 1952 6984
rect 1719 6953 1731 6956
rect 1673 6947 1731 6953
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 2682 6944 2688 6996
rect 2740 6984 2746 6996
rect 7374 6984 7380 6996
rect 2740 6956 7144 6984
rect 7335 6956 7380 6984
rect 2740 6944 2746 6956
rect 5350 6916 5356 6928
rect 4448 6888 5356 6916
rect 2314 6848 2320 6860
rect 2275 6820 2320 6848
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 4448 6857 4476 6888
rect 5350 6876 5356 6888
rect 5408 6876 5414 6928
rect 7116 6916 7144 6956
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 9125 6987 9183 6993
rect 9125 6984 9137 6987
rect 7616 6956 9137 6984
rect 7616 6944 7622 6956
rect 9125 6953 9137 6956
rect 9171 6953 9183 6987
rect 9125 6947 9183 6953
rect 9508 6956 10824 6984
rect 9398 6916 9404 6928
rect 6656 6888 7052 6916
rect 7116 6888 9404 6916
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6817 3387 6851
rect 3329 6811 3387 6817
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6817 4491 6851
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 4433 6811 4491 6817
rect 5368 6820 5641 6848
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 2832 6752 3065 6780
rect 2832 6740 2838 6752
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 3344 6780 3372 6811
rect 5368 6780 5396 6820
rect 5629 6817 5641 6820
rect 5675 6848 5687 6851
rect 6656 6848 6684 6888
rect 5675 6820 6684 6848
rect 5675 6817 5687 6820
rect 5629 6811 5687 6817
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 6788 6820 6837 6848
rect 6788 6808 6794 6820
rect 6825 6817 6837 6820
rect 6871 6817 6883 6851
rect 6825 6811 6883 6817
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6817 6975 6851
rect 6917 6811 6975 6817
rect 3344 6752 5396 6780
rect 5445 6783 5503 6789
rect 3053 6743 3111 6749
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 6362 6780 6368 6792
rect 5491 6752 6368 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 6932 6780 6960 6811
rect 6696 6752 6960 6780
rect 7024 6780 7052 6888
rect 9398 6876 9404 6888
rect 9456 6876 9462 6928
rect 7282 6808 7288 6860
rect 7340 6848 7346 6860
rect 8021 6851 8079 6857
rect 8021 6848 8033 6851
rect 7340 6820 8033 6848
rect 7340 6808 7346 6820
rect 8021 6817 8033 6820
rect 8067 6848 8079 6851
rect 8570 6848 8576 6860
rect 8067 6820 8576 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 9508 6848 9536 6956
rect 8720 6820 9536 6848
rect 10505 6851 10563 6857
rect 8720 6808 8726 6820
rect 10505 6817 10517 6851
rect 10551 6848 10563 6851
rect 10686 6848 10692 6860
rect 10551 6820 10692 6848
rect 10551 6817 10563 6820
rect 10505 6811 10563 6817
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 9766 6780 9772 6792
rect 7024 6752 9772 6780
rect 6696 6740 6702 6752
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 10249 6783 10307 6789
rect 10249 6749 10261 6783
rect 10295 6780 10307 6783
rect 10796 6780 10824 6956
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12124 6956 12480 6984
rect 12124 6944 12130 6956
rect 12452 6857 12480 6956
rect 14458 6944 14464 6996
rect 14516 6984 14522 6996
rect 14642 6984 14648 6996
rect 14516 6956 14648 6984
rect 14516 6944 14522 6956
rect 14642 6944 14648 6956
rect 14700 6984 14706 6996
rect 15381 6987 15439 6993
rect 15381 6984 15393 6987
rect 14700 6956 15393 6984
rect 14700 6944 14706 6956
rect 15381 6953 15393 6956
rect 15427 6984 15439 6987
rect 17034 6984 17040 6996
rect 15427 6956 17040 6984
rect 15427 6953 15439 6956
rect 15381 6947 15439 6953
rect 17034 6944 17040 6956
rect 17092 6944 17098 6996
rect 17862 6944 17868 6996
rect 17920 6984 17926 6996
rect 21266 6984 21272 6996
rect 17920 6956 21272 6984
rect 17920 6944 17926 6956
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 16868 6888 17540 6916
rect 12437 6851 12495 6857
rect 12437 6817 12449 6851
rect 12483 6848 12495 6851
rect 12802 6848 12808 6860
rect 12483 6820 12808 6848
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 14274 6808 14280 6860
rect 14332 6848 14338 6860
rect 14369 6851 14427 6857
rect 14369 6848 14381 6851
rect 14332 6820 14381 6848
rect 14332 6808 14338 6820
rect 14369 6817 14381 6820
rect 14415 6848 14427 6851
rect 15562 6848 15568 6860
rect 14415 6820 15568 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 15838 6808 15844 6860
rect 15896 6848 15902 6860
rect 15933 6851 15991 6857
rect 15933 6848 15945 6851
rect 15896 6820 15945 6848
rect 15896 6808 15902 6820
rect 15933 6817 15945 6820
rect 15979 6817 15991 6851
rect 16114 6848 16120 6860
rect 16075 6820 16120 6848
rect 15933 6811 15991 6817
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 16298 6808 16304 6860
rect 16356 6848 16362 6860
rect 16868 6848 16896 6888
rect 17402 6848 17408 6860
rect 16356 6820 16896 6848
rect 16960 6820 17264 6848
rect 17363 6820 17408 6848
rect 16356 6808 16362 6820
rect 10962 6780 10968 6792
rect 10295 6752 10968 6780
rect 10295 6749 10307 6752
rect 10249 6743 10307 6749
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 14645 6783 14703 6789
rect 14645 6780 14657 6783
rect 11112 6752 14657 6780
rect 11112 6740 11118 6752
rect 14645 6749 14657 6752
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 14826 6740 14832 6792
rect 14884 6740 14890 6792
rect 15102 6740 15108 6792
rect 15160 6780 15166 6792
rect 16960 6780 16988 6820
rect 15160 6752 16988 6780
rect 17037 6783 17095 6789
rect 15160 6740 15166 6752
rect 17037 6749 17049 6783
rect 17083 6749 17095 6783
rect 17236 6780 17264 6820
rect 17402 6808 17408 6820
rect 17460 6808 17466 6860
rect 17512 6848 17540 6888
rect 17586 6876 17592 6928
rect 17644 6916 17650 6928
rect 17644 6888 18460 6916
rect 17644 6876 17650 6888
rect 18432 6860 18460 6888
rect 17512 6820 17816 6848
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 17236 6752 17693 6780
rect 17037 6743 17095 6749
rect 17681 6749 17693 6752
rect 17727 6749 17739 6783
rect 17788 6780 17816 6820
rect 18230 6808 18236 6860
rect 18288 6848 18294 6860
rect 18325 6851 18383 6857
rect 18325 6848 18337 6851
rect 18288 6820 18337 6848
rect 18288 6808 18294 6820
rect 18325 6817 18337 6820
rect 18371 6817 18383 6851
rect 18325 6811 18383 6817
rect 18414 6808 18420 6860
rect 18472 6848 18478 6860
rect 18472 6820 19012 6848
rect 18472 6808 18478 6820
rect 18877 6783 18935 6789
rect 18877 6780 18889 6783
rect 17788 6752 18889 6780
rect 17681 6743 17739 6749
rect 18877 6749 18889 6752
rect 18923 6749 18935 6783
rect 18984 6780 19012 6820
rect 20898 6808 20904 6860
rect 20956 6848 20962 6860
rect 21085 6851 21143 6857
rect 21085 6848 21097 6851
rect 20956 6820 21097 6848
rect 20956 6808 20962 6820
rect 21085 6817 21097 6820
rect 21131 6817 21143 6851
rect 21085 6811 21143 6817
rect 20358 6783 20416 6789
rect 20358 6780 20370 6783
rect 18984 6752 20370 6780
rect 18877 6743 18935 6749
rect 20358 6749 20370 6752
rect 20404 6749 20416 6783
rect 20622 6780 20628 6792
rect 20583 6752 20628 6780
rect 20358 6743 20416 6749
rect 2041 6715 2099 6721
rect 2041 6681 2053 6715
rect 2087 6712 2099 6715
rect 3418 6712 3424 6724
rect 2087 6684 3424 6712
rect 2087 6681 2099 6684
rect 2041 6675 2099 6681
rect 3418 6672 3424 6684
rect 3476 6672 3482 6724
rect 4614 6672 4620 6724
rect 4672 6712 4678 6724
rect 4890 6712 4896 6724
rect 4672 6684 4896 6712
rect 4672 6672 4678 6684
rect 4890 6672 4896 6684
rect 4948 6712 4954 6724
rect 6733 6715 6791 6721
rect 4948 6684 6500 6712
rect 4948 6672 4954 6684
rect 2130 6644 2136 6656
rect 2091 6616 2136 6644
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 2682 6644 2688 6656
rect 2643 6616 2688 6644
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 3142 6604 3148 6656
rect 3200 6644 3206 6656
rect 3786 6644 3792 6656
rect 3200 6616 3245 6644
rect 3747 6616 3792 6644
rect 3200 6604 3206 6616
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 4154 6644 4160 6656
rect 4115 6616 4160 6644
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 5074 6644 5080 6656
rect 4304 6616 4349 6644
rect 5035 6616 5080 6644
rect 4304 6604 4310 6616
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 5537 6647 5595 6653
rect 5537 6613 5549 6647
rect 5583 6644 5595 6647
rect 6365 6647 6423 6653
rect 6365 6644 6377 6647
rect 5583 6616 6377 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 6365 6613 6377 6616
rect 6411 6613 6423 6647
rect 6472 6644 6500 6684
rect 6733 6681 6745 6715
rect 6779 6712 6791 6715
rect 7374 6712 7380 6724
rect 6779 6684 7380 6712
rect 6779 6681 6791 6684
rect 6733 6675 6791 6681
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 8573 6715 8631 6721
rect 7484 6684 8340 6712
rect 7484 6644 7512 6684
rect 7742 6644 7748 6656
rect 6472 6616 7512 6644
rect 7703 6616 7748 6644
rect 6365 6607 6423 6613
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 7837 6647 7895 6653
rect 7837 6613 7849 6647
rect 7883 6644 7895 6647
rect 8202 6644 8208 6656
rect 7883 6616 8208 6644
rect 7883 6613 7895 6616
rect 7837 6607 7895 6613
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8312 6644 8340 6684
rect 8573 6681 8585 6715
rect 8619 6712 8631 6715
rect 9858 6712 9864 6724
rect 8619 6684 9864 6712
rect 8619 6681 8631 6684
rect 8573 6675 8631 6681
rect 9858 6672 9864 6684
rect 9916 6672 9922 6724
rect 10069 6684 12112 6712
rect 10069 6644 10097 6684
rect 8312 6616 10097 6644
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 11057 6647 11115 6653
rect 11057 6644 11069 6647
rect 10192 6616 11069 6644
rect 10192 6604 10198 6616
rect 11057 6613 11069 6616
rect 11103 6644 11115 6647
rect 11974 6644 11980 6656
rect 11103 6616 11980 6644
rect 11103 6613 11115 6616
rect 11057 6607 11115 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 12084 6644 12112 6684
rect 12158 6672 12164 6724
rect 12216 6721 12222 6724
rect 12216 6712 12228 6721
rect 12216 6684 12261 6712
rect 12216 6675 12228 6684
rect 12216 6672 12222 6675
rect 12342 6672 12348 6724
rect 12400 6712 12406 6724
rect 14844 6712 14872 6740
rect 12400 6684 14872 6712
rect 12400 6672 12406 6684
rect 15378 6672 15384 6724
rect 15436 6712 15442 6724
rect 17052 6712 17080 6743
rect 20622 6740 20628 6752
rect 20680 6740 20686 6792
rect 17494 6712 17500 6724
rect 15436 6684 17500 6712
rect 15436 6672 15442 6684
rect 17494 6672 17500 6684
rect 17552 6672 17558 6724
rect 19610 6712 19616 6724
rect 18064 6684 19616 6712
rect 12526 6644 12532 6656
rect 12084 6616 12532 6644
rect 12526 6604 12532 6616
rect 12584 6604 12590 6656
rect 12802 6644 12808 6656
rect 12763 6616 12808 6644
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 13078 6644 13084 6656
rect 13039 6616 13084 6644
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 13630 6644 13636 6656
rect 13591 6616 13636 6644
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 14553 6647 14611 6653
rect 14553 6613 14565 6647
rect 14599 6644 14611 6647
rect 14826 6644 14832 6656
rect 14599 6616 14832 6644
rect 14599 6613 14611 6616
rect 14553 6607 14611 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15010 6644 15016 6656
rect 14971 6616 15016 6644
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 16206 6644 16212 6656
rect 16167 6616 16212 6644
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 16574 6644 16580 6656
rect 16535 6616 16580 6644
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6644 16911 6647
rect 16942 6644 16948 6656
rect 16899 6616 16948 6644
rect 16899 6613 16911 6616
rect 16853 6607 16911 6613
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 17586 6604 17592 6656
rect 17644 6644 17650 6656
rect 18064 6653 18092 6684
rect 19610 6672 19616 6684
rect 19668 6672 19674 6724
rect 20530 6672 20536 6724
rect 20588 6712 20594 6724
rect 21269 6715 21327 6721
rect 21269 6712 21281 6715
rect 20588 6684 21281 6712
rect 20588 6672 20594 6684
rect 21269 6681 21281 6684
rect 21315 6681 21327 6715
rect 21269 6675 21327 6681
rect 18049 6647 18107 6653
rect 17644 6616 17689 6644
rect 17644 6604 17650 6616
rect 18049 6613 18061 6647
rect 18095 6613 18107 6647
rect 18690 6644 18696 6656
rect 18651 6616 18696 6644
rect 18049 6607 18107 6613
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 19242 6644 19248 6656
rect 19203 6616 19248 6644
rect 19242 6604 19248 6616
rect 19300 6604 19306 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2685 6443 2743 6449
rect 2685 6440 2697 6443
rect 2188 6412 2697 6440
rect 2188 6400 2194 6412
rect 2685 6409 2697 6412
rect 2731 6409 2743 6443
rect 2685 6403 2743 6409
rect 3053 6443 3111 6449
rect 3053 6409 3065 6443
rect 3099 6440 3111 6443
rect 3142 6440 3148 6452
rect 3099 6412 3148 6440
rect 3099 6409 3111 6412
rect 3053 6403 3111 6409
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3878 6400 3884 6452
rect 3936 6440 3942 6452
rect 3973 6443 4031 6449
rect 3973 6440 3985 6443
rect 3936 6412 3985 6440
rect 3936 6400 3942 6412
rect 3973 6409 3985 6412
rect 4019 6409 4031 6443
rect 3973 6403 4031 6409
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 4982 6440 4988 6452
rect 4387 6412 4988 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 5350 6400 5356 6452
rect 5408 6440 5414 6452
rect 6546 6440 6552 6452
rect 5408 6412 6408 6440
rect 6507 6412 6552 6440
rect 5408 6400 5414 6412
rect 1486 6372 1492 6384
rect 1447 6344 1492 6372
rect 1486 6332 1492 6344
rect 1544 6332 1550 6384
rect 1670 6332 1676 6384
rect 1728 6372 1734 6384
rect 2593 6375 2651 6381
rect 2593 6372 2605 6375
rect 1728 6344 2605 6372
rect 1728 6332 1734 6344
rect 2593 6341 2605 6344
rect 2639 6372 2651 6375
rect 6270 6372 6276 6384
rect 2639 6344 6276 6372
rect 2639 6341 2651 6344
rect 2593 6335 2651 6341
rect 6270 6332 6276 6344
rect 6328 6332 6334 6384
rect 2130 6264 2136 6316
rect 2188 6304 2194 6316
rect 2958 6304 2964 6316
rect 2188 6276 2964 6304
rect 2188 6264 2194 6276
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 4430 6304 4436 6316
rect 4343 6276 4436 6304
rect 4430 6264 4436 6276
rect 4488 6304 4494 6316
rect 4798 6304 4804 6316
rect 4488 6276 4804 6304
rect 4488 6264 4494 6276
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 4982 6304 4988 6316
rect 4943 6276 4988 6304
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 5810 6304 5816 6316
rect 5771 6276 5816 6304
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 6380 6313 6408 6412
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 7098 6440 7104 6452
rect 7059 6412 7104 6440
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6440 8999 6443
rect 8987 6412 9674 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 7558 6332 7564 6384
rect 7616 6372 7622 6384
rect 8110 6372 8116 6384
rect 7616 6344 8116 6372
rect 7616 6332 7622 6344
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 7282 6264 7288 6316
rect 7340 6304 7346 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 7340 6276 7481 6304
rect 7340 6264 7346 6276
rect 7469 6273 7481 6276
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 2547 6208 2581 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 1762 6128 1768 6180
rect 1820 6168 1826 6180
rect 2516 6168 2544 6199
rect 3050 6196 3056 6248
rect 3108 6236 3114 6248
rect 3329 6239 3387 6245
rect 3329 6236 3341 6239
rect 3108 6208 3341 6236
rect 3108 6196 3114 6208
rect 3329 6205 3341 6208
rect 3375 6205 3387 6239
rect 4614 6236 4620 6248
rect 4575 6208 4620 6236
rect 3329 6199 3387 6205
rect 4614 6196 4620 6208
rect 4672 6196 4678 6248
rect 5537 6239 5595 6245
rect 5000 6208 5304 6236
rect 5000 6168 5028 6208
rect 5166 6168 5172 6180
rect 1820 6140 5028 6168
rect 5127 6140 5172 6168
rect 1820 6128 1826 6140
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 5276 6168 5304 6208
rect 5537 6205 5549 6239
rect 5583 6236 5595 6239
rect 7374 6236 7380 6248
rect 5583 6208 7380 6236
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7558 6236 7564 6248
rect 7519 6208 7564 6236
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 7668 6245 7696 6344
rect 8110 6332 8116 6344
rect 8168 6332 8174 6384
rect 9122 6332 9128 6384
rect 9180 6372 9186 6384
rect 9398 6372 9404 6384
rect 9180 6344 9404 6372
rect 9180 6332 9186 6344
rect 9398 6332 9404 6344
rect 9456 6332 9462 6384
rect 9646 6372 9674 6412
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 12066 6440 12072 6452
rect 9824 6412 12072 6440
rect 9824 6400 9830 6412
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 12621 6443 12679 6449
rect 12621 6409 12633 6443
rect 12667 6440 12679 6443
rect 12802 6440 12808 6452
rect 12667 6412 12808 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 12986 6440 12992 6452
rect 12947 6412 12992 6440
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 16761 6443 16819 6449
rect 16761 6440 16773 6443
rect 14608 6412 16773 6440
rect 14608 6400 14614 6412
rect 16761 6409 16773 6412
rect 16807 6409 16819 6443
rect 16761 6403 16819 6409
rect 17218 6400 17224 6452
rect 17276 6440 17282 6452
rect 19797 6443 19855 6449
rect 19797 6440 19809 6443
rect 17276 6412 19809 6440
rect 17276 6400 17282 6412
rect 19797 6409 19809 6412
rect 19843 6440 19855 6443
rect 20898 6440 20904 6452
rect 19843 6412 20904 6440
rect 19843 6409 19855 6412
rect 19797 6403 19855 6409
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 9646 6344 10640 6372
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 10612 6313 10640 6344
rect 11698 6332 11704 6384
rect 11756 6372 11762 6384
rect 14102 6375 14160 6381
rect 14102 6372 14114 6375
rect 11756 6344 14114 6372
rect 11756 6332 11762 6344
rect 14102 6341 14114 6344
rect 14148 6372 14160 6375
rect 14274 6372 14280 6384
rect 14148 6344 14280 6372
rect 14148 6341 14160 6344
rect 14102 6335 14160 6341
rect 14274 6332 14280 6344
rect 14332 6332 14338 6384
rect 15010 6332 15016 6384
rect 15068 6372 15074 6384
rect 15068 6344 16252 6372
rect 15068 6332 15074 6344
rect 10341 6307 10399 6313
rect 10341 6304 10353 6307
rect 8628 6276 10353 6304
rect 8628 6264 8634 6276
rect 10341 6273 10353 6276
rect 10387 6304 10399 6307
rect 10597 6307 10655 6313
rect 10387 6276 10548 6304
rect 10387 6273 10399 6276
rect 10341 6267 10399 6273
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6205 7711 6239
rect 10520 6236 10548 6276
rect 10597 6273 10609 6307
rect 10643 6304 10655 6307
rect 10962 6304 10968 6316
rect 10643 6276 10968 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 10962 6264 10968 6276
rect 11020 6304 11026 6316
rect 11609 6307 11667 6313
rect 11609 6304 11621 6307
rect 11020 6276 11621 6304
rect 11020 6264 11026 6276
rect 11609 6273 11621 6276
rect 11655 6304 11667 6307
rect 12802 6304 12808 6316
rect 11655 6276 12808 6304
rect 11655 6273 11667 6276
rect 11609 6267 11667 6273
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 14369 6307 14427 6313
rect 14369 6273 14381 6307
rect 14415 6304 14427 6307
rect 14458 6304 14464 6316
rect 14415 6276 14464 6304
rect 14415 6273 14427 6276
rect 14369 6267 14427 6273
rect 14458 6264 14464 6276
rect 14516 6264 14522 6316
rect 16022 6264 16028 6316
rect 16080 6313 16086 6316
rect 16080 6304 16092 6313
rect 16080 6276 16125 6304
rect 16080 6267 16092 6276
rect 16080 6264 16086 6267
rect 11238 6236 11244 6248
rect 10520 6208 11244 6236
rect 7653 6199 7711 6205
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 16224 6236 16252 6344
rect 17034 6332 17040 6384
rect 17092 6372 17098 6384
rect 20622 6372 20628 6384
rect 17092 6344 20628 6372
rect 17092 6332 17098 6344
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 17052 6304 17080 6332
rect 17586 6304 17592 6316
rect 16347 6276 17080 6304
rect 17144 6276 17592 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 17144 6236 17172 6276
rect 17586 6264 17592 6276
rect 17644 6264 17650 6316
rect 17862 6264 17868 6316
rect 17920 6313 17926 6316
rect 17920 6304 17932 6313
rect 17920 6276 17965 6304
rect 17920 6267 17932 6276
rect 17920 6264 17926 6267
rect 18046 6264 18052 6316
rect 18104 6264 18110 6316
rect 18156 6313 18184 6344
rect 20622 6332 20628 6344
rect 20680 6332 20686 6384
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6273 18199 6307
rect 18506 6304 18512 6316
rect 18467 6276 18512 6304
rect 18141 6267 18199 6273
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19153 6307 19211 6313
rect 19153 6304 19165 6307
rect 19024 6276 19165 6304
rect 19024 6264 19030 6276
rect 19153 6273 19165 6276
rect 19199 6273 19211 6307
rect 19889 6307 19947 6313
rect 19889 6304 19901 6307
rect 19153 6267 19211 6273
rect 19260 6276 19901 6304
rect 16224 6208 17172 6236
rect 18064 6236 18092 6264
rect 19260 6236 19288 6276
rect 19889 6273 19901 6276
rect 19935 6273 19947 6307
rect 19889 6267 19947 6273
rect 19978 6264 19984 6316
rect 20036 6304 20042 6316
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20036 6276 20821 6304
rect 20036 6264 20042 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 19610 6236 19616 6248
rect 18064 6208 19288 6236
rect 19571 6208 19616 6236
rect 19610 6196 19616 6208
rect 19668 6196 19674 6248
rect 20533 6239 20591 6245
rect 20533 6236 20545 6239
rect 19720 6208 20545 6236
rect 5997 6171 6055 6177
rect 5276 6140 5764 6168
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 2041 6103 2099 6109
rect 2041 6069 2053 6103
rect 2087 6100 2099 6103
rect 3142 6100 3148 6112
rect 2087 6072 3148 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 3142 6060 3148 6072
rect 3200 6100 3206 6112
rect 5350 6100 5356 6112
rect 3200 6072 5356 6100
rect 3200 6060 3206 6072
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 5736 6100 5764 6140
rect 5997 6137 6009 6171
rect 6043 6168 6055 6171
rect 6822 6168 6828 6180
rect 6043 6140 6828 6168
rect 6043 6137 6055 6140
rect 5997 6131 6055 6137
rect 6822 6128 6828 6140
rect 6880 6128 6886 6180
rect 6932 6140 9260 6168
rect 6730 6100 6736 6112
rect 5736 6072 6736 6100
rect 6730 6060 6736 6072
rect 6788 6100 6794 6112
rect 6932 6100 6960 6140
rect 8570 6100 8576 6112
rect 6788 6072 6960 6100
rect 8531 6072 8576 6100
rect 6788 6060 6794 6072
rect 8570 6060 8576 6072
rect 8628 6060 8634 6112
rect 9232 6109 9260 6140
rect 18598 6128 18604 6180
rect 18656 6168 18662 6180
rect 18656 6140 19564 6168
rect 18656 6128 18662 6140
rect 9217 6103 9275 6109
rect 9217 6069 9229 6103
rect 9263 6100 9275 6103
rect 10686 6100 10692 6112
rect 9263 6072 10692 6100
rect 9263 6069 9275 6072
rect 9217 6063 9275 6069
rect 10686 6060 10692 6072
rect 10744 6060 10750 6112
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11238 6100 11244 6112
rect 11112 6072 11244 6100
rect 11112 6060 11118 6072
rect 11238 6060 11244 6072
rect 11296 6060 11302 6112
rect 12250 6100 12256 6112
rect 12211 6072 12256 6100
rect 12250 6060 12256 6072
rect 12308 6060 12314 6112
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 14921 6103 14979 6109
rect 14921 6100 14933 6103
rect 13044 6072 14933 6100
rect 13044 6060 13050 6072
rect 14921 6069 14933 6072
rect 14967 6069 14979 6103
rect 14921 6063 14979 6069
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 18966 6100 18972 6112
rect 18739 6072 18972 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 19061 6103 19119 6109
rect 19061 6069 19073 6103
rect 19107 6100 19119 6103
rect 19242 6100 19248 6112
rect 19107 6072 19248 6100
rect 19107 6069 19119 6072
rect 19061 6063 19119 6069
rect 19242 6060 19248 6072
rect 19300 6060 19306 6112
rect 19536 6100 19564 6140
rect 19720 6100 19748 6208
rect 20533 6205 20545 6208
rect 20579 6236 20591 6239
rect 20714 6236 20720 6248
rect 20579 6208 20720 6236
rect 20579 6205 20591 6208
rect 20533 6199 20591 6205
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 19536 6072 19748 6100
rect 19886 6060 19892 6112
rect 19944 6100 19950 6112
rect 20257 6103 20315 6109
rect 20257 6100 20269 6103
rect 19944 6072 20269 6100
rect 19944 6060 19950 6072
rect 20257 6069 20269 6072
rect 20303 6069 20315 6103
rect 20257 6063 20315 6069
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2498 5896 2504 5908
rect 2455 5868 2504 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 4154 5896 4160 5908
rect 3467 5868 4160 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 4154 5856 4160 5868
rect 4212 5856 4218 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5592 5868 6316 5896
rect 5592 5856 5598 5868
rect 14 5788 20 5840
rect 72 5828 78 5840
rect 934 5828 940 5840
rect 72 5800 940 5828
rect 72 5788 78 5800
rect 934 5788 940 5800
rect 992 5788 998 5840
rect 5074 5828 5080 5840
rect 1964 5800 5080 5828
rect 1854 5760 1860 5772
rect 1815 5732 1860 5760
rect 1854 5720 1860 5732
rect 1912 5720 1918 5772
rect 1964 5769 1992 5800
rect 5074 5788 5080 5800
rect 5132 5788 5138 5840
rect 5166 5788 5172 5840
rect 5224 5828 5230 5840
rect 5626 5828 5632 5840
rect 5224 5800 5632 5828
rect 5224 5788 5230 5800
rect 5626 5788 5632 5800
rect 5684 5828 5690 5840
rect 5721 5831 5779 5837
rect 5721 5828 5733 5831
rect 5684 5800 5733 5828
rect 5684 5788 5690 5800
rect 5721 5797 5733 5800
rect 5767 5797 5779 5831
rect 5721 5791 5779 5797
rect 6181 5831 6239 5837
rect 6181 5797 6193 5831
rect 6227 5797 6239 5831
rect 6288 5828 6316 5868
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 9122 5896 9128 5908
rect 8628 5868 9128 5896
rect 8628 5856 8634 5868
rect 9122 5856 9128 5868
rect 9180 5896 9186 5908
rect 9674 5896 9680 5908
rect 9180 5868 9680 5896
rect 9180 5856 9186 5868
rect 9674 5856 9680 5868
rect 9732 5856 9738 5908
rect 12345 5899 12403 5905
rect 12345 5865 12357 5899
rect 12391 5896 12403 5899
rect 12526 5896 12532 5908
rect 12391 5868 12532 5896
rect 12391 5865 12403 5868
rect 12345 5859 12403 5865
rect 12526 5856 12532 5868
rect 12584 5896 12590 5908
rect 13262 5896 13268 5908
rect 12584 5868 13268 5896
rect 12584 5856 12590 5868
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 14185 5899 14243 5905
rect 14185 5865 14197 5899
rect 14231 5896 14243 5899
rect 14274 5896 14280 5908
rect 14231 5868 14280 5896
rect 14231 5865 14243 5868
rect 14185 5859 14243 5865
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 16301 5899 16359 5905
rect 16301 5865 16313 5899
rect 16347 5896 16359 5899
rect 17218 5896 17224 5908
rect 16347 5868 17224 5896
rect 16347 5865 16359 5868
rect 16301 5859 16359 5865
rect 17218 5856 17224 5868
rect 17276 5856 17282 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 19334 5896 19340 5908
rect 17460 5868 19340 5896
rect 17460 5856 17466 5868
rect 19334 5856 19340 5868
rect 19392 5856 19398 5908
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 19576 5868 19932 5896
rect 19576 5856 19582 5868
rect 7101 5831 7159 5837
rect 7101 5828 7113 5831
rect 6288 5800 7113 5828
rect 6181 5791 6239 5797
rect 7101 5797 7113 5800
rect 7147 5797 7159 5831
rect 7101 5791 7159 5797
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5729 2007 5763
rect 2774 5760 2780 5772
rect 2735 5732 2780 5760
rect 1949 5723 2007 5729
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 2958 5720 2964 5772
rect 3016 5760 3022 5772
rect 4798 5760 4804 5772
rect 3016 5732 4568 5760
rect 4759 5732 4804 5760
rect 3016 5720 3022 5732
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2682 5692 2688 5704
rect 2087 5664 2688 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 3050 5692 3056 5704
rect 3011 5664 3056 5692
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3418 5652 3424 5704
rect 3476 5692 3482 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3476 5664 3801 5692
rect 3476 5652 3482 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 4338 5692 4344 5704
rect 3789 5655 3847 5661
rect 3896 5664 4344 5692
rect 2498 5584 2504 5636
rect 2556 5624 2562 5636
rect 3896 5624 3924 5664
rect 4338 5652 4344 5664
rect 4396 5692 4402 5704
rect 4433 5695 4491 5701
rect 4433 5692 4445 5695
rect 4396 5664 4445 5692
rect 4396 5652 4402 5664
rect 4433 5661 4445 5664
rect 4479 5661 4491 5695
rect 4540 5692 4568 5732
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 6196 5760 6224 5791
rect 15654 5788 15660 5840
rect 15712 5828 15718 5840
rect 15712 5800 16988 5828
rect 15712 5788 15718 5800
rect 4908 5732 6224 5760
rect 4908 5692 4936 5732
rect 8202 5720 8208 5772
rect 8260 5760 8266 5772
rect 8570 5760 8576 5772
rect 8260 5732 8576 5760
rect 8260 5720 8266 5732
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 10502 5760 10508 5772
rect 10459 5732 10508 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 10502 5720 10508 5732
rect 10560 5760 10566 5772
rect 10962 5760 10968 5772
rect 10560 5732 10968 5760
rect 10560 5720 10566 5732
rect 10962 5720 10968 5732
rect 11020 5720 11026 5772
rect 12802 5760 12808 5772
rect 12715 5732 12808 5760
rect 12802 5720 12808 5732
rect 12860 5760 12866 5772
rect 13265 5763 13323 5769
rect 13265 5760 13277 5763
rect 12860 5732 13277 5760
rect 12860 5720 12866 5732
rect 13265 5729 13277 5732
rect 13311 5760 13323 5763
rect 14458 5760 14464 5772
rect 13311 5732 14464 5760
rect 13311 5729 13323 5732
rect 13265 5723 13323 5729
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 16850 5760 16856 5772
rect 15948 5732 16856 5760
rect 4540 5664 4936 5692
rect 4433 5655 4491 5661
rect 5442 5652 5448 5704
rect 5500 5692 5506 5704
rect 5500 5664 5856 5692
rect 5500 5652 5506 5664
rect 5828 5636 5856 5664
rect 5902 5652 5908 5704
rect 5960 5692 5966 5704
rect 6362 5692 6368 5704
rect 5960 5664 6005 5692
rect 6323 5664 6368 5692
rect 5960 5652 5966 5664
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 6696 5664 6837 5692
rect 6696 5652 6702 5664
rect 6825 5661 6837 5664
rect 6871 5692 6883 5695
rect 6914 5692 6920 5704
rect 6871 5664 6920 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 7190 5652 7196 5704
rect 7248 5692 7254 5704
rect 7285 5695 7343 5701
rect 7285 5692 7297 5695
rect 7248 5664 7297 5692
rect 7248 5652 7254 5664
rect 7285 5661 7297 5664
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 7892 5664 7941 5692
rect 7892 5652 7898 5664
rect 7929 5661 7941 5664
rect 7975 5692 7987 5695
rect 8297 5695 8355 5701
rect 8297 5692 8309 5695
rect 7975 5664 8309 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8297 5661 8309 5664
rect 8343 5692 8355 5695
rect 9030 5692 9036 5704
rect 8343 5664 9036 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 14728 5695 14786 5701
rect 14728 5692 14740 5695
rect 14660 5664 14740 5692
rect 5077 5627 5135 5633
rect 5077 5624 5089 5627
rect 2556 5596 3924 5624
rect 3988 5596 5089 5624
rect 2556 5584 2562 5596
rect 3988 5565 4016 5596
rect 5077 5593 5089 5596
rect 5123 5593 5135 5627
rect 5077 5587 5135 5593
rect 5810 5584 5816 5636
rect 5868 5624 5874 5636
rect 5868 5596 9076 5624
rect 5868 5584 5874 5596
rect 3973 5559 4031 5565
rect 3973 5525 3985 5559
rect 4019 5525 4031 5559
rect 3973 5519 4031 5525
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4249 5559 4307 5565
rect 4249 5556 4261 5559
rect 4120 5528 4261 5556
rect 4120 5516 4126 5528
rect 4249 5525 4261 5528
rect 4295 5525 4307 5559
rect 4249 5519 4307 5525
rect 4985 5559 5043 5565
rect 4985 5525 4997 5559
rect 5031 5556 5043 5559
rect 5258 5556 5264 5568
rect 5031 5528 5264 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 5442 5556 5448 5568
rect 5403 5528 5448 5556
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 6270 5516 6276 5568
rect 6328 5556 6334 5568
rect 9048 5565 9076 5596
rect 9858 5584 9864 5636
rect 9916 5624 9922 5636
rect 10042 5624 10048 5636
rect 9916 5596 10048 5624
rect 9916 5584 9922 5596
rect 10042 5584 10048 5596
rect 10100 5584 10106 5636
rect 10168 5627 10226 5633
rect 10168 5593 10180 5627
rect 10214 5624 10226 5627
rect 11054 5624 11060 5636
rect 10214 5596 11060 5624
rect 10214 5593 10226 5596
rect 10168 5587 10226 5593
rect 11054 5584 11060 5596
rect 11112 5584 11118 5636
rect 11232 5627 11290 5633
rect 11232 5624 11244 5627
rect 11164 5596 11244 5624
rect 6641 5559 6699 5565
rect 6641 5556 6653 5559
rect 6328 5528 6653 5556
rect 6328 5516 6334 5528
rect 6641 5525 6653 5528
rect 6687 5525 6699 5559
rect 6641 5519 6699 5525
rect 9033 5559 9091 5565
rect 9033 5525 9045 5559
rect 9079 5556 9091 5559
rect 11164 5556 11192 5596
rect 11232 5593 11244 5596
rect 11278 5593 11290 5627
rect 11232 5587 11290 5593
rect 11698 5584 11704 5636
rect 11756 5624 11762 5636
rect 14660 5624 14688 5664
rect 14728 5661 14740 5664
rect 14774 5692 14786 5695
rect 15948 5692 15976 5732
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 16960 5704 16988 5800
rect 19150 5788 19156 5840
rect 19208 5828 19214 5840
rect 19794 5828 19800 5840
rect 19208 5800 19800 5828
rect 19208 5788 19214 5800
rect 19794 5788 19800 5800
rect 19852 5788 19858 5840
rect 17034 5720 17040 5772
rect 17092 5760 17098 5772
rect 17092 5732 17137 5760
rect 17092 5720 17098 5732
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 19705 5763 19763 5769
rect 18196 5732 18920 5760
rect 18196 5720 18202 5732
rect 18892 5704 18920 5732
rect 19705 5729 19717 5763
rect 19751 5760 19763 5763
rect 19904 5760 19932 5868
rect 20162 5856 20168 5908
rect 20220 5896 20226 5908
rect 20533 5899 20591 5905
rect 20533 5896 20545 5899
rect 20220 5868 20545 5896
rect 20220 5856 20226 5868
rect 20533 5865 20545 5868
rect 20579 5865 20591 5899
rect 20533 5859 20591 5865
rect 20257 5831 20315 5837
rect 20257 5797 20269 5831
rect 20303 5828 20315 5831
rect 20346 5828 20352 5840
rect 20303 5800 20352 5828
rect 20303 5797 20315 5800
rect 20257 5791 20315 5797
rect 20346 5788 20352 5800
rect 20404 5788 20410 5840
rect 20530 5760 20536 5772
rect 19751 5732 20536 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 20530 5720 20536 5732
rect 20588 5720 20594 5772
rect 21177 5763 21235 5769
rect 21177 5729 21189 5763
rect 21223 5760 21235 5763
rect 21266 5760 21272 5772
rect 21223 5732 21272 5760
rect 21223 5729 21235 5732
rect 21177 5723 21235 5729
rect 21266 5720 21272 5732
rect 21324 5720 21330 5772
rect 16114 5692 16120 5704
rect 14774 5664 15976 5692
rect 16075 5664 16120 5692
rect 14774 5661 14786 5664
rect 14728 5655 14786 5661
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 16577 5695 16635 5701
rect 16577 5661 16589 5695
rect 16623 5661 16635 5695
rect 16942 5692 16948 5704
rect 16855 5664 16948 5692
rect 16577 5655 16635 5661
rect 11756 5596 14688 5624
rect 16592 5624 16620 5655
rect 16942 5652 16948 5664
rect 17000 5692 17006 5704
rect 17293 5695 17351 5701
rect 17293 5692 17305 5695
rect 17000 5664 17305 5692
rect 17000 5652 17006 5664
rect 17293 5661 17305 5664
rect 17339 5661 17351 5695
rect 17293 5655 17351 5661
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 19886 5692 19892 5704
rect 18932 5664 19025 5692
rect 19847 5664 19892 5692
rect 18932 5652 18938 5664
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 20993 5695 21051 5701
rect 20993 5661 21005 5695
rect 21039 5692 21051 5695
rect 21542 5692 21548 5704
rect 21039 5664 21548 5692
rect 21039 5661 21051 5664
rect 20993 5655 21051 5661
rect 21542 5652 21548 5664
rect 21600 5652 21606 5704
rect 16592 5596 18664 5624
rect 11756 5584 11762 5596
rect 9079 5528 11192 5556
rect 9079 5525 9091 5528
rect 9033 5519 9091 5525
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12710 5556 12716 5568
rect 12032 5528 12716 5556
rect 12032 5516 12038 5528
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 13722 5556 13728 5568
rect 13683 5528 13728 5556
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 15562 5516 15568 5568
rect 15620 5556 15626 5568
rect 15841 5559 15899 5565
rect 15841 5556 15853 5559
rect 15620 5528 15853 5556
rect 15620 5516 15626 5528
rect 15841 5525 15853 5528
rect 15887 5556 15899 5559
rect 15930 5556 15936 5568
rect 15887 5528 15936 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 16761 5559 16819 5565
rect 16761 5525 16773 5559
rect 16807 5556 16819 5559
rect 17862 5556 17868 5568
rect 16807 5528 17868 5556
rect 16807 5525 16819 5528
rect 16761 5519 16819 5525
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18417 5559 18475 5565
rect 18417 5556 18429 5559
rect 18012 5528 18429 5556
rect 18012 5516 18018 5528
rect 18417 5525 18429 5528
rect 18463 5525 18475 5559
rect 18636 5556 18664 5596
rect 19242 5584 19248 5636
rect 19300 5624 19306 5636
rect 19978 5624 19984 5636
rect 19300 5596 19984 5624
rect 19300 5584 19306 5596
rect 19978 5584 19984 5596
rect 20036 5584 20042 5636
rect 20898 5624 20904 5636
rect 20859 5596 20904 5624
rect 20898 5584 20904 5596
rect 20956 5584 20962 5636
rect 18693 5559 18751 5565
rect 18693 5556 18705 5559
rect 18636 5528 18705 5556
rect 18417 5519 18475 5525
rect 18693 5525 18705 5528
rect 18739 5525 18751 5559
rect 19794 5556 19800 5568
rect 19755 5528 19800 5556
rect 18693 5519 18751 5525
rect 19794 5516 19800 5528
rect 19852 5516 19858 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 2501 5355 2559 5361
rect 2501 5321 2513 5355
rect 2547 5352 2559 5355
rect 3145 5355 3203 5361
rect 3145 5352 3157 5355
rect 2547 5324 3157 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 3145 5321 3157 5324
rect 3191 5321 3203 5355
rect 3145 5315 3203 5321
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4982 5352 4988 5364
rect 4295 5324 4988 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 5629 5355 5687 5361
rect 5629 5321 5641 5355
rect 5675 5352 5687 5355
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 5675 5324 6469 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 7469 5355 7527 5361
rect 7469 5352 7481 5355
rect 6871 5324 7481 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 7469 5321 7481 5324
rect 7515 5321 7527 5355
rect 7469 5315 7527 5321
rect 7837 5355 7895 5361
rect 7837 5321 7849 5355
rect 7883 5352 7895 5355
rect 8018 5352 8024 5364
rect 7883 5324 8024 5352
rect 7883 5321 7895 5324
rect 7837 5315 7895 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 9125 5355 9183 5361
rect 9125 5352 9137 5355
rect 9088 5324 9137 5352
rect 9088 5312 9094 5324
rect 9125 5321 9137 5324
rect 9171 5352 9183 5355
rect 9582 5352 9588 5364
rect 9171 5324 9588 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 10962 5312 10968 5364
rect 11020 5352 11026 5364
rect 13909 5355 13967 5361
rect 11020 5324 13492 5352
rect 11020 5312 11026 5324
rect 934 5244 940 5296
rect 992 5284 998 5296
rect 1489 5287 1547 5293
rect 1489 5284 1501 5287
rect 992 5256 1501 5284
rect 992 5244 998 5256
rect 1489 5253 1501 5256
rect 1535 5253 1547 5287
rect 1670 5284 1676 5296
rect 1631 5256 1676 5284
rect 1489 5247 1547 5253
rect 1670 5244 1676 5256
rect 1728 5244 1734 5296
rect 2593 5287 2651 5293
rect 2593 5253 2605 5287
rect 2639 5284 2651 5287
rect 2639 5256 4292 5284
rect 2639 5253 2651 5256
rect 2593 5247 2651 5253
rect 3326 5216 3332 5228
rect 3287 5188 3332 5216
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 3418 5176 3424 5228
rect 3476 5216 3482 5228
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3476 5188 4077 5216
rect 3476 5176 3482 5188
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4264 5216 4292 5256
rect 4338 5244 4344 5296
rect 4396 5284 4402 5296
rect 4396 5256 10364 5284
rect 4396 5244 4402 5256
rect 4430 5216 4436 5228
rect 4264 5188 4436 5216
rect 4065 5179 4123 5185
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5216 5595 5219
rect 5902 5216 5908 5228
rect 5583 5188 5908 5216
rect 5583 5185 5595 5188
rect 5537 5179 5595 5185
rect 2682 5148 2688 5160
rect 2643 5120 2688 5148
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 3234 5108 3240 5160
rect 3292 5148 3298 5160
rect 3605 5151 3663 5157
rect 3605 5148 3617 5151
rect 3292 5120 3617 5148
rect 3292 5108 3298 5120
rect 3605 5117 3617 5120
rect 3651 5117 3663 5151
rect 4540 5148 4568 5179
rect 5902 5176 5908 5188
rect 5960 5176 5966 5228
rect 8478 5216 8484 5228
rect 8439 5188 8484 5216
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 9490 5176 9496 5228
rect 9548 5216 9554 5228
rect 10238 5219 10296 5225
rect 10238 5216 10250 5219
rect 9548 5188 10250 5216
rect 9548 5176 9554 5188
rect 10238 5185 10250 5188
rect 10284 5185 10296 5219
rect 10336 5216 10364 5256
rect 11790 5244 11796 5296
rect 11848 5284 11854 5296
rect 12342 5284 12348 5296
rect 11848 5256 12348 5284
rect 11848 5244 11854 5256
rect 12342 5244 12348 5256
rect 12400 5244 12406 5296
rect 10336 5188 10456 5216
rect 10238 5179 10296 5185
rect 5810 5148 5816 5160
rect 3605 5111 3663 5117
rect 3712 5120 4568 5148
rect 5771 5120 5816 5148
rect 842 5040 848 5092
rect 900 5080 906 5092
rect 3326 5080 3332 5092
rect 900 5052 3332 5080
rect 900 5040 906 5052
rect 3326 5040 3332 5052
rect 3384 5080 3390 5092
rect 3712 5080 3740 5120
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 6917 5151 6975 5157
rect 6917 5148 6929 5151
rect 5920 5120 6929 5148
rect 3384 5052 3740 5080
rect 3384 5040 3390 5052
rect 3878 5040 3884 5092
rect 3936 5080 3942 5092
rect 3936 5052 4844 5080
rect 3936 5040 3942 5052
rect 106 4972 112 5024
rect 164 5012 170 5024
rect 934 5012 940 5024
rect 164 4984 940 5012
rect 164 4972 170 4984
rect 934 4972 940 4984
rect 992 4972 998 5024
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 3786 4972 3792 5024
rect 3844 5012 3850 5024
rect 3970 5012 3976 5024
rect 3844 4984 3976 5012
rect 3844 4972 3850 4984
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 4816 5012 4844 5052
rect 4890 5040 4896 5092
rect 4948 5080 4954 5092
rect 5920 5080 5948 5120
rect 6917 5117 6929 5120
rect 6963 5117 6975 5151
rect 6917 5111 6975 5117
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 7116 5080 7144 5111
rect 7650 5108 7656 5160
rect 7708 5148 7714 5160
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7708 5120 7941 5148
rect 7708 5108 7714 5120
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 8110 5148 8116 5160
rect 8071 5120 8116 5148
rect 7929 5111 7987 5117
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 10428 5148 10456 5188
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 10560 5188 10793 5216
rect 10560 5176 10566 5188
rect 10781 5185 10793 5188
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 12066 5176 12072 5228
rect 12124 5216 12130 5228
rect 13274 5219 13332 5225
rect 13274 5216 13286 5219
rect 12124 5188 13286 5216
rect 12124 5176 12130 5188
rect 13274 5185 13286 5188
rect 13320 5185 13332 5219
rect 13274 5179 13332 5185
rect 11790 5148 11796 5160
rect 10428 5120 11796 5148
rect 11790 5108 11796 5120
rect 11848 5108 11854 5160
rect 13464 5148 13492 5324
rect 13909 5321 13921 5355
rect 13955 5352 13967 5355
rect 14458 5352 14464 5364
rect 13955 5324 14464 5352
rect 13955 5321 13967 5324
rect 13909 5315 13967 5321
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5216 13599 5219
rect 13924 5216 13952 5315
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 15841 5355 15899 5361
rect 15841 5321 15853 5355
rect 15887 5352 15899 5355
rect 16298 5352 16304 5364
rect 15887 5324 16304 5352
rect 15887 5321 15899 5324
rect 15841 5315 15899 5321
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17402 5352 17408 5364
rect 17184 5324 17408 5352
rect 17184 5312 17190 5324
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17586 5352 17592 5364
rect 17547 5324 17592 5352
rect 17586 5312 17592 5324
rect 17644 5312 17650 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 19150 5352 19156 5364
rect 18012 5324 19156 5352
rect 18012 5312 18018 5324
rect 19150 5312 19156 5324
rect 19208 5312 19214 5364
rect 19334 5352 19340 5364
rect 19295 5324 19340 5352
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 19702 5312 19708 5364
rect 19760 5352 19766 5364
rect 20530 5352 20536 5364
rect 19760 5324 20536 5352
rect 19760 5312 19766 5324
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 16206 5284 16212 5296
rect 13587 5188 13952 5216
rect 14016 5256 16212 5284
rect 13587 5185 13599 5188
rect 13541 5179 13599 5185
rect 14016 5148 14044 5256
rect 16206 5244 16212 5256
rect 16264 5244 16270 5296
rect 20162 5284 20168 5296
rect 16868 5256 20168 5284
rect 14277 5219 14335 5225
rect 14277 5185 14289 5219
rect 14323 5185 14335 5219
rect 14918 5216 14924 5228
rect 14879 5188 14924 5216
rect 14277 5179 14335 5185
rect 13464 5120 14044 5148
rect 14292 5148 14320 5179
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 14292 5120 14872 5148
rect 4948 5052 5948 5080
rect 6288 5052 8800 5080
rect 4948 5040 4954 5052
rect 5169 5015 5227 5021
rect 5169 5012 5181 5015
rect 4816 4984 5181 5012
rect 5169 4981 5181 4984
rect 5215 4981 5227 5015
rect 5169 4975 5227 4981
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 6288 5012 6316 5052
rect 5592 4984 6316 5012
rect 5592 4972 5598 4984
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 8018 5012 8024 5024
rect 6972 4984 8024 5012
rect 6972 4972 6978 4984
rect 8018 4972 8024 4984
rect 8076 4972 8082 5024
rect 8662 5012 8668 5024
rect 8623 4984 8668 5012
rect 8662 4972 8668 4984
rect 8720 4972 8726 5024
rect 8772 5012 8800 5052
rect 9306 5040 9312 5092
rect 9364 5080 9370 5092
rect 9490 5080 9496 5092
rect 9364 5052 9496 5080
rect 9364 5040 9370 5052
rect 9490 5040 9496 5052
rect 9548 5040 9554 5092
rect 12158 5080 12164 5092
rect 12119 5052 12164 5080
rect 12158 5040 12164 5052
rect 12216 5040 12222 5092
rect 13630 5040 13636 5092
rect 13688 5080 13694 5092
rect 14292 5080 14320 5120
rect 14458 5080 14464 5092
rect 13688 5052 14320 5080
rect 14419 5052 14464 5080
rect 13688 5040 13694 5052
rect 14458 5040 14464 5052
rect 14516 5040 14522 5092
rect 11054 5012 11060 5024
rect 8772 4984 11060 5012
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 14550 4972 14556 5024
rect 14608 5012 14614 5024
rect 14737 5015 14795 5021
rect 14737 5012 14749 5015
rect 14608 4984 14749 5012
rect 14608 4972 14614 4984
rect 14737 4981 14749 4984
rect 14783 4981 14795 5015
rect 14844 5012 14872 5120
rect 15212 5080 15240 5179
rect 15672 5148 15700 5179
rect 15746 5176 15752 5228
rect 15804 5216 15810 5228
rect 16117 5219 16175 5225
rect 16117 5216 16129 5219
rect 15804 5188 16129 5216
rect 15804 5176 15810 5188
rect 16117 5185 16129 5188
rect 16163 5216 16175 5219
rect 16298 5216 16304 5228
rect 16163 5188 16304 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 16868 5148 16896 5256
rect 20162 5244 20168 5256
rect 20220 5244 20226 5296
rect 20254 5244 20260 5296
rect 20312 5284 20318 5296
rect 20622 5284 20628 5296
rect 20312 5256 20628 5284
rect 20312 5244 20318 5256
rect 20622 5244 20628 5256
rect 20680 5284 20686 5296
rect 21269 5287 21327 5293
rect 20680 5256 20760 5284
rect 20680 5244 20686 5256
rect 17126 5216 17132 5228
rect 17087 5188 17132 5216
rect 17126 5176 17132 5188
rect 17184 5176 17190 5228
rect 17221 5220 17279 5225
rect 17310 5220 17316 5228
rect 17221 5219 17316 5220
rect 17221 5185 17233 5219
rect 17267 5192 17316 5219
rect 17267 5185 17279 5192
rect 17221 5179 17279 5185
rect 17310 5176 17316 5192
rect 17368 5176 17374 5228
rect 17770 5176 17776 5228
rect 17828 5216 17834 5228
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 17828 5188 17877 5216
rect 17828 5176 17834 5188
rect 17865 5185 17877 5188
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 18417 5219 18475 5225
rect 18417 5216 18429 5219
rect 18196 5188 18429 5216
rect 18196 5176 18202 5188
rect 18417 5185 18429 5188
rect 18463 5185 18475 5219
rect 19058 5216 19064 5228
rect 19019 5188 19064 5216
rect 18417 5179 18475 5185
rect 19058 5176 19064 5188
rect 19116 5216 19122 5228
rect 19886 5216 19892 5228
rect 19116 5188 19892 5216
rect 19116 5176 19122 5188
rect 19886 5176 19892 5188
rect 19944 5176 19950 5228
rect 19978 5176 19984 5228
rect 20036 5216 20042 5228
rect 20732 5225 20760 5256
rect 21269 5253 21281 5287
rect 21315 5284 21327 5287
rect 21358 5284 21364 5296
rect 21315 5256 21364 5284
rect 21315 5253 21327 5256
rect 21269 5247 21327 5253
rect 21358 5244 21364 5256
rect 21416 5244 21422 5296
rect 20450 5219 20508 5225
rect 20450 5216 20462 5219
rect 20036 5188 20462 5216
rect 20036 5176 20042 5188
rect 20450 5185 20462 5188
rect 20496 5185 20508 5219
rect 20450 5179 20508 5185
rect 20717 5219 20775 5225
rect 20717 5185 20729 5219
rect 20763 5185 20775 5219
rect 20717 5179 20775 5185
rect 15672 5120 16896 5148
rect 17037 5151 17095 5157
rect 17037 5117 17049 5151
rect 17083 5148 17095 5151
rect 19702 5148 19708 5160
rect 17083 5120 19708 5148
rect 17083 5117 17095 5120
rect 17037 5111 17095 5117
rect 19702 5108 19708 5120
rect 19760 5108 19766 5160
rect 18877 5083 18935 5089
rect 18877 5080 18889 5083
rect 15212 5052 18889 5080
rect 18877 5049 18889 5052
rect 18923 5049 18935 5083
rect 21082 5080 21088 5092
rect 21043 5052 21088 5080
rect 18877 5043 18935 5049
rect 21082 5040 21088 5052
rect 21140 5040 21146 5092
rect 15194 5012 15200 5024
rect 14844 4984 15200 5012
rect 14737 4975 14795 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15378 5012 15384 5024
rect 15339 4984 15384 5012
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 17954 5012 17960 5024
rect 16347 4984 17960 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 17954 4972 17960 4984
rect 18012 4972 18018 5024
rect 18049 5015 18107 5021
rect 18049 4981 18061 5015
rect 18095 5012 18107 5015
rect 18506 5012 18512 5024
rect 18095 4984 18512 5012
rect 18095 4981 18107 4984
rect 18049 4975 18107 4981
rect 18506 4972 18512 4984
rect 18564 4972 18570 5024
rect 18601 5015 18659 5021
rect 18601 4981 18613 5015
rect 18647 5012 18659 5015
rect 20070 5012 20076 5024
rect 18647 4984 20076 5012
rect 18647 4981 18659 4984
rect 18601 4975 18659 4981
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 4890 4808 4896 4820
rect 2832 4780 4752 4808
rect 4851 4780 4896 4808
rect 2832 4768 2838 4780
rect 3786 4740 3792 4752
rect 2240 4712 3792 4740
rect 1394 4632 1400 4684
rect 1452 4672 1458 4684
rect 1949 4675 2007 4681
rect 1949 4672 1961 4675
rect 1452 4644 1961 4672
rect 1452 4632 1458 4644
rect 1949 4641 1961 4644
rect 1995 4641 2007 4675
rect 1949 4635 2007 4641
rect 2240 4616 2268 4712
rect 3786 4700 3792 4712
rect 3844 4700 3850 4752
rect 4724 4740 4752 4780
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5902 4808 5908 4820
rect 5863 4780 5908 4808
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 7650 4808 7656 4820
rect 6012 4780 7656 4808
rect 4982 4740 4988 4752
rect 4724 4712 4988 4740
rect 4982 4700 4988 4712
rect 5040 4700 5046 4752
rect 5534 4740 5540 4752
rect 5276 4712 5540 4740
rect 2314 4632 2320 4684
rect 2372 4672 2378 4684
rect 2593 4675 2651 4681
rect 2593 4672 2605 4675
rect 2372 4644 2605 4672
rect 2372 4632 2378 4644
rect 2593 4641 2605 4644
rect 2639 4672 2651 4675
rect 2682 4672 2688 4684
rect 2639 4644 2688 4672
rect 2639 4641 2651 4644
rect 2593 4635 2651 4641
rect 2682 4632 2688 4644
rect 2740 4672 2746 4684
rect 4249 4675 4307 4681
rect 2740 4632 2774 4672
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4798 4672 4804 4684
rect 4295 4644 4804 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 5276 4681 5304 4712
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 5261 4675 5319 4681
rect 5261 4641 5273 4675
rect 5307 4641 5319 4675
rect 5442 4672 5448 4684
rect 5403 4644 5448 4672
rect 5261 4635 5319 4641
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 2222 4604 2228 4616
rect 2183 4576 2228 4604
rect 2222 4564 2228 4576
rect 2280 4564 2286 4616
rect 2746 4604 2774 4632
rect 4338 4604 4344 4616
rect 2746 4576 4344 4604
rect 4338 4564 4344 4576
rect 4396 4564 4402 4616
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4614 4604 4620 4616
rect 4479 4576 4620 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 6012 4604 6040 4780
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 7929 4811 7987 4817
rect 7929 4808 7941 4811
rect 7800 4780 7941 4808
rect 7800 4768 7806 4780
rect 7929 4777 7941 4780
rect 7975 4777 7987 4811
rect 7929 4771 7987 4777
rect 7944 4740 7972 4771
rect 8110 4768 8116 4820
rect 8168 4808 8174 4820
rect 8478 4808 8484 4820
rect 8168 4780 8484 4808
rect 8168 4768 8174 4780
rect 8478 4768 8484 4780
rect 8536 4808 8542 4820
rect 9858 4808 9864 4820
rect 8536 4780 9864 4808
rect 8536 4768 8542 4780
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10502 4808 10508 4820
rect 10463 4780 10508 4808
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 10781 4811 10839 4817
rect 10781 4808 10793 4811
rect 10652 4780 10793 4808
rect 10652 4768 10658 4780
rect 10781 4777 10793 4780
rect 10827 4777 10839 4811
rect 11238 4808 11244 4820
rect 11199 4780 11244 4808
rect 10781 4771 10839 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 12860 4780 12909 4808
rect 12860 4768 12866 4780
rect 12897 4777 12909 4780
rect 12943 4777 12955 4811
rect 12897 4771 12955 4777
rect 17126 4768 17132 4820
rect 17184 4808 17190 4820
rect 20257 4811 20315 4817
rect 20257 4808 20269 4811
rect 17184 4780 20269 4808
rect 17184 4768 17190 4780
rect 20257 4777 20269 4780
rect 20303 4777 20315 4811
rect 20257 4771 20315 4777
rect 9677 4743 9735 4749
rect 7944 4712 9352 4740
rect 6454 4632 6460 4684
rect 6512 4672 6518 4684
rect 6549 4675 6607 4681
rect 6549 4672 6561 4675
rect 6512 4644 6561 4672
rect 6512 4632 6518 4644
rect 6549 4641 6561 4644
rect 6595 4641 6607 4675
rect 6549 4635 6607 4641
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 8018 4672 8024 4684
rect 7432 4644 8024 4672
rect 7432 4632 7438 4644
rect 8018 4632 8024 4644
rect 8076 4672 8082 4684
rect 9122 4672 9128 4684
rect 8076 4644 8340 4672
rect 9083 4644 9128 4672
rect 8076 4632 8082 4644
rect 4764 4576 6040 4604
rect 6273 4607 6331 4613
rect 4764 4564 4770 4576
rect 6273 4573 6285 4607
rect 6319 4604 6331 4607
rect 6472 4604 6500 4632
rect 6319 4576 6500 4604
rect 7285 4607 7343 4613
rect 6319 4573 6331 4576
rect 6273 4567 6331 4573
rect 7285 4573 7297 4607
rect 7331 4604 7343 4607
rect 7466 4604 7472 4616
rect 7331 4576 7472 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 7742 4604 7748 4616
rect 7703 4576 7748 4604
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 8312 4600 8340 4644
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 9324 4613 9352 4712
rect 9677 4709 9689 4743
rect 9723 4740 9735 4743
rect 10962 4740 10968 4752
rect 9723 4712 10968 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 10410 4632 10416 4684
rect 10468 4672 10474 4684
rect 10594 4672 10600 4684
rect 10468 4644 10600 4672
rect 10468 4632 10474 4644
rect 10594 4632 10600 4644
rect 10652 4672 10658 4684
rect 12621 4675 12679 4681
rect 10652 4644 11468 4672
rect 10652 4632 10658 4644
rect 8389 4607 8447 4613
rect 8389 4600 8401 4607
rect 8312 4573 8401 4600
rect 8435 4573 8447 4607
rect 8312 4572 8447 4573
rect 8389 4567 8447 4572
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 9953 4607 10011 4613
rect 9953 4573 9965 4607
rect 9999 4573 10011 4607
rect 9953 4567 10011 4573
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4604 11023 4607
rect 11146 4604 11152 4616
rect 11011 4576 11152 4604
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 3418 4536 3424 4548
rect 2832 4508 2877 4536
rect 3068 4508 3424 4536
rect 2832 4496 2838 4508
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 3068 4468 3096 4508
rect 3418 4496 3424 4508
rect 3476 4536 3482 4548
rect 3881 4539 3939 4545
rect 3476 4508 3832 4536
rect 3476 4496 3482 4508
rect 2915 4440 3096 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 3142 4428 3148 4480
rect 3200 4468 3206 4480
rect 3237 4471 3295 4477
rect 3237 4468 3249 4471
rect 3200 4440 3249 4468
rect 3200 4428 3206 4440
rect 3237 4437 3249 4440
rect 3283 4437 3295 4471
rect 3804 4468 3832 4508
rect 3881 4505 3893 4539
rect 3927 4536 3939 4539
rect 7760 4536 7788 4564
rect 3927 4508 7788 4536
rect 3927 4505 3939 4508
rect 3881 4499 3939 4505
rect 8110 4496 8116 4548
rect 8168 4536 8174 4548
rect 9968 4536 9996 4567
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 8168 4508 9996 4536
rect 11440 4536 11468 4644
rect 12621 4641 12633 4675
rect 12667 4672 12679 4675
rect 12820 4672 12848 4768
rect 16117 4743 16175 4749
rect 16117 4709 16129 4743
rect 16163 4709 16175 4743
rect 16117 4703 16175 4709
rect 16577 4743 16635 4749
rect 16577 4709 16589 4743
rect 16623 4740 16635 4743
rect 17770 4740 17776 4752
rect 16623 4712 17776 4740
rect 16623 4709 16635 4712
rect 16577 4703 16635 4709
rect 13262 4672 13268 4684
rect 12667 4644 13268 4672
rect 12667 4641 12679 4644
rect 12621 4635 12679 4641
rect 13262 4632 13268 4644
rect 13320 4672 13326 4684
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 13320 4644 14105 4672
rect 13320 4632 13326 4644
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 16132 4672 16160 4703
rect 17770 4700 17776 4712
rect 17828 4700 17834 4752
rect 19337 4743 19395 4749
rect 19337 4709 19349 4743
rect 19383 4740 19395 4743
rect 19610 4740 19616 4752
rect 19383 4712 19616 4740
rect 19383 4709 19395 4712
rect 19337 4703 19395 4709
rect 19610 4700 19616 4712
rect 19668 4700 19674 4752
rect 19886 4700 19892 4752
rect 19944 4740 19950 4752
rect 20162 4740 20168 4752
rect 19944 4712 20168 4740
rect 19944 4700 19950 4712
rect 20162 4700 20168 4712
rect 20220 4740 20226 4752
rect 21269 4743 21327 4749
rect 21269 4740 21281 4743
rect 20220 4712 21281 4740
rect 20220 4700 20226 4712
rect 21269 4709 21281 4712
rect 21315 4709 21327 4743
rect 21269 4703 21327 4709
rect 17126 4672 17132 4684
rect 16132 4644 17132 4672
rect 14093 4635 14151 4641
rect 11790 4564 11796 4616
rect 11848 4604 11854 4616
rect 13170 4604 13176 4616
rect 11848 4576 13176 4604
rect 11848 4564 11854 4576
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 13722 4604 13728 4616
rect 13587 4576 13728 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 14108 4604 14136 4635
rect 17126 4632 17132 4644
rect 17184 4632 17190 4684
rect 18877 4675 18935 4681
rect 18877 4641 18889 4675
rect 18923 4672 18935 4675
rect 20254 4672 20260 4684
rect 18923 4644 20260 4672
rect 18923 4641 18935 4644
rect 18877 4635 18935 4641
rect 20254 4632 20260 4644
rect 20312 4632 20318 4684
rect 20806 4672 20812 4684
rect 20767 4644 20812 4672
rect 20806 4632 20812 4644
rect 20864 4632 20870 4684
rect 14734 4604 14740 4616
rect 14108 4576 14740 4604
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 15930 4604 15936 4616
rect 15891 4576 15936 4604
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 16850 4604 16856 4616
rect 16439 4576 16856 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4604 17003 4607
rect 17218 4604 17224 4616
rect 16991 4576 17224 4604
rect 16991 4573 17003 4576
rect 16945 4567 17003 4573
rect 17218 4564 17224 4576
rect 17276 4564 17282 4616
rect 18138 4564 18144 4616
rect 18196 4604 18202 4616
rect 18621 4607 18679 4613
rect 18621 4604 18633 4607
rect 18196 4576 18633 4604
rect 18196 4564 18202 4576
rect 18621 4573 18633 4576
rect 18667 4604 18679 4607
rect 18782 4604 18788 4616
rect 18667 4576 18788 4604
rect 18667 4573 18679 4576
rect 18621 4567 18679 4573
rect 18782 4564 18788 4576
rect 18840 4564 18846 4616
rect 19150 4564 19156 4616
rect 19208 4604 19214 4616
rect 19613 4607 19671 4613
rect 19613 4604 19625 4607
rect 19208 4576 19625 4604
rect 19208 4564 19214 4576
rect 19613 4573 19625 4576
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 20070 4564 20076 4616
rect 20128 4604 20134 4616
rect 20717 4607 20775 4613
rect 20717 4604 20729 4607
rect 20128 4576 20729 4604
rect 20128 4564 20134 4576
rect 20717 4573 20729 4576
rect 20763 4573 20775 4607
rect 20717 4567 20775 4573
rect 12354 4539 12412 4545
rect 12354 4536 12366 4539
rect 11440 4508 12366 4536
rect 8168 4496 8174 4508
rect 12354 4505 12366 4508
rect 12400 4505 12412 4539
rect 13188 4536 13216 4564
rect 14338 4539 14396 4545
rect 14338 4536 14350 4539
rect 13188 4508 14350 4536
rect 12354 4499 12412 4505
rect 14338 4505 14350 4508
rect 14384 4505 14396 4539
rect 14338 4499 14396 4505
rect 15378 4496 15384 4548
rect 15436 4536 15442 4548
rect 18874 4536 18880 4548
rect 15436 4508 18880 4536
rect 15436 4496 15442 4508
rect 18874 4496 18880 4508
rect 18932 4496 18938 4548
rect 19058 4496 19064 4548
rect 19116 4536 19122 4548
rect 19702 4536 19708 4548
rect 19116 4508 19708 4536
rect 19116 4496 19122 4508
rect 19702 4496 19708 4508
rect 19760 4496 19766 4548
rect 3970 4468 3976 4480
rect 3804 4440 3976 4468
rect 3237 4431 3295 4437
rect 3970 4428 3976 4440
rect 4028 4428 4034 4480
rect 4525 4471 4583 4477
rect 4525 4437 4537 4471
rect 4571 4468 4583 4471
rect 4614 4468 4620 4480
rect 4571 4440 4620 4468
rect 4571 4437 4583 4440
rect 4525 4431 4583 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 5534 4468 5540 4480
rect 5495 4440 5540 4468
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 7469 4471 7527 4477
rect 7469 4437 7481 4471
rect 7515 4468 7527 4471
rect 7558 4468 7564 4480
rect 7515 4440 7564 4468
rect 7515 4437 7527 4440
rect 7469 4431 7527 4437
rect 7558 4428 7564 4440
rect 7616 4428 7622 4480
rect 8202 4468 8208 4480
rect 8163 4440 8208 4468
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 9122 4428 9128 4480
rect 9180 4468 9186 4480
rect 9217 4471 9275 4477
rect 9217 4468 9229 4471
rect 9180 4440 9229 4468
rect 9180 4428 9186 4440
rect 9217 4437 9229 4440
rect 9263 4437 9275 4471
rect 9217 4431 9275 4437
rect 10137 4471 10195 4477
rect 10137 4437 10149 4471
rect 10183 4468 10195 4471
rect 13170 4468 13176 4480
rect 10183 4440 13176 4468
rect 10183 4437 10195 4440
rect 10137 4431 10195 4437
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 13725 4471 13783 4477
rect 13725 4437 13737 4471
rect 13771 4468 13783 4471
rect 14918 4468 14924 4480
rect 13771 4440 14924 4468
rect 13771 4437 13783 4440
rect 13725 4431 13783 4437
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15473 4471 15531 4477
rect 15473 4468 15485 4471
rect 15160 4440 15485 4468
rect 15160 4428 15166 4440
rect 15473 4437 15485 4440
rect 15519 4437 15531 4471
rect 15473 4431 15531 4437
rect 17129 4471 17187 4477
rect 17129 4437 17141 4471
rect 17175 4468 17187 4471
rect 17218 4468 17224 4480
rect 17175 4440 17224 4468
rect 17175 4437 17187 4440
rect 17129 4431 17187 4437
rect 17218 4428 17224 4440
rect 17276 4428 17282 4480
rect 17494 4468 17500 4480
rect 17455 4440 17500 4468
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 19150 4468 19156 4480
rect 17736 4440 19156 4468
rect 17736 4428 17742 4440
rect 19150 4428 19156 4440
rect 19208 4428 19214 4480
rect 19518 4428 19524 4480
rect 19576 4468 19582 4480
rect 19797 4471 19855 4477
rect 19797 4468 19809 4471
rect 19576 4440 19809 4468
rect 19576 4428 19582 4440
rect 19797 4437 19809 4440
rect 19843 4437 19855 4471
rect 20622 4468 20628 4480
rect 20583 4440 20628 4468
rect 19797 4431 19855 4437
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 1670 4224 1676 4276
rect 1728 4264 1734 4276
rect 1765 4267 1823 4273
rect 1765 4264 1777 4267
rect 1728 4236 1777 4264
rect 1728 4224 1734 4236
rect 1765 4233 1777 4236
rect 1811 4233 1823 4267
rect 1765 4227 1823 4233
rect 1857 4267 1915 4273
rect 1857 4233 1869 4267
rect 1903 4264 1915 4267
rect 3234 4264 3240 4276
rect 1903 4236 3240 4264
rect 1903 4233 1915 4236
rect 1857 4227 1915 4233
rect 3234 4224 3240 4236
rect 3292 4224 3298 4276
rect 4617 4267 4675 4273
rect 4617 4233 4629 4267
rect 4663 4233 4675 4267
rect 5994 4264 6000 4276
rect 5955 4236 6000 4264
rect 4617 4227 4675 4233
rect 4632 4196 4660 4227
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 7466 4224 7472 4276
rect 7524 4224 7530 4276
rect 8110 4264 8116 4276
rect 8071 4236 8116 4264
rect 8110 4224 8116 4236
rect 8168 4224 8174 4276
rect 9766 4264 9772 4276
rect 8220 4236 9772 4264
rect 7484 4196 7512 4224
rect 4632 4168 7512 4196
rect 7558 4156 7564 4208
rect 7616 4196 7622 4208
rect 8220 4196 8248 4236
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 10594 4224 10600 4276
rect 10652 4264 10658 4276
rect 10689 4267 10747 4273
rect 10689 4264 10701 4267
rect 10652 4236 10701 4264
rect 10652 4224 10658 4236
rect 10689 4233 10701 4236
rect 10735 4233 10747 4267
rect 10689 4227 10747 4233
rect 11054 4224 11060 4276
rect 11112 4264 11118 4276
rect 11701 4267 11759 4273
rect 11701 4264 11713 4267
rect 11112 4236 11713 4264
rect 11112 4224 11118 4236
rect 11701 4233 11713 4236
rect 11747 4233 11759 4267
rect 11701 4227 11759 4233
rect 15930 4224 15936 4276
rect 15988 4264 15994 4276
rect 16117 4267 16175 4273
rect 16117 4264 16129 4267
rect 15988 4236 16129 4264
rect 15988 4224 15994 4236
rect 16117 4233 16129 4236
rect 16163 4233 16175 4267
rect 16117 4227 16175 4233
rect 18874 4224 18880 4276
rect 18932 4264 18938 4276
rect 19058 4264 19064 4276
rect 18932 4236 19064 4264
rect 18932 4224 18938 4236
rect 19058 4224 19064 4236
rect 19116 4224 19122 4276
rect 10502 4196 10508 4208
rect 7616 4168 8248 4196
rect 9324 4168 10508 4196
rect 7616 4156 7622 4168
rect 2314 4128 2320 4140
rect 1688 4100 2320 4128
rect 1688 4069 1716 4100
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2866 4128 2872 4140
rect 2827 4100 2872 4128
rect 2866 4088 2872 4100
rect 2924 4088 2930 4140
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3252 4100 3893 4128
rect 1673 4063 1731 4069
rect 1673 4029 1685 4063
rect 1719 4029 1731 4063
rect 1673 4023 1731 4029
rect 2593 4063 2651 4069
rect 2593 4029 2605 4063
rect 2639 4029 2651 4063
rect 2593 4023 2651 4029
rect 2608 3992 2636 4023
rect 2682 4020 2688 4072
rect 2740 4060 2746 4072
rect 2777 4063 2835 4069
rect 2777 4060 2789 4063
rect 2740 4032 2789 4060
rect 2740 4020 2746 4032
rect 2777 4029 2789 4032
rect 2823 4029 2835 4063
rect 2777 4023 2835 4029
rect 3050 3992 3056 4004
rect 2608 3964 3056 3992
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 3252 4001 3280 4100
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 3881 4091 3939 4097
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4128 4491 4131
rect 4614 4128 4620 4140
rect 4479 4100 4620 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 4893 4131 4951 4137
rect 4893 4097 4905 4131
rect 4939 4097 4951 4131
rect 4893 4091 4951 4097
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4128 5411 4131
rect 5626 4128 5632 4140
rect 5399 4100 5632 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 4908 4060 4936 4091
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 5718 4060 5724 4072
rect 4908 4032 5724 4060
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 5828 4060 5856 4091
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 5960 4100 7021 4128
rect 5960 4088 5966 4100
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 7466 4128 7472 4140
rect 7427 4100 7472 4128
rect 7009 4091 7067 4097
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 7926 4128 7932 4140
rect 7887 4100 7932 4128
rect 7926 4088 7932 4100
rect 7984 4088 7990 4140
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4097 8631 4131
rect 8573 4091 8631 4097
rect 5994 4060 6000 4072
rect 5828 4032 6000 4060
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6546 4060 6552 4072
rect 6507 4032 6552 4060
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 8588 4060 8616 4091
rect 8662 4088 8668 4140
rect 8720 4128 8726 4140
rect 9324 4137 9352 4168
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 13538 4156 13544 4208
rect 13596 4205 13602 4208
rect 13596 4199 13660 4205
rect 13596 4165 13614 4199
rect 13648 4165 13660 4199
rect 13596 4159 13660 4165
rect 13596 4156 13602 4159
rect 15194 4156 15200 4208
rect 15252 4196 15258 4208
rect 18598 4196 18604 4208
rect 15252 4168 18604 4196
rect 15252 4156 15258 4168
rect 18598 4156 18604 4168
rect 18656 4156 18662 4208
rect 20806 4196 20812 4208
rect 19352 4168 19656 4196
rect 20767 4168 20812 4196
rect 9582 4137 9588 4140
rect 8849 4131 8907 4137
rect 8849 4128 8861 4131
rect 8720 4100 8861 4128
rect 8720 4088 8726 4100
rect 8849 4097 8861 4100
rect 8895 4097 8907 4131
rect 8849 4091 8907 4097
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 9576 4091 9588 4137
rect 9640 4128 9646 4140
rect 9640 4100 9676 4128
rect 9582 4088 9588 4091
rect 9640 4088 9646 4100
rect 9858 4088 9864 4140
rect 9916 4128 9922 4140
rect 12825 4131 12883 4137
rect 12825 4128 12837 4131
rect 9916 4100 12837 4128
rect 9916 4088 9922 4100
rect 12825 4097 12837 4100
rect 12871 4128 12883 4131
rect 12986 4128 12992 4140
rect 12871 4100 12992 4128
rect 12871 4097 12883 4100
rect 12825 4091 12883 4097
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 13081 4131 13139 4137
rect 13081 4097 13093 4131
rect 13127 4128 13139 4131
rect 13262 4128 13268 4140
rect 13127 4100 13268 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 13262 4088 13268 4100
rect 13320 4128 13326 4140
rect 13357 4131 13415 4137
rect 13357 4128 13369 4131
rect 13320 4100 13369 4128
rect 13320 4088 13326 4100
rect 13357 4097 13369 4100
rect 13403 4097 13415 4131
rect 13357 4091 13415 4097
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 15013 4131 15071 4137
rect 15013 4128 15025 4131
rect 14424 4100 15025 4128
rect 14424 4088 14430 4100
rect 15013 4097 15025 4100
rect 15059 4097 15071 4131
rect 15470 4128 15476 4140
rect 15431 4100 15476 4128
rect 15013 4091 15071 4097
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 15930 4128 15936 4140
rect 15891 4100 15936 4128
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 17034 4128 17040 4140
rect 16995 4100 17040 4128
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 18049 4131 18107 4137
rect 18049 4097 18061 4131
rect 18095 4128 18107 4131
rect 18690 4128 18696 4140
rect 18095 4100 18696 4128
rect 18095 4097 18107 4100
rect 18049 4091 18107 4097
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 18966 4088 18972 4140
rect 19024 4128 19030 4140
rect 19352 4128 19380 4168
rect 19024 4100 19380 4128
rect 19024 4088 19030 4100
rect 19426 4088 19432 4140
rect 19484 4137 19490 4140
rect 19484 4128 19496 4137
rect 19628 4128 19656 4168
rect 20806 4156 20812 4168
rect 20864 4156 20870 4208
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 19484 4100 19529 4128
rect 19628 4100 20177 4128
rect 19484 4091 19496 4100
rect 20165 4097 20177 4100
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 19484 4088 19490 4091
rect 20438 4088 20444 4140
rect 20496 4128 20502 4140
rect 20901 4131 20959 4137
rect 20901 4128 20913 4131
rect 20496 4100 20913 4128
rect 20496 4088 20502 4100
rect 20901 4097 20913 4100
rect 20947 4097 20959 4131
rect 20901 4091 20959 4097
rect 9122 4060 9128 4072
rect 7116 4032 9128 4060
rect 3237 3995 3295 4001
rect 3237 3961 3249 3995
rect 3283 3961 3295 3995
rect 3237 3955 3295 3961
rect 3605 3995 3663 4001
rect 3605 3961 3617 3995
rect 3651 3992 3663 3995
rect 5537 3995 5595 4001
rect 3651 3964 5488 3992
rect 3651 3961 3663 3964
rect 3605 3955 3663 3961
rect 2038 3884 2044 3936
rect 2096 3924 2102 3936
rect 2225 3927 2283 3933
rect 2225 3924 2237 3927
rect 2096 3896 2237 3924
rect 2096 3884 2102 3896
rect 2225 3893 2237 3896
rect 2271 3893 2283 3927
rect 4062 3924 4068 3936
rect 4023 3896 4068 3924
rect 2225 3887 2283 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 5074 3924 5080 3936
rect 5035 3896 5080 3924
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5460 3924 5488 3964
rect 5537 3961 5549 3995
rect 5583 3992 5595 3995
rect 6086 3992 6092 4004
rect 5583 3964 6092 3992
rect 5583 3961 5595 3964
rect 5537 3955 5595 3961
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 7116 3924 7144 4032
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 15838 4060 15844 4072
rect 14752 4032 15844 4060
rect 7193 3995 7251 4001
rect 7193 3961 7205 3995
rect 7239 3992 7251 3995
rect 7558 3992 7564 4004
rect 7239 3964 7564 3992
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 7558 3952 7564 3964
rect 7616 3952 7622 4004
rect 8294 3952 8300 4004
rect 8352 3992 8358 4004
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 8352 3964 8401 3992
rect 8352 3952 8358 3964
rect 8389 3961 8401 3964
rect 8435 3961 8447 3995
rect 8389 3955 8447 3961
rect 10410 3952 10416 4004
rect 10468 3992 10474 4004
rect 14752 4001 14780 4032
rect 15838 4020 15844 4032
rect 15896 4020 15902 4072
rect 17129 4063 17187 4069
rect 17129 4029 17141 4063
rect 17175 4029 17187 4063
rect 17129 4023 17187 4029
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4060 17371 4063
rect 17494 4060 17500 4072
rect 17359 4032 17500 4060
rect 17359 4029 17371 4032
rect 17313 4023 17371 4029
rect 14737 3995 14795 4001
rect 10468 3964 11836 3992
rect 10468 3952 10474 3964
rect 7650 3924 7656 3936
rect 5460 3896 7144 3924
rect 7611 3896 7656 3924
rect 7650 3884 7656 3896
rect 7708 3884 7714 3936
rect 9033 3927 9091 3933
rect 9033 3893 9045 3927
rect 9079 3924 9091 3927
rect 10594 3924 10600 3936
rect 9079 3896 10600 3924
rect 9079 3893 9091 3896
rect 9033 3887 9091 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11149 3927 11207 3933
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 11606 3924 11612 3936
rect 11195 3896 11612 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 11808 3924 11836 3964
rect 14737 3961 14749 3995
rect 14783 3961 14795 3995
rect 14737 3955 14795 3961
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 16669 3995 16727 4001
rect 16669 3992 16681 3995
rect 14884 3964 16681 3992
rect 14884 3952 14890 3964
rect 16669 3961 16681 3964
rect 16715 3961 16727 3995
rect 17144 3992 17172 4023
rect 17494 4020 17500 4032
rect 17552 4020 17558 4072
rect 19705 4063 19763 4069
rect 19705 4029 19717 4063
rect 19751 4060 19763 4063
rect 20254 4060 20260 4072
rect 19751 4032 20260 4060
rect 19751 4029 19763 4032
rect 19705 4023 19763 4029
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 20993 4063 21051 4069
rect 20993 4060 21005 4063
rect 20588 4032 21005 4060
rect 20588 4020 20594 4032
rect 20993 4029 21005 4032
rect 21039 4029 21051 4063
rect 20993 4023 21051 4029
rect 18690 3992 18696 4004
rect 17144 3964 18696 3992
rect 16669 3955 16727 3961
rect 18690 3952 18696 3964
rect 18748 3952 18754 4004
rect 20438 3992 20444 4004
rect 20399 3964 20444 3992
rect 20438 3952 20444 3964
rect 20496 3952 20502 4004
rect 12710 3924 12716 3936
rect 11808 3896 12716 3924
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 15194 3924 15200 3936
rect 15155 3896 15200 3924
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 15657 3927 15715 3933
rect 15657 3893 15669 3927
rect 15703 3924 15715 3927
rect 16574 3924 16580 3936
rect 15703 3896 16580 3924
rect 15703 3893 15715 3896
rect 15657 3887 15715 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 17865 3927 17923 3933
rect 17865 3893 17877 3927
rect 17911 3924 17923 3927
rect 18230 3924 18236 3936
rect 17911 3896 18236 3924
rect 17911 3893 17923 3896
rect 17865 3887 17923 3893
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 18325 3927 18383 3933
rect 18325 3893 18337 3927
rect 18371 3924 18383 3927
rect 18414 3924 18420 3936
rect 18371 3896 18420 3924
rect 18371 3893 18383 3896
rect 18325 3887 18383 3893
rect 18414 3884 18420 3896
rect 18472 3884 18478 3936
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 19981 3927 20039 3933
rect 19981 3924 19993 3927
rect 18840 3896 19993 3924
rect 18840 3884 18846 3896
rect 19981 3893 19993 3896
rect 20027 3893 20039 3927
rect 19981 3887 20039 3893
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 2682 3720 2688 3732
rect 2643 3692 2688 3720
rect 2682 3680 2688 3692
rect 2740 3680 2746 3732
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 4154 3720 4160 3732
rect 3108 3692 4160 3720
rect 3108 3680 3114 3692
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4246 3680 4252 3732
rect 4304 3720 4310 3732
rect 4893 3723 4951 3729
rect 4893 3720 4905 3723
rect 4304 3692 4905 3720
rect 4304 3680 4310 3692
rect 4893 3689 4905 3692
rect 4939 3689 4951 3723
rect 4893 3683 4951 3689
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 6181 3723 6239 3729
rect 6181 3720 6193 3723
rect 5592 3692 6193 3720
rect 5592 3680 5598 3692
rect 6181 3689 6193 3692
rect 6227 3689 6239 3723
rect 6181 3683 6239 3689
rect 6288 3692 6684 3720
rect 2409 3655 2467 3661
rect 2409 3621 2421 3655
rect 2455 3652 2467 3655
rect 2866 3652 2872 3664
rect 2455 3624 2872 3652
rect 2455 3621 2467 3624
rect 2409 3615 2467 3621
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 4798 3612 4804 3664
rect 4856 3652 4862 3664
rect 6288 3652 6316 3692
rect 4856 3624 6316 3652
rect 6656 3652 6684 3692
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 6788 3692 7205 3720
rect 6788 3680 6794 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 7193 3683 7251 3689
rect 7650 3680 7656 3732
rect 7708 3720 7714 3732
rect 10410 3720 10416 3732
rect 7708 3692 10416 3720
rect 7708 3680 7714 3692
rect 10410 3680 10416 3692
rect 10468 3680 10474 3732
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 12805 3723 12863 3729
rect 10652 3692 12434 3720
rect 10652 3680 10658 3692
rect 8478 3652 8484 3664
rect 6656 3624 8484 3652
rect 4856 3612 4862 3624
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2130 3584 2136 3596
rect 1995 3556 2136 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 1872 3516 1900 3547
rect 2130 3544 2136 3556
rect 2188 3544 2194 3596
rect 3142 3584 3148 3596
rect 3103 3556 3148 3584
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 3329 3587 3387 3593
rect 3329 3553 3341 3587
rect 3375 3584 3387 3587
rect 4154 3584 4160 3596
rect 3375 3556 4160 3584
rect 3375 3553 3387 3556
rect 3329 3547 3387 3553
rect 3344 3516 3372 3547
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 4338 3584 4344 3596
rect 4299 3556 4344 3584
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 4982 3544 4988 3596
rect 5040 3584 5046 3596
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 5040 3556 5457 3584
rect 5040 3544 5046 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 5534 3544 5540 3596
rect 5592 3584 5598 3596
rect 6270 3584 6276 3596
rect 5592 3556 6276 3584
rect 5592 3544 5598 3556
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 6840 3593 6868 3624
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 9033 3655 9091 3661
rect 9033 3621 9045 3655
rect 9079 3652 9091 3655
rect 9398 3652 9404 3664
rect 9079 3624 9404 3652
rect 9079 3621 9091 3624
rect 9033 3615 9091 3621
rect 9398 3612 9404 3624
rect 9456 3612 9462 3664
rect 12066 3652 12072 3664
rect 12027 3624 12072 3652
rect 12066 3612 12072 3624
rect 12124 3612 12130 3664
rect 6825 3587 6883 3593
rect 6825 3553 6837 3587
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 7466 3544 7472 3596
rect 7524 3584 7530 3596
rect 7653 3587 7711 3593
rect 7653 3584 7665 3587
rect 7524 3556 7665 3584
rect 7524 3544 7530 3556
rect 7653 3553 7665 3556
rect 7699 3553 7711 3587
rect 7653 3547 7711 3553
rect 7837 3587 7895 3593
rect 7837 3553 7849 3587
rect 7883 3584 7895 3587
rect 10413 3587 10471 3593
rect 7883 3556 9444 3584
rect 7883 3553 7895 3556
rect 7837 3547 7895 3553
rect 1872 3488 3372 3516
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 5166 3516 5172 3528
rect 4295 3488 5172 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 5166 3476 5172 3488
rect 5224 3476 5230 3528
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 5350 3516 5356 3528
rect 5307 3488 5356 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 7561 3519 7619 3525
rect 6604 3488 6649 3516
rect 6604 3476 6610 3488
rect 7561 3485 7573 3519
rect 7607 3516 7619 3519
rect 8202 3516 8208 3528
rect 7607 3488 8208 3516
rect 7607 3485 7619 3488
rect 7561 3479 7619 3485
rect 7668 3460 7696 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8386 3516 8392 3528
rect 8347 3488 8392 3516
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 9416 3516 9444 3556
rect 10413 3553 10425 3587
rect 10459 3584 10471 3587
rect 10502 3584 10508 3596
rect 10459 3556 10508 3584
rect 10459 3553 10471 3556
rect 10413 3547 10471 3553
rect 10502 3544 10508 3556
rect 10560 3584 10566 3596
rect 10689 3587 10747 3593
rect 10689 3584 10701 3587
rect 10560 3556 10701 3584
rect 10560 3544 10566 3556
rect 10689 3553 10701 3556
rect 10735 3553 10747 3587
rect 12406 3584 12434 3692
rect 12805 3689 12817 3723
rect 12851 3720 12863 3723
rect 12894 3720 12900 3732
rect 12851 3692 12900 3720
rect 12851 3689 12863 3692
rect 12805 3683 12863 3689
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 15746 3720 15752 3732
rect 13228 3692 15752 3720
rect 13228 3680 13234 3692
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 16114 3720 16120 3732
rect 16075 3692 16120 3720
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16577 3723 16635 3729
rect 16577 3689 16589 3723
rect 16623 3720 16635 3723
rect 16942 3720 16948 3732
rect 16623 3692 16948 3720
rect 16623 3689 16635 3692
rect 16577 3683 16635 3689
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 17034 3680 17040 3732
rect 17092 3720 17098 3732
rect 17497 3723 17555 3729
rect 17497 3720 17509 3723
rect 17092 3692 17509 3720
rect 17092 3680 17098 3692
rect 17497 3689 17509 3692
rect 17543 3689 17555 3723
rect 17497 3683 17555 3689
rect 18230 3680 18236 3732
rect 18288 3720 18294 3732
rect 18288 3692 19012 3720
rect 18288 3680 18294 3692
rect 13541 3655 13599 3661
rect 13541 3621 13553 3655
rect 13587 3652 13599 3655
rect 14642 3652 14648 3664
rect 13587 3624 14648 3652
rect 13587 3621 13599 3624
rect 13541 3615 13599 3621
rect 14642 3612 14648 3624
rect 14700 3612 14706 3664
rect 17862 3612 17868 3664
rect 17920 3652 17926 3664
rect 17920 3624 18920 3652
rect 17920 3612 17926 3624
rect 14366 3584 14372 3596
rect 12406 3556 14372 3584
rect 10689 3547 10747 3553
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 14734 3584 14740 3596
rect 14695 3556 14740 3584
rect 14734 3544 14740 3556
rect 14792 3544 14798 3596
rect 18138 3584 18144 3596
rect 18099 3556 18144 3584
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 10134 3516 10140 3528
rect 10192 3525 10198 3528
rect 9416 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3516 10204 3525
rect 11974 3516 11980 3528
rect 10192 3488 10237 3516
rect 10336 3488 11980 3516
rect 10192 3479 10204 3488
rect 10192 3476 10198 3479
rect 2038 3448 2044 3460
rect 1999 3420 2044 3448
rect 2038 3408 2044 3420
rect 2096 3408 2102 3460
rect 3053 3451 3111 3457
rect 3053 3417 3065 3451
rect 3099 3448 3111 3451
rect 3099 3420 3832 3448
rect 3099 3417 3111 3420
rect 3053 3411 3111 3417
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3418 3380 3424 3392
rect 3016 3352 3424 3380
rect 3016 3340 3022 3352
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 3804 3389 3832 3420
rect 4614 3408 4620 3460
rect 4672 3448 4678 3460
rect 6641 3451 6699 3457
rect 6641 3448 6653 3451
rect 4672 3420 6653 3448
rect 4672 3408 4678 3420
rect 6641 3417 6653 3420
rect 6687 3417 6699 3451
rect 6641 3411 6699 3417
rect 7650 3408 7656 3460
rect 7708 3408 7714 3460
rect 10336 3448 10364 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 12250 3476 12256 3528
rect 12308 3516 12314 3528
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 12308 3488 12541 3516
rect 12308 3476 12314 3488
rect 12529 3485 12541 3488
rect 12575 3485 12587 3519
rect 12529 3479 12587 3485
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 14274 3516 14280 3528
rect 13403 3488 14136 3516
rect 14235 3488 14280 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 7760 3420 10364 3448
rect 3789 3383 3847 3389
rect 3789 3349 3801 3383
rect 3835 3349 3847 3383
rect 4154 3380 4160 3392
rect 4115 3352 4160 3380
rect 3789 3343 3847 3349
rect 4154 3340 4160 3352
rect 4212 3380 4218 3392
rect 4522 3380 4528 3392
rect 4212 3352 4528 3380
rect 4212 3340 4218 3352
rect 4522 3340 4528 3352
rect 4580 3340 4586 3392
rect 5350 3340 5356 3392
rect 5408 3380 5414 3392
rect 5408 3352 5453 3380
rect 5408 3340 5414 3352
rect 5626 3340 5632 3392
rect 5684 3380 5690 3392
rect 5994 3380 6000 3392
rect 5684 3352 6000 3380
rect 5684 3340 5690 3352
rect 5994 3340 6000 3352
rect 6052 3380 6058 3392
rect 7760 3380 7788 3420
rect 10686 3408 10692 3460
rect 10744 3448 10750 3460
rect 10934 3451 10992 3457
rect 10934 3448 10946 3451
rect 10744 3420 10946 3448
rect 10744 3408 10750 3420
rect 10934 3417 10946 3420
rect 10980 3417 10992 3451
rect 10934 3411 10992 3417
rect 11606 3408 11612 3460
rect 11664 3448 11670 3460
rect 11790 3448 11796 3460
rect 11664 3420 11796 3448
rect 11664 3408 11670 3420
rect 11790 3408 11796 3420
rect 11848 3448 11854 3460
rect 13004 3448 13032 3479
rect 11848 3420 13032 3448
rect 11848 3408 11854 3420
rect 8570 3380 8576 3392
rect 6052 3352 7788 3380
rect 8531 3352 8576 3380
rect 6052 3340 6058 3352
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 9030 3340 9036 3392
rect 9088 3380 9094 3392
rect 9490 3380 9496 3392
rect 9088 3352 9496 3380
rect 9088 3340 9094 3352
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 11698 3380 11704 3392
rect 9732 3352 11704 3380
rect 9732 3340 9738 3352
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 12342 3380 12348 3392
rect 12303 3352 12348 3380
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 14108 3389 14136 3488
rect 14274 3476 14280 3488
rect 14332 3476 14338 3528
rect 16390 3516 16396 3528
rect 16351 3488 16396 3516
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16632 3488 16865 3516
rect 16632 3476 16638 3488
rect 16853 3485 16865 3488
rect 16899 3485 16911 3519
rect 17310 3516 17316 3528
rect 16853 3479 16911 3485
rect 16960 3488 17316 3516
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 14982 3451 15040 3457
rect 14982 3448 14994 3451
rect 14884 3420 14994 3448
rect 14884 3408 14890 3420
rect 14982 3417 14994 3420
rect 15028 3448 15040 3451
rect 15102 3448 15108 3460
rect 15028 3420 15108 3448
rect 15028 3417 15040 3420
rect 14982 3411 15040 3417
rect 15102 3408 15108 3420
rect 15160 3408 15166 3460
rect 14093 3383 14151 3389
rect 14093 3349 14105 3383
rect 14139 3349 14151 3383
rect 14093 3343 14151 3349
rect 14182 3340 14188 3392
rect 14240 3380 14246 3392
rect 16960 3380 16988 3488
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17865 3519 17923 3525
rect 17865 3485 17877 3519
rect 17911 3516 17923 3519
rect 17954 3516 17960 3528
rect 17911 3488 17960 3516
rect 17911 3485 17923 3488
rect 17865 3479 17923 3485
rect 17954 3476 17960 3488
rect 18012 3476 18018 3528
rect 18782 3516 18788 3528
rect 18743 3488 18788 3516
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 18892 3516 18920 3624
rect 18984 3584 19012 3692
rect 19794 3680 19800 3732
rect 19852 3720 19858 3732
rect 20625 3723 20683 3729
rect 20625 3720 20637 3723
rect 19852 3692 20637 3720
rect 19852 3680 19858 3692
rect 20625 3689 20637 3692
rect 20671 3689 20683 3723
rect 20625 3683 20683 3689
rect 19058 3612 19064 3664
rect 19116 3652 19122 3664
rect 19981 3655 20039 3661
rect 19981 3652 19993 3655
rect 19116 3624 19993 3652
rect 19116 3612 19122 3624
rect 19981 3621 19993 3624
rect 20027 3621 20039 3655
rect 19981 3615 20039 3621
rect 20162 3584 20168 3596
rect 18984 3556 20168 3584
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 20898 3544 20904 3596
rect 20956 3584 20962 3596
rect 21177 3587 21235 3593
rect 21177 3584 21189 3587
rect 20956 3556 21189 3584
rect 20956 3544 20962 3556
rect 21177 3553 21189 3556
rect 21223 3553 21235 3587
rect 21177 3547 21235 3553
rect 19245 3519 19303 3525
rect 19245 3516 19257 3519
rect 18892 3488 19257 3516
rect 19245 3485 19257 3488
rect 19291 3485 19303 3519
rect 19245 3479 19303 3485
rect 19702 3476 19708 3528
rect 19760 3516 19766 3528
rect 19797 3519 19855 3525
rect 19797 3516 19809 3519
rect 19760 3488 19809 3516
rect 19760 3476 19766 3488
rect 19797 3485 19809 3488
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 21085 3519 21143 3525
rect 21085 3485 21097 3519
rect 21131 3516 21143 3519
rect 21542 3516 21548 3528
rect 21131 3488 21548 3516
rect 21131 3485 21143 3488
rect 21085 3479 21143 3485
rect 21542 3476 21548 3488
rect 21600 3476 21606 3528
rect 18322 3448 18328 3460
rect 17052 3420 18328 3448
rect 17052 3389 17080 3420
rect 18322 3408 18328 3420
rect 18380 3408 18386 3460
rect 18414 3408 18420 3460
rect 18472 3408 18478 3460
rect 19150 3408 19156 3460
rect 19208 3448 19214 3460
rect 20993 3451 21051 3457
rect 20993 3448 21005 3451
rect 19208 3420 21005 3448
rect 19208 3408 19214 3420
rect 20993 3417 21005 3420
rect 21039 3417 21051 3451
rect 20993 3411 21051 3417
rect 14240 3352 16988 3380
rect 17037 3383 17095 3389
rect 14240 3340 14246 3352
rect 17037 3349 17049 3383
rect 17083 3349 17095 3383
rect 17037 3343 17095 3349
rect 17862 3340 17868 3392
rect 17920 3380 17926 3392
rect 17957 3383 18015 3389
rect 17957 3380 17969 3383
rect 17920 3352 17969 3380
rect 17920 3340 17926 3352
rect 17957 3349 17969 3352
rect 18003 3349 18015 3383
rect 18432 3380 18460 3408
rect 18601 3383 18659 3389
rect 18601 3380 18613 3383
rect 18432 3352 18613 3380
rect 17957 3343 18015 3349
rect 18601 3349 18613 3352
rect 18647 3349 18659 3383
rect 18601 3343 18659 3349
rect 18782 3340 18788 3392
rect 18840 3380 18846 3392
rect 19429 3383 19487 3389
rect 19429 3380 19441 3383
rect 18840 3352 19441 3380
rect 18840 3340 18846 3352
rect 19429 3349 19441 3352
rect 19475 3349 19487 3383
rect 19429 3343 19487 3349
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 1854 3136 1860 3188
rect 1912 3176 1918 3188
rect 4154 3176 4160 3188
rect 1912 3148 4160 3176
rect 1912 3136 1918 3148
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 5997 3179 6055 3185
rect 5997 3176 6009 3179
rect 5868 3148 6009 3176
rect 5868 3136 5874 3148
rect 5997 3145 6009 3148
rect 6043 3145 6055 3179
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 5997 3139 6055 3145
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 7650 3176 7656 3188
rect 7611 3148 7656 3176
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 8849 3179 8907 3185
rect 8849 3176 8861 3179
rect 8496 3148 8861 3176
rect 1210 3068 1216 3120
rect 1268 3108 1274 3120
rect 3970 3108 3976 3120
rect 1268 3080 3976 3108
rect 1268 3068 1274 3080
rect 3970 3068 3976 3080
rect 4028 3068 4034 3120
rect 5074 3068 5080 3120
rect 5132 3108 5138 3120
rect 7466 3108 7472 3120
rect 5132 3080 7472 3108
rect 5132 3068 5138 3080
rect 7466 3068 7472 3080
rect 7524 3108 7530 3120
rect 7561 3111 7619 3117
rect 7561 3108 7573 3111
rect 7524 3080 7573 3108
rect 7524 3068 7530 3080
rect 7561 3077 7573 3080
rect 7607 3077 7619 3111
rect 7561 3071 7619 3077
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2406 3040 2412 3052
rect 2271 3012 2412 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2590 3000 2596 3052
rect 2648 3040 2654 3052
rect 2685 3043 2743 3049
rect 2685 3040 2697 3043
rect 2648 3012 2697 3040
rect 2648 3000 2654 3012
rect 2685 3009 2697 3012
rect 2731 3009 2743 3043
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 2685 3003 2743 3009
rect 2884 3012 3157 3040
rect 2884 2913 2912 3012
rect 3145 3009 3157 3012
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 3878 3040 3884 3052
rect 3651 3012 3884 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 4062 3040 4068 3052
rect 4023 3012 4068 3040
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 4488 3012 5365 3040
rect 4488 3000 4494 3012
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 6086 3040 6092 3052
rect 5859 3012 6092 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6362 3040 6368 3052
rect 6323 3012 6368 3040
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6638 3040 6644 3052
rect 6512 3012 6644 3040
rect 6512 3000 6518 3012
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 8496 3040 8524 3148
rect 8849 3145 8861 3148
rect 8895 3176 8907 3179
rect 11698 3176 11704 3188
rect 8895 3148 11704 3176
rect 8895 3145 8907 3148
rect 8849 3139 8907 3145
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 15841 3179 15899 3185
rect 12176 3148 14228 3176
rect 8570 3068 8576 3120
rect 8628 3108 8634 3120
rect 12176 3108 12204 3148
rect 8628 3080 12204 3108
rect 8628 3068 8634 3080
rect 13446 3068 13452 3120
rect 13504 3108 13510 3120
rect 13541 3111 13599 3117
rect 13541 3108 13553 3111
rect 13504 3080 13553 3108
rect 13504 3068 13510 3080
rect 13541 3077 13553 3080
rect 13587 3077 13599 3111
rect 13541 3071 13599 3077
rect 7024 3012 8524 3040
rect 8941 3043 8999 3049
rect 4522 2932 4528 2984
rect 4580 2972 4586 2984
rect 5077 2975 5135 2981
rect 5077 2972 5089 2975
rect 4580 2944 5089 2972
rect 4580 2932 4586 2944
rect 5077 2941 5089 2944
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 2869 2907 2927 2913
rect 2869 2873 2881 2907
rect 2915 2873 2927 2907
rect 2869 2867 2927 2873
rect 3789 2907 3847 2913
rect 3789 2873 3801 2907
rect 3835 2904 3847 2907
rect 5902 2904 5908 2916
rect 3835 2876 5908 2904
rect 3835 2873 3847 2876
rect 3789 2867 3847 2873
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 6549 2907 6607 2913
rect 6549 2873 6561 2907
rect 6595 2904 6607 2907
rect 7024 2904 7052 3012
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 9306 3040 9312 3052
rect 8987 3012 9312 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 9674 3040 9680 3052
rect 9600 3012 9680 3040
rect 7469 2975 7527 2981
rect 7469 2941 7481 2975
rect 7515 2972 7527 2975
rect 9030 2972 9036 2984
rect 7515 2944 8524 2972
rect 8991 2944 9036 2972
rect 7515 2941 7527 2944
rect 7469 2935 7527 2941
rect 6595 2876 7052 2904
rect 8496 2904 8524 2944
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 9600 2981 9628 3012
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 9858 3040 9864 3052
rect 9819 3012 9864 3040
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 10778 3000 10784 3052
rect 10836 3040 10842 3052
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10836 3012 10885 3040
rect 10836 3000 10842 3012
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 11054 3040 11060 3052
rect 11015 3012 11060 3040
rect 10873 3003 10931 3009
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11974 3040 11980 3052
rect 11440 3012 11836 3040
rect 11935 3012 11980 3040
rect 9585 2975 9643 2981
rect 9585 2941 9597 2975
rect 9631 2941 9643 2975
rect 9766 2972 9772 2984
rect 9727 2944 9772 2972
rect 9585 2935 9643 2941
rect 9766 2932 9772 2944
rect 9824 2932 9830 2984
rect 11440 2904 11468 3012
rect 8496 2876 11468 2904
rect 11808 2904 11836 3012
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 12069 3043 12127 3049
rect 12069 3009 12081 3043
rect 12115 3040 12127 3043
rect 12526 3040 12532 3052
rect 12115 3012 12532 3040
rect 12115 3009 12127 3012
rect 12069 3003 12127 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12710 3040 12716 3052
rect 12671 3012 12716 3040
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 14200 3049 14228 3148
rect 15841 3145 15853 3179
rect 15887 3176 15899 3179
rect 17865 3179 17923 3185
rect 17865 3176 17877 3179
rect 15887 3148 17877 3176
rect 15887 3145 15899 3148
rect 15841 3139 15899 3145
rect 17865 3145 17877 3148
rect 17911 3145 17923 3179
rect 17865 3139 17923 3145
rect 17954 3136 17960 3188
rect 18012 3176 18018 3188
rect 18233 3179 18291 3185
rect 18233 3176 18245 3179
rect 18012 3148 18245 3176
rect 18012 3136 18018 3148
rect 18233 3145 18245 3148
rect 18279 3145 18291 3179
rect 18233 3139 18291 3145
rect 18690 3136 18696 3188
rect 18748 3176 18754 3188
rect 18877 3179 18935 3185
rect 18877 3176 18889 3179
rect 18748 3148 18889 3176
rect 18748 3136 18754 3148
rect 18877 3145 18889 3148
rect 18923 3145 18935 3179
rect 18877 3139 18935 3145
rect 19242 3136 19248 3188
rect 19300 3176 19306 3188
rect 19337 3179 19395 3185
rect 19337 3176 19349 3179
rect 19300 3148 19349 3176
rect 19300 3136 19306 3148
rect 19337 3145 19349 3148
rect 19383 3145 19395 3179
rect 19337 3139 19395 3145
rect 14642 3068 14648 3120
rect 14700 3108 14706 3120
rect 14700 3080 16712 3108
rect 14700 3068 14706 3080
rect 14185 3043 14243 3049
rect 14185 3009 14197 3043
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14424 3012 14841 3040
rect 14424 3000 14430 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 15930 3040 15936 3052
rect 15891 3012 15936 3040
rect 14829 3003 14887 3009
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 16684 3049 16712 3080
rect 17586 3068 17592 3120
rect 17644 3108 17650 3120
rect 18966 3108 18972 3120
rect 17644 3080 18972 3108
rect 17644 3068 17650 3080
rect 18966 3068 18972 3080
rect 19024 3068 19030 3120
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 17221 3043 17279 3049
rect 17221 3040 17233 3043
rect 17184 3012 17233 3040
rect 17184 3000 17190 3012
rect 17221 3009 17233 3012
rect 17267 3009 17279 3043
rect 17221 3003 17279 3009
rect 18325 3043 18383 3049
rect 18325 3009 18337 3043
rect 18371 3040 18383 3043
rect 18874 3040 18880 3052
rect 18371 3012 18880 3040
rect 18371 3009 18383 3012
rect 18325 3003 18383 3009
rect 18874 3000 18880 3012
rect 18932 3040 18938 3052
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 18932 3012 19257 3040
rect 18932 3000 18938 3012
rect 19245 3009 19257 3012
rect 19291 3009 19303 3043
rect 19978 3040 19984 3052
rect 19939 3012 19984 3040
rect 19245 3003 19303 3009
rect 19978 3000 19984 3012
rect 20036 3040 20042 3052
rect 20622 3040 20628 3052
rect 20036 3012 20628 3040
rect 20036 3000 20042 3012
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 20990 3000 20996 3052
rect 21048 3040 21054 3052
rect 21361 3043 21419 3049
rect 21361 3040 21373 3043
rect 21048 3012 21373 3040
rect 21048 3000 21054 3012
rect 21361 3009 21373 3012
rect 21407 3009 21419 3043
rect 21361 3003 21419 3009
rect 12161 2975 12219 2981
rect 12161 2941 12173 2975
rect 12207 2972 12219 2975
rect 13078 2972 13084 2984
rect 12207 2944 13084 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 12176 2904 12204 2935
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 13354 2972 13360 2984
rect 13315 2944 13360 2972
rect 13354 2932 13360 2944
rect 13412 2932 13418 2984
rect 13449 2975 13507 2981
rect 13449 2941 13461 2975
rect 13495 2941 13507 2975
rect 13449 2935 13507 2941
rect 13464 2904 13492 2935
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 15657 2975 15715 2981
rect 15657 2972 15669 2975
rect 15620 2944 15669 2972
rect 15620 2932 15626 2944
rect 15657 2941 15669 2944
rect 15703 2941 15715 2975
rect 16574 2972 16580 2984
rect 15657 2935 15715 2941
rect 15764 2944 16580 2972
rect 15764 2904 15792 2944
rect 16574 2932 16580 2944
rect 16632 2932 16638 2984
rect 18230 2932 18236 2984
rect 18288 2972 18294 2984
rect 18417 2975 18475 2981
rect 18417 2972 18429 2975
rect 18288 2944 18429 2972
rect 18288 2932 18294 2944
rect 18417 2941 18429 2944
rect 18463 2941 18475 2975
rect 18417 2935 18475 2941
rect 19429 2975 19487 2981
rect 19429 2941 19441 2975
rect 19475 2941 19487 2975
rect 20254 2972 20260 2984
rect 20215 2944 20260 2972
rect 19429 2935 19487 2941
rect 16853 2907 16911 2913
rect 16853 2904 16865 2907
rect 11808 2876 12204 2904
rect 12406 2876 13492 2904
rect 13832 2876 15792 2904
rect 15856 2876 16865 2904
rect 6595 2873 6607 2876
rect 6549 2867 6607 2873
rect 1118 2796 1124 2848
rect 1176 2836 1182 2848
rect 2774 2836 2780 2848
rect 1176 2808 2780 2836
rect 1176 2796 1182 2808
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 3329 2839 3387 2845
rect 3329 2805 3341 2839
rect 3375 2836 3387 2839
rect 3418 2836 3424 2848
rect 3375 2808 3424 2836
rect 3375 2805 3387 2808
rect 3329 2799 3387 2805
rect 3418 2796 3424 2808
rect 3476 2796 3482 2848
rect 4249 2839 4307 2845
rect 4249 2805 4261 2839
rect 4295 2836 4307 2839
rect 4338 2836 4344 2848
rect 4295 2808 4344 2836
rect 4295 2805 4307 2808
rect 4249 2799 4307 2805
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 8018 2836 8024 2848
rect 7979 2808 8024 2836
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 8481 2839 8539 2845
rect 8481 2805 8493 2839
rect 8527 2836 8539 2839
rect 8570 2836 8576 2848
rect 8527 2808 8576 2836
rect 8527 2805 8539 2808
rect 8481 2799 8539 2805
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 10229 2839 10287 2845
rect 10229 2805 10241 2839
rect 10275 2836 10287 2839
rect 10318 2836 10324 2848
rect 10275 2808 10324 2836
rect 10275 2805 10287 2808
rect 10229 2799 10287 2805
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 11606 2836 11612 2848
rect 11567 2808 11612 2836
rect 11606 2796 11612 2808
rect 11664 2796 11670 2848
rect 11698 2796 11704 2848
rect 11756 2836 11762 2848
rect 12406 2836 12434 2876
rect 11756 2808 12434 2836
rect 12897 2839 12955 2845
rect 11756 2796 11762 2808
rect 12897 2805 12909 2839
rect 12943 2836 12955 2839
rect 13832 2836 13860 2876
rect 15856 2848 15884 2876
rect 16853 2873 16865 2876
rect 16899 2873 16911 2907
rect 16853 2867 16911 2873
rect 18138 2864 18144 2916
rect 18196 2904 18202 2916
rect 19444 2904 19472 2935
rect 20254 2932 20260 2944
rect 20312 2932 20318 2984
rect 18196 2876 19472 2904
rect 18196 2864 18202 2876
rect 12943 2808 13860 2836
rect 13909 2839 13967 2845
rect 12943 2805 12955 2808
rect 12897 2799 12955 2805
rect 13909 2805 13921 2839
rect 13955 2836 13967 2839
rect 14182 2836 14188 2848
rect 13955 2808 14188 2836
rect 13955 2805 13967 2808
rect 13909 2799 13967 2805
rect 14182 2796 14188 2808
rect 14240 2796 14246 2848
rect 14274 2796 14280 2848
rect 14332 2836 14338 2848
rect 14369 2839 14427 2845
rect 14369 2836 14381 2839
rect 14332 2808 14381 2836
rect 14332 2796 14338 2808
rect 14369 2805 14381 2808
rect 14415 2805 14427 2839
rect 14369 2799 14427 2805
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 15013 2839 15071 2845
rect 15013 2836 15025 2839
rect 14792 2808 15025 2836
rect 14792 2796 14798 2808
rect 15013 2805 15025 2808
rect 15059 2805 15071 2839
rect 15013 2799 15071 2805
rect 15838 2796 15844 2848
rect 15896 2796 15902 2848
rect 16298 2836 16304 2848
rect 16259 2808 16304 2836
rect 16298 2796 16304 2808
rect 16356 2796 16362 2848
rect 16942 2796 16948 2848
rect 17000 2836 17006 2848
rect 17405 2839 17463 2845
rect 17405 2836 17417 2839
rect 17000 2808 17417 2836
rect 17000 2796 17006 2808
rect 17405 2805 17417 2808
rect 17451 2805 17463 2839
rect 17405 2799 17463 2805
rect 20070 2796 20076 2848
rect 20128 2836 20134 2848
rect 21177 2839 21235 2845
rect 21177 2836 21189 2839
rect 20128 2808 21189 2836
rect 20128 2796 20134 2808
rect 21177 2805 21189 2808
rect 21223 2805 21235 2839
rect 21177 2799 21235 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 1854 2632 1860 2644
rect 1815 2604 1860 2632
rect 1854 2592 1860 2604
rect 1912 2592 1918 2644
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 4522 2632 4528 2644
rect 2915 2604 4528 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 5350 2592 5356 2644
rect 5408 2632 5414 2644
rect 6825 2635 6883 2641
rect 5408 2604 6776 2632
rect 5408 2592 5414 2604
rect 2409 2567 2467 2573
rect 2409 2533 2421 2567
rect 2455 2564 2467 2567
rect 2958 2564 2964 2576
rect 2455 2536 2964 2564
rect 2455 2533 2467 2536
rect 2409 2527 2467 2533
rect 2958 2524 2964 2536
rect 3016 2524 3022 2576
rect 3970 2524 3976 2576
rect 4028 2564 4034 2576
rect 6454 2564 6460 2576
rect 4028 2536 6460 2564
rect 4028 2524 4034 2536
rect 6454 2524 6460 2536
rect 6512 2524 6518 2576
rect 6748 2564 6776 2604
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 7282 2632 7288 2644
rect 6871 2604 7288 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 7282 2592 7288 2604
rect 7340 2632 7346 2644
rect 9858 2632 9864 2644
rect 7340 2604 9864 2632
rect 7340 2592 7346 2604
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 12250 2632 12256 2644
rect 12211 2604 12256 2632
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 12406 2604 13584 2632
rect 6748 2536 6960 2564
rect 3694 2496 3700 2508
rect 1688 2468 3700 2496
rect 1210 2388 1216 2440
rect 1268 2428 1274 2440
rect 1688 2437 1716 2468
rect 3694 2456 3700 2468
rect 3752 2456 3758 2508
rect 4154 2456 4160 2508
rect 4212 2496 4218 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4212 2468 4629 2496
rect 4212 2456 4218 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 5166 2456 5172 2508
rect 5224 2496 5230 2508
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 5224 2468 5457 2496
rect 5224 2456 5230 2468
rect 5445 2465 5457 2468
rect 5491 2465 5503 2499
rect 6730 2496 6736 2508
rect 5445 2459 5503 2465
rect 5644 2468 6736 2496
rect 1673 2431 1731 2437
rect 1673 2428 1685 2431
rect 1268 2400 1685 2428
rect 1268 2388 1274 2400
rect 1673 2397 1685 2400
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 2056 2400 2636 2428
rect 658 2320 664 2372
rect 716 2360 722 2372
rect 2056 2360 2084 2400
rect 2222 2360 2228 2372
rect 716 2332 2084 2360
rect 2183 2332 2228 2360
rect 716 2320 722 2332
rect 2222 2320 2228 2332
rect 2280 2320 2286 2372
rect 2608 2360 2636 2400
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 3234 2428 3240 2440
rect 2832 2400 2877 2428
rect 3195 2400 3240 2428
rect 2832 2388 2838 2400
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 5644 2428 5672 2468
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 4387 2400 5672 2428
rect 5721 2431 5779 2437
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 5721 2397 5733 2431
rect 5767 2397 5779 2431
rect 5721 2391 5779 2397
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 6822 2428 6828 2440
rect 6687 2400 6828 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 3252 2360 3280 2388
rect 2608 2332 3280 2360
rect 4798 2320 4804 2372
rect 4856 2360 4862 2372
rect 5736 2360 5764 2391
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 4856 2332 5764 2360
rect 6932 2360 6960 2536
rect 7006 2524 7012 2576
rect 7064 2564 7070 2576
rect 12406 2564 12434 2604
rect 7064 2536 12434 2564
rect 7064 2524 7070 2536
rect 7650 2496 7656 2508
rect 7611 2468 7656 2496
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 8018 2456 8024 2508
rect 8076 2496 8082 2508
rect 9493 2499 9551 2505
rect 8076 2468 9444 2496
rect 8076 2456 8082 2468
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7064 2400 7941 2428
rect 7064 2388 7070 2400
rect 7929 2397 7941 2400
rect 7975 2428 7987 2431
rect 8202 2428 8208 2440
rect 7975 2400 8208 2428
rect 7975 2397 7987 2400
rect 7929 2391 7987 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2428 9275 2431
rect 9306 2428 9312 2440
rect 9263 2400 9312 2428
rect 9263 2397 9275 2400
rect 9217 2391 9275 2397
rect 6932 2332 7972 2360
rect 4856 2320 4862 2332
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 3476 2264 3521 2292
rect 3476 2252 3482 2264
rect 3970 2252 3976 2304
rect 4028 2292 4034 2304
rect 7098 2292 7104 2304
rect 4028 2264 7104 2292
rect 4028 2252 4034 2264
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 7944 2292 7972 2332
rect 8386 2292 8392 2304
rect 7944 2264 8392 2292
rect 8386 2252 8392 2264
rect 8444 2252 8450 2304
rect 8588 2292 8616 2391
rect 9306 2388 9312 2400
rect 9364 2388 9370 2440
rect 9416 2360 9444 2468
rect 9493 2465 9505 2499
rect 9539 2496 9551 2499
rect 10134 2496 10140 2508
rect 9539 2468 10140 2496
rect 9539 2465 9551 2468
rect 9493 2459 9551 2465
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 10594 2496 10600 2508
rect 10555 2468 10600 2496
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 11701 2499 11759 2505
rect 11701 2465 11713 2499
rect 11747 2496 11759 2499
rect 12434 2496 12440 2508
rect 11747 2468 12440 2496
rect 11747 2465 11759 2468
rect 11701 2459 11759 2465
rect 12434 2456 12440 2468
rect 12492 2456 12498 2508
rect 13556 2496 13584 2604
rect 14918 2592 14924 2644
rect 14976 2632 14982 2644
rect 18874 2632 18880 2644
rect 14976 2604 18880 2632
rect 14976 2592 14982 2604
rect 18874 2592 18880 2604
rect 18932 2592 18938 2644
rect 20625 2635 20683 2641
rect 20625 2601 20637 2635
rect 20671 2632 20683 2635
rect 20806 2632 20812 2644
rect 20671 2604 20812 2632
rect 20671 2601 20683 2604
rect 20625 2595 20683 2601
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 13630 2524 13636 2576
rect 13688 2564 13694 2576
rect 14829 2567 14887 2573
rect 14829 2564 14841 2567
rect 13688 2536 14841 2564
rect 13688 2524 13694 2536
rect 14829 2533 14841 2536
rect 14875 2533 14887 2567
rect 14829 2527 14887 2533
rect 15102 2524 15108 2576
rect 15160 2564 15166 2576
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 15160 2536 15945 2564
rect 15160 2524 15166 2536
rect 15933 2533 15945 2536
rect 15979 2533 15991 2567
rect 15933 2527 15991 2533
rect 17126 2524 17132 2576
rect 17184 2564 17190 2576
rect 17957 2567 18015 2573
rect 17957 2564 17969 2567
rect 17184 2536 17969 2564
rect 17184 2524 17190 2536
rect 17957 2533 17969 2536
rect 18003 2533 18015 2567
rect 17957 2527 18015 2533
rect 18046 2524 18052 2576
rect 18104 2564 18110 2576
rect 19889 2567 19947 2573
rect 19889 2564 19901 2567
rect 18104 2536 19901 2564
rect 18104 2524 18110 2536
rect 19889 2533 19901 2536
rect 19935 2533 19947 2567
rect 19889 2527 19947 2533
rect 20898 2524 20904 2576
rect 20956 2564 20962 2576
rect 20956 2536 21220 2564
rect 20956 2524 20962 2536
rect 13556 2468 14688 2496
rect 10042 2388 10048 2440
rect 10100 2428 10106 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 10100 2400 10333 2428
rect 10100 2388 10106 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 11664 2400 11805 2428
rect 11664 2388 11670 2400
rect 11793 2397 11805 2400
rect 11839 2397 11851 2431
rect 12618 2428 12624 2440
rect 12579 2400 12624 2428
rect 11793 2391 11851 2397
rect 12618 2388 12624 2400
rect 12676 2388 12682 2440
rect 13170 2428 13176 2440
rect 13131 2400 13176 2428
rect 13170 2388 13176 2400
rect 13228 2388 13234 2440
rect 14660 2437 14688 2468
rect 18874 2456 18880 2508
rect 18932 2496 18938 2508
rect 21192 2505 21220 2536
rect 21177 2499 21235 2505
rect 18932 2468 21036 2496
rect 18932 2456 18938 2468
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 14645 2431 14703 2437
rect 14645 2397 14657 2431
rect 14691 2397 14703 2431
rect 15194 2428 15200 2440
rect 15155 2400 15200 2428
rect 14645 2391 14703 2397
rect 11885 2363 11943 2369
rect 11885 2360 11897 2363
rect 9416 2332 11897 2360
rect 11885 2329 11897 2332
rect 11931 2329 11943 2363
rect 11885 2323 11943 2329
rect 12250 2320 12256 2372
rect 12308 2360 12314 2372
rect 14108 2360 14136 2391
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 15746 2428 15752 2440
rect 15707 2400 15752 2428
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16574 2388 16580 2440
rect 16632 2428 16638 2440
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 16632 2400 16681 2428
rect 16632 2388 16638 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 17218 2428 17224 2440
rect 17179 2400 17224 2428
rect 16669 2391 16727 2397
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 17770 2428 17776 2440
rect 17731 2400 17776 2428
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 18322 2428 18328 2440
rect 18283 2400 18328 2428
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 18564 2400 19257 2428
rect 18564 2388 18570 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 20070 2428 20076 2440
rect 20031 2400 20076 2428
rect 19245 2391 19303 2397
rect 20070 2388 20076 2400
rect 20128 2388 20134 2440
rect 21008 2437 21036 2468
rect 21177 2465 21189 2499
rect 21223 2465 21235 2499
rect 21177 2459 21235 2465
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 12308 2332 14136 2360
rect 12308 2320 12314 2332
rect 14366 2320 14372 2372
rect 14424 2360 14430 2372
rect 14424 2332 15424 2360
rect 14424 2320 14430 2332
rect 11238 2292 11244 2304
rect 8588 2264 11244 2292
rect 11238 2252 11244 2264
rect 11296 2292 11302 2304
rect 11974 2292 11980 2304
rect 11296 2264 11980 2292
rect 11296 2252 11302 2264
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 12434 2292 12440 2304
rect 12124 2264 12440 2292
rect 12124 2252 12130 2264
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 12526 2252 12532 2304
rect 12584 2292 12590 2304
rect 12805 2295 12863 2301
rect 12805 2292 12817 2295
rect 12584 2264 12817 2292
rect 12584 2252 12590 2264
rect 12805 2261 12817 2264
rect 12851 2261 12863 2295
rect 12805 2255 12863 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13357 2295 13415 2301
rect 13357 2292 13369 2295
rect 12952 2264 13369 2292
rect 12952 2252 12958 2264
rect 13357 2261 13369 2264
rect 13403 2261 13415 2295
rect 13357 2255 13415 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 15396 2301 15424 2332
rect 16206 2320 16212 2372
rect 16264 2360 16270 2372
rect 16264 2332 17448 2360
rect 16264 2320 16270 2332
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13596 2264 14289 2292
rect 13596 2252 13602 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 15381 2295 15439 2301
rect 15381 2261 15393 2295
rect 15427 2261 15439 2295
rect 15381 2255 15439 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 17420 2301 17448 2332
rect 17678 2320 17684 2372
rect 17736 2360 17742 2372
rect 21085 2363 21143 2369
rect 17736 2332 19472 2360
rect 17736 2320 17742 2332
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 15528 2264 16865 2292
rect 15528 2252 15534 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 17405 2295 17463 2301
rect 17405 2261 17417 2295
rect 17451 2261 17463 2295
rect 17405 2255 17463 2261
rect 17586 2252 17592 2304
rect 17644 2292 17650 2304
rect 19444 2301 19472 2332
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 21174 2360 21180 2372
rect 21131 2332 21180 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 21174 2320 21180 2332
rect 21232 2320 21238 2372
rect 18509 2295 18567 2301
rect 18509 2292 18521 2295
rect 17644 2264 18521 2292
rect 17644 2252 17650 2264
rect 18509 2261 18521 2264
rect 18555 2261 18567 2295
rect 18509 2255 18567 2261
rect 19429 2295 19487 2301
rect 19429 2261 19441 2295
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 750 2048 756 2100
rect 808 2088 814 2100
rect 4798 2088 4804 2100
rect 808 2060 4804 2088
rect 808 2048 814 2060
rect 4798 2048 4804 2060
rect 4856 2048 4862 2100
rect 6822 2048 6828 2100
rect 6880 2088 6886 2100
rect 9950 2088 9956 2100
rect 6880 2060 9956 2088
rect 6880 2048 6886 2060
rect 9950 2048 9956 2060
rect 10008 2088 10014 2100
rect 10962 2088 10968 2100
rect 10008 2060 10968 2088
rect 10008 2048 10014 2060
rect 10962 2048 10968 2060
rect 11020 2048 11026 2100
rect 12434 2048 12440 2100
rect 12492 2088 12498 2100
rect 13446 2088 13452 2100
rect 12492 2060 13452 2088
rect 12492 2048 12498 2060
rect 13446 2048 13452 2060
rect 13504 2048 13510 2100
rect 13722 2048 13728 2100
rect 13780 2088 13786 2100
rect 19242 2088 19248 2100
rect 13780 2060 19248 2088
rect 13780 2048 13786 2060
rect 19242 2048 19248 2060
rect 19300 2048 19306 2100
rect 3234 1980 3240 2032
rect 3292 2020 3298 2032
rect 6270 2020 6276 2032
rect 3292 1992 6276 2020
rect 3292 1980 3298 1992
rect 6270 1980 6276 1992
rect 6328 1980 6334 2032
rect 7558 1980 7564 2032
rect 7616 2020 7622 2032
rect 13170 2020 13176 2032
rect 7616 1992 13176 2020
rect 7616 1980 7622 1992
rect 13170 1980 13176 1992
rect 13228 1980 13234 2032
rect 3418 1912 3424 1964
rect 3476 1952 3482 1964
rect 9490 1952 9496 1964
rect 3476 1924 9496 1952
rect 3476 1912 3482 1924
rect 9490 1912 9496 1924
rect 9548 1912 9554 1964
rect 8386 1844 8392 1896
rect 8444 1884 8450 1896
rect 12066 1884 12072 1896
rect 8444 1856 12072 1884
rect 8444 1844 8450 1856
rect 12066 1844 12072 1856
rect 12124 1844 12130 1896
rect 3510 1776 3516 1828
rect 3568 1816 3574 1828
rect 12250 1816 12256 1828
rect 3568 1788 12256 1816
rect 3568 1776 3574 1788
rect 12250 1776 12256 1788
rect 12308 1776 12314 1828
rect 4338 1708 4344 1760
rect 4396 1748 4402 1760
rect 12618 1748 12624 1760
rect 4396 1720 12624 1748
rect 4396 1708 4402 1720
rect 12618 1708 12624 1720
rect 12676 1708 12682 1760
<< via1 >>
rect 16120 20748 16172 20800
rect 17960 20748 18012 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 2044 20587 2096 20596
rect 2044 20553 2053 20587
rect 2053 20553 2087 20587
rect 2087 20553 2096 20587
rect 2044 20544 2096 20553
rect 5724 20544 5776 20596
rect 1676 20451 1728 20460
rect 1676 20417 1685 20451
rect 1685 20417 1719 20451
rect 1719 20417 1728 20451
rect 1676 20408 1728 20417
rect 2596 20408 2648 20460
rect 2964 20451 3016 20460
rect 2964 20417 2973 20451
rect 2973 20417 3007 20451
rect 3007 20417 3016 20451
rect 2964 20408 3016 20417
rect 5172 20340 5224 20392
rect 4712 20272 4764 20324
rect 12072 20476 12124 20528
rect 17224 20544 17276 20596
rect 21640 20544 21692 20596
rect 19892 20476 19944 20528
rect 7472 20408 7524 20460
rect 16120 20451 16172 20460
rect 7564 20340 7616 20392
rect 7012 20272 7064 20324
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 2228 20204 2280 20256
rect 3424 20204 3476 20256
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 4160 20247 4212 20256
rect 4160 20213 4169 20247
rect 4169 20213 4203 20247
rect 4203 20213 4212 20247
rect 4160 20204 4212 20213
rect 5264 20247 5316 20256
rect 5264 20213 5273 20247
rect 5273 20213 5307 20247
rect 5307 20213 5316 20247
rect 5264 20204 5316 20213
rect 7656 20204 7708 20256
rect 13452 20383 13504 20392
rect 8300 20247 8352 20256
rect 8300 20213 8309 20247
rect 8309 20213 8343 20247
rect 8343 20213 8352 20247
rect 8300 20204 8352 20213
rect 10324 20247 10376 20256
rect 10324 20213 10333 20247
rect 10333 20213 10367 20247
rect 10367 20213 10376 20247
rect 10324 20204 10376 20213
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 13452 20349 13461 20383
rect 13461 20349 13495 20383
rect 13495 20349 13504 20383
rect 13452 20340 13504 20349
rect 15384 20340 15436 20392
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 16304 20340 16356 20392
rect 13820 20272 13872 20324
rect 14648 20272 14700 20324
rect 12716 20204 12768 20256
rect 13544 20204 13596 20256
rect 14924 20204 14976 20256
rect 19708 20451 19760 20460
rect 19708 20417 19717 20451
rect 19717 20417 19751 20451
rect 19751 20417 19760 20451
rect 19708 20408 19760 20417
rect 19800 20408 19852 20460
rect 18236 20383 18288 20392
rect 18236 20349 18245 20383
rect 18245 20349 18279 20383
rect 18279 20349 18288 20383
rect 18236 20340 18288 20349
rect 18880 20383 18932 20392
rect 18880 20349 18889 20383
rect 18889 20349 18923 20383
rect 18923 20349 18932 20383
rect 18880 20340 18932 20349
rect 17224 20204 17276 20256
rect 19524 20247 19576 20256
rect 19524 20213 19533 20247
rect 19533 20213 19567 20247
rect 19567 20213 19576 20247
rect 19524 20204 19576 20213
rect 20168 20247 20220 20256
rect 20168 20213 20177 20247
rect 20177 20213 20211 20247
rect 20211 20213 20220 20247
rect 20168 20204 20220 20213
rect 20720 20247 20772 20256
rect 20720 20213 20729 20247
rect 20729 20213 20763 20247
rect 20763 20213 20772 20247
rect 20720 20204 20772 20213
rect 21272 20247 21324 20256
rect 21272 20213 21281 20247
rect 21281 20213 21315 20247
rect 21315 20213 21324 20247
rect 21272 20204 21324 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 1676 20000 1728 20052
rect 2596 20000 2648 20052
rect 10876 20000 10928 20052
rect 19708 20000 19760 20052
rect 20628 20000 20680 20052
rect 1952 19932 2004 19984
rect 4344 19864 4396 19916
rect 13360 19932 13412 19984
rect 19800 19932 19852 19984
rect 10784 19864 10836 19916
rect 11704 19864 11756 19916
rect 11888 19864 11940 19916
rect 13820 19864 13872 19916
rect 14648 19864 14700 19916
rect 15200 19907 15252 19916
rect 15200 19873 15209 19907
rect 15209 19873 15243 19907
rect 15243 19873 15252 19907
rect 15200 19864 15252 19873
rect 16304 19864 16356 19916
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 2688 19839 2740 19848
rect 2688 19805 2697 19839
rect 2697 19805 2731 19839
rect 2731 19805 2740 19839
rect 2688 19796 2740 19805
rect 3792 19796 3844 19848
rect 4436 19796 4488 19848
rect 6920 19796 6972 19848
rect 8300 19796 8352 19848
rect 8484 19796 8536 19848
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 12072 19796 12124 19805
rect 12624 19796 12676 19848
rect 13544 19796 13596 19848
rect 15384 19839 15436 19848
rect 7472 19728 7524 19780
rect 15384 19805 15393 19839
rect 15393 19805 15427 19839
rect 15427 19805 15436 19839
rect 15384 19796 15436 19805
rect 16212 19796 16264 19848
rect 20444 19864 20496 19916
rect 17500 19796 17552 19848
rect 18880 19796 18932 19848
rect 19800 19796 19852 19848
rect 20536 19839 20588 19848
rect 20536 19805 20545 19839
rect 20545 19805 20579 19839
rect 20579 19805 20588 19839
rect 20536 19796 20588 19805
rect 20812 19796 20864 19848
rect 17224 19728 17276 19780
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 4528 19703 4580 19712
rect 4528 19669 4537 19703
rect 4537 19669 4571 19703
rect 4571 19669 4580 19703
rect 4528 19660 4580 19669
rect 5356 19660 5408 19712
rect 6000 19660 6052 19712
rect 7012 19660 7064 19712
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7564 19660 7616 19669
rect 9312 19660 9364 19712
rect 11244 19703 11296 19712
rect 11244 19669 11253 19703
rect 11253 19669 11287 19703
rect 11287 19669 11296 19703
rect 11244 19660 11296 19669
rect 11980 19660 12032 19712
rect 13820 19660 13872 19712
rect 15752 19703 15804 19712
rect 15752 19669 15761 19703
rect 15761 19669 15795 19703
rect 15795 19669 15804 19703
rect 15752 19660 15804 19669
rect 15844 19660 15896 19712
rect 16396 19703 16448 19712
rect 16396 19669 16405 19703
rect 16405 19669 16439 19703
rect 16439 19669 16448 19703
rect 16396 19660 16448 19669
rect 17040 19703 17092 19712
rect 17040 19669 17049 19703
rect 17049 19669 17083 19703
rect 17083 19669 17092 19703
rect 17040 19660 17092 19669
rect 17592 19660 17644 19712
rect 18604 19660 18656 19712
rect 19984 19660 20036 19712
rect 21272 19703 21324 19712
rect 21272 19669 21281 19703
rect 21281 19669 21315 19703
rect 21315 19669 21324 19703
rect 21272 19660 21324 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 4620 19456 4672 19508
rect 5356 19499 5408 19508
rect 5356 19465 5365 19499
rect 5365 19465 5399 19499
rect 5399 19465 5408 19499
rect 5356 19456 5408 19465
rect 10048 19456 10100 19508
rect 10600 19499 10652 19508
rect 10600 19465 10609 19499
rect 10609 19465 10643 19499
rect 10643 19465 10652 19499
rect 10600 19456 10652 19465
rect 11244 19456 11296 19508
rect 13452 19499 13504 19508
rect 13452 19465 13461 19499
rect 13461 19465 13495 19499
rect 13495 19465 13504 19499
rect 13452 19456 13504 19465
rect 15844 19456 15896 19508
rect 16396 19456 16448 19508
rect 2688 19388 2740 19440
rect 3148 19388 3200 19440
rect 9956 19431 10008 19440
rect 9956 19397 9965 19431
rect 9965 19397 9999 19431
rect 9999 19397 10008 19431
rect 9956 19388 10008 19397
rect 16948 19431 17000 19440
rect 2228 19363 2280 19372
rect 2228 19329 2237 19363
rect 2237 19329 2271 19363
rect 2271 19329 2280 19363
rect 2228 19320 2280 19329
rect 2504 19363 2556 19372
rect 2504 19329 2513 19363
rect 2513 19329 2547 19363
rect 2547 19329 2556 19363
rect 2504 19320 2556 19329
rect 3424 19320 3476 19372
rect 4252 19320 4304 19372
rect 6736 19320 6788 19372
rect 11796 19363 11848 19372
rect 5632 19295 5684 19304
rect 2044 19227 2096 19236
rect 2044 19193 2053 19227
rect 2053 19193 2087 19227
rect 2087 19193 2096 19227
rect 2044 19184 2096 19193
rect 5632 19261 5641 19295
rect 5641 19261 5675 19295
rect 5675 19261 5684 19295
rect 5632 19252 5684 19261
rect 4344 19227 4396 19236
rect 4344 19193 4353 19227
rect 4353 19193 4387 19227
rect 4387 19193 4396 19227
rect 4344 19184 4396 19193
rect 7932 19252 7984 19304
rect 8392 19295 8444 19304
rect 8392 19261 8401 19295
rect 8401 19261 8435 19295
rect 8435 19261 8444 19295
rect 8392 19252 8444 19261
rect 10416 19295 10468 19304
rect 10416 19261 10425 19295
rect 10425 19261 10459 19295
rect 10459 19261 10468 19295
rect 10416 19252 10468 19261
rect 11796 19329 11805 19363
rect 11805 19329 11839 19363
rect 11839 19329 11848 19363
rect 11796 19320 11848 19329
rect 12532 19363 12584 19372
rect 11244 19252 11296 19304
rect 12532 19329 12541 19363
rect 12541 19329 12575 19363
rect 12575 19329 12584 19363
rect 12532 19320 12584 19329
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 3056 19116 3108 19168
rect 4988 19159 5040 19168
rect 4988 19125 4997 19159
rect 4997 19125 5031 19159
rect 5031 19125 5040 19159
rect 4988 19116 5040 19125
rect 6736 19159 6788 19168
rect 6736 19125 6745 19159
rect 6745 19125 6779 19159
rect 6779 19125 6788 19159
rect 6736 19116 6788 19125
rect 7564 19184 7616 19236
rect 11980 19252 12032 19304
rect 16948 19397 16957 19431
rect 16957 19397 16991 19431
rect 16991 19397 17000 19431
rect 16948 19388 17000 19397
rect 17500 19456 17552 19508
rect 18236 19499 18288 19508
rect 18236 19465 18245 19499
rect 18245 19465 18279 19499
rect 18279 19465 18288 19499
rect 18236 19456 18288 19465
rect 19064 19456 19116 19508
rect 19800 19456 19852 19508
rect 19984 19499 20036 19508
rect 19984 19465 19993 19499
rect 19993 19465 20027 19499
rect 20027 19465 20036 19499
rect 19984 19456 20036 19465
rect 20628 19456 20680 19508
rect 20812 19388 20864 19440
rect 14280 19320 14332 19372
rect 7748 19116 7800 19168
rect 7932 19116 7984 19168
rect 9220 19159 9272 19168
rect 9220 19125 9229 19159
rect 9229 19125 9263 19159
rect 9263 19125 9272 19159
rect 9220 19116 9272 19125
rect 10968 19159 11020 19168
rect 10968 19125 10977 19159
rect 10977 19125 11011 19159
rect 11011 19125 11020 19159
rect 10968 19116 11020 19125
rect 11888 19184 11940 19236
rect 12256 19227 12308 19236
rect 12256 19193 12265 19227
rect 12265 19193 12299 19227
rect 12299 19193 12308 19227
rect 12256 19184 12308 19193
rect 12440 19116 12492 19168
rect 12900 19252 12952 19304
rect 13544 19295 13596 19304
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 15200 19320 15252 19372
rect 15384 19320 15436 19372
rect 13452 19184 13504 19236
rect 15476 19252 15528 19304
rect 18880 19320 18932 19372
rect 20720 19320 20772 19372
rect 17132 19252 17184 19304
rect 18052 19184 18104 19236
rect 19616 19252 19668 19304
rect 21548 19184 21600 19236
rect 16304 19116 16356 19168
rect 17868 19159 17920 19168
rect 17868 19125 17877 19159
rect 17877 19125 17911 19159
rect 17911 19125 17920 19159
rect 17868 19116 17920 19125
rect 18512 19116 18564 19168
rect 19616 19116 19668 19168
rect 21364 19116 21416 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 2228 18912 2280 18964
rect 2504 18912 2556 18964
rect 5080 18912 5132 18964
rect 9956 18912 10008 18964
rect 10416 18912 10468 18964
rect 12532 18912 12584 18964
rect 12624 18912 12676 18964
rect 14740 18912 14792 18964
rect 15476 18955 15528 18964
rect 15476 18921 15485 18955
rect 15485 18921 15519 18955
rect 15519 18921 15528 18955
rect 15476 18912 15528 18921
rect 15568 18912 15620 18964
rect 18512 18912 18564 18964
rect 18880 18955 18932 18964
rect 18880 18921 18889 18955
rect 18889 18921 18923 18955
rect 18923 18921 18932 18955
rect 18880 18912 18932 18921
rect 19340 18912 19392 18964
rect 20536 18912 20588 18964
rect 1676 18844 1728 18896
rect 4712 18844 4764 18896
rect 9680 18887 9732 18896
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 3056 18751 3108 18760
rect 3056 18717 3065 18751
rect 3065 18717 3099 18751
rect 3099 18717 3108 18751
rect 3056 18708 3108 18717
rect 4988 18708 5040 18760
rect 2780 18640 2832 18692
rect 7840 18776 7892 18828
rect 8668 18776 8720 18828
rect 5632 18708 5684 18760
rect 6552 18708 6604 18760
rect 8392 18708 8444 18760
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 1676 18572 1728 18624
rect 3056 18572 3108 18624
rect 5540 18640 5592 18692
rect 7288 18640 7340 18692
rect 8300 18640 8352 18692
rect 9680 18853 9689 18887
rect 9689 18853 9723 18887
rect 9723 18853 9732 18887
rect 9680 18844 9732 18853
rect 14188 18844 14240 18896
rect 16948 18844 17000 18896
rect 10600 18819 10652 18828
rect 10600 18785 10609 18819
rect 10609 18785 10643 18819
rect 10643 18785 10652 18819
rect 10600 18776 10652 18785
rect 12808 18776 12860 18828
rect 14832 18776 14884 18828
rect 9496 18708 9548 18760
rect 13544 18708 13596 18760
rect 15108 18776 15160 18828
rect 19340 18776 19392 18828
rect 16396 18708 16448 18760
rect 17224 18708 17276 18760
rect 17592 18708 17644 18760
rect 18420 18751 18472 18760
rect 12808 18640 12860 18692
rect 16120 18640 16172 18692
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 4896 18572 4948 18624
rect 5816 18572 5868 18624
rect 6644 18615 6696 18624
rect 6644 18581 6653 18615
rect 6653 18581 6687 18615
rect 6687 18581 6696 18615
rect 6644 18572 6696 18581
rect 7012 18615 7064 18624
rect 7012 18581 7021 18615
rect 7021 18581 7055 18615
rect 7055 18581 7064 18615
rect 7012 18572 7064 18581
rect 7472 18615 7524 18624
rect 7472 18581 7481 18615
rect 7481 18581 7515 18615
rect 7515 18581 7524 18615
rect 7472 18572 7524 18581
rect 8024 18572 8076 18624
rect 8576 18615 8628 18624
rect 8576 18581 8585 18615
rect 8585 18581 8619 18615
rect 8619 18581 8628 18615
rect 8576 18572 8628 18581
rect 8944 18615 8996 18624
rect 8944 18581 8953 18615
rect 8953 18581 8987 18615
rect 8987 18581 8996 18615
rect 8944 18572 8996 18581
rect 11152 18572 11204 18624
rect 11980 18572 12032 18624
rect 12900 18572 12952 18624
rect 13636 18615 13688 18624
rect 13636 18581 13645 18615
rect 13645 18581 13679 18615
rect 13679 18581 13688 18615
rect 13636 18572 13688 18581
rect 14372 18615 14424 18624
rect 14372 18581 14381 18615
rect 14381 18581 14415 18615
rect 14415 18581 14424 18615
rect 14372 18572 14424 18581
rect 17960 18615 18012 18624
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 17960 18572 18012 18581
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 19524 18751 19576 18760
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 20628 18751 20680 18760
rect 20628 18717 20637 18751
rect 20637 18717 20671 18751
rect 20671 18717 20680 18751
rect 20628 18708 20680 18717
rect 19984 18615 20036 18624
rect 19984 18581 19993 18615
rect 19993 18581 20027 18615
rect 20027 18581 20036 18615
rect 19984 18572 20036 18581
rect 20076 18572 20128 18624
rect 21272 18615 21324 18624
rect 21272 18581 21281 18615
rect 21281 18581 21315 18615
rect 21315 18581 21324 18615
rect 21272 18572 21324 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 2136 18411 2188 18420
rect 2136 18377 2145 18411
rect 2145 18377 2179 18411
rect 2179 18377 2188 18411
rect 2136 18368 2188 18377
rect 2780 18368 2832 18420
rect 4528 18368 4580 18420
rect 8576 18368 8628 18420
rect 10140 18368 10192 18420
rect 11244 18368 11296 18420
rect 11980 18411 12032 18420
rect 11980 18377 11989 18411
rect 11989 18377 12023 18411
rect 12023 18377 12032 18411
rect 11980 18368 12032 18377
rect 12808 18411 12860 18420
rect 12808 18377 12817 18411
rect 12817 18377 12851 18411
rect 12851 18377 12860 18411
rect 12808 18368 12860 18377
rect 15752 18368 15804 18420
rect 4620 18343 4672 18352
rect 4620 18309 4629 18343
rect 4629 18309 4663 18343
rect 4663 18309 4672 18343
rect 4620 18300 4672 18309
rect 7012 18300 7064 18352
rect 8208 18300 8260 18352
rect 10048 18300 10100 18352
rect 15660 18300 15712 18352
rect 19524 18368 19576 18420
rect 20996 18368 21048 18420
rect 1952 18275 2004 18284
rect 1952 18241 1961 18275
rect 1961 18241 1995 18275
rect 1995 18241 2004 18275
rect 1952 18232 2004 18241
rect 2964 18232 3016 18284
rect 3056 18275 3108 18284
rect 3056 18241 3065 18275
rect 3065 18241 3099 18275
rect 3099 18241 3108 18275
rect 3056 18232 3108 18241
rect 7564 18232 7616 18284
rect 7748 18232 7800 18284
rect 8116 18207 8168 18216
rect 5632 18096 5684 18148
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8116 18164 8168 18173
rect 9128 18232 9180 18284
rect 14464 18275 14516 18284
rect 8576 18164 8628 18216
rect 8944 18164 8996 18216
rect 9864 18207 9916 18216
rect 9864 18173 9873 18207
rect 9873 18173 9907 18207
rect 9907 18173 9916 18207
rect 9864 18164 9916 18173
rect 13176 18207 13228 18216
rect 13176 18173 13185 18207
rect 13185 18173 13219 18207
rect 13219 18173 13228 18207
rect 13176 18164 13228 18173
rect 13360 18207 13412 18216
rect 13360 18173 13369 18207
rect 13369 18173 13403 18207
rect 13403 18173 13412 18207
rect 13360 18164 13412 18173
rect 14188 18207 14240 18216
rect 14188 18173 14197 18207
rect 14197 18173 14231 18207
rect 14231 18173 14240 18207
rect 14188 18164 14240 18173
rect 14464 18241 14473 18275
rect 14473 18241 14507 18275
rect 14507 18241 14516 18275
rect 14464 18232 14516 18241
rect 15108 18232 15160 18284
rect 16120 18275 16172 18284
rect 15568 18164 15620 18216
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 17408 18232 17460 18284
rect 18328 18232 18380 18284
rect 19064 18232 19116 18284
rect 20076 18232 20128 18284
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20812 18275 20864 18284
rect 20168 18232 20220 18241
rect 20812 18241 20821 18275
rect 20821 18241 20855 18275
rect 20855 18241 20864 18275
rect 20812 18232 20864 18241
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 3240 18028 3292 18080
rect 3976 18028 4028 18080
rect 5356 18071 5408 18080
rect 5356 18037 5365 18071
rect 5365 18037 5399 18071
rect 5399 18037 5408 18071
rect 5356 18028 5408 18037
rect 5724 18071 5776 18080
rect 5724 18037 5733 18071
rect 5733 18037 5767 18071
rect 5767 18037 5776 18071
rect 5724 18028 5776 18037
rect 5816 18028 5868 18080
rect 8576 18028 8628 18080
rect 9772 18096 9824 18148
rect 11796 18096 11848 18148
rect 17408 18096 17460 18148
rect 19524 18164 19576 18216
rect 18328 18096 18380 18148
rect 20720 18164 20772 18216
rect 21088 18096 21140 18148
rect 12072 18028 12124 18080
rect 18420 18028 18472 18080
rect 20260 18028 20312 18080
rect 21364 18028 21416 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 20 17824 72 17876
rect 1032 17824 1084 17876
rect 2780 17824 2832 17876
rect 6828 17867 6880 17876
rect 6828 17833 6837 17867
rect 6837 17833 6871 17867
rect 6871 17833 6880 17867
rect 6828 17824 6880 17833
rect 7380 17824 7432 17876
rect 8116 17824 8168 17876
rect 8392 17824 8444 17876
rect 11060 17824 11112 17876
rect 1860 17756 1912 17808
rect 4068 17756 4120 17808
rect 8760 17756 8812 17808
rect 17224 17824 17276 17876
rect 18236 17824 18288 17876
rect 18420 17867 18472 17876
rect 18420 17833 18429 17867
rect 18429 17833 18463 17867
rect 18463 17833 18472 17867
rect 18420 17824 18472 17833
rect 19524 17824 19576 17876
rect 12532 17756 12584 17808
rect 16120 17756 16172 17808
rect 16396 17756 16448 17808
rect 2228 17663 2280 17672
rect 2228 17629 2237 17663
rect 2237 17629 2271 17663
rect 2271 17629 2280 17663
rect 2228 17620 2280 17629
rect 3976 17688 4028 17740
rect 5356 17688 5408 17740
rect 5448 17688 5500 17740
rect 8392 17688 8444 17740
rect 10232 17688 10284 17740
rect 10416 17688 10468 17740
rect 11060 17731 11112 17740
rect 11060 17697 11069 17731
rect 11069 17697 11103 17731
rect 11103 17697 11112 17731
rect 11060 17688 11112 17697
rect 3240 17620 3292 17672
rect 6000 17620 6052 17672
rect 7380 17620 7432 17672
rect 12716 17731 12768 17740
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 2044 17527 2096 17536
rect 2044 17493 2053 17527
rect 2053 17493 2087 17527
rect 2087 17493 2096 17527
rect 2044 17484 2096 17493
rect 3976 17527 4028 17536
rect 3976 17493 3985 17527
rect 3985 17493 4019 17527
rect 4019 17493 4028 17527
rect 3976 17484 4028 17493
rect 4436 17527 4488 17536
rect 4436 17493 4445 17527
rect 4445 17493 4479 17527
rect 4479 17493 4488 17527
rect 4436 17484 4488 17493
rect 7932 17552 7984 17604
rect 10508 17552 10560 17604
rect 12256 17620 12308 17672
rect 12716 17697 12725 17731
rect 12725 17697 12759 17731
rect 12759 17697 12768 17731
rect 12716 17688 12768 17697
rect 15844 17688 15896 17740
rect 17960 17756 18012 17808
rect 12440 17620 12492 17672
rect 14556 17620 14608 17672
rect 11980 17552 12032 17604
rect 12348 17552 12400 17604
rect 17040 17552 17092 17604
rect 18144 17688 18196 17740
rect 17868 17620 17920 17672
rect 19616 17688 19668 17740
rect 19800 17688 19852 17740
rect 20444 17688 20496 17740
rect 18512 17620 18564 17672
rect 17592 17552 17644 17604
rect 18604 17552 18656 17604
rect 7012 17484 7064 17536
rect 7380 17484 7432 17536
rect 8208 17484 8260 17536
rect 9680 17527 9732 17536
rect 9680 17493 9689 17527
rect 9689 17493 9723 17527
rect 9723 17493 9732 17527
rect 9680 17484 9732 17493
rect 10140 17527 10192 17536
rect 10140 17493 10149 17527
rect 10149 17493 10183 17527
rect 10183 17493 10192 17527
rect 10140 17484 10192 17493
rect 12164 17527 12216 17536
rect 12164 17493 12173 17527
rect 12173 17493 12207 17527
rect 12207 17493 12216 17527
rect 12164 17484 12216 17493
rect 13544 17484 13596 17536
rect 14372 17527 14424 17536
rect 14372 17493 14381 17527
rect 14381 17493 14415 17527
rect 14415 17493 14424 17527
rect 14372 17484 14424 17493
rect 14648 17484 14700 17536
rect 14924 17484 14976 17536
rect 15200 17527 15252 17536
rect 15200 17493 15209 17527
rect 15209 17493 15243 17527
rect 15243 17493 15252 17527
rect 15200 17484 15252 17493
rect 15568 17484 15620 17536
rect 16396 17484 16448 17536
rect 17224 17527 17276 17536
rect 17224 17493 17233 17527
rect 17233 17493 17267 17527
rect 17267 17493 17276 17527
rect 17224 17484 17276 17493
rect 17684 17527 17736 17536
rect 17684 17493 17693 17527
rect 17693 17493 17727 17527
rect 17727 17493 17736 17527
rect 17684 17484 17736 17493
rect 19708 17595 19760 17604
rect 19708 17561 19717 17595
rect 19717 17561 19751 17595
rect 19751 17561 19760 17595
rect 19708 17552 19760 17561
rect 20352 17484 20404 17536
rect 20720 17527 20772 17536
rect 20720 17493 20729 17527
rect 20729 17493 20763 17527
rect 20763 17493 20772 17527
rect 20720 17484 20772 17493
rect 21456 17484 21508 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1952 17280 2004 17332
rect 2504 17144 2556 17196
rect 2688 17187 2740 17196
rect 2688 17153 2697 17187
rect 2697 17153 2731 17187
rect 2731 17153 2740 17187
rect 2688 17144 2740 17153
rect 5448 17280 5500 17332
rect 5632 17323 5684 17332
rect 5632 17289 5641 17323
rect 5641 17289 5675 17323
rect 5675 17289 5684 17323
rect 5632 17280 5684 17289
rect 5816 17280 5868 17332
rect 6828 17280 6880 17332
rect 7564 17323 7616 17332
rect 7564 17289 7573 17323
rect 7573 17289 7607 17323
rect 7607 17289 7616 17323
rect 7564 17280 7616 17289
rect 7932 17323 7984 17332
rect 7932 17289 7941 17323
rect 7941 17289 7975 17323
rect 7975 17289 7984 17323
rect 7932 17280 7984 17289
rect 9680 17280 9732 17332
rect 10324 17323 10376 17332
rect 10324 17289 10333 17323
rect 10333 17289 10367 17323
rect 10367 17289 10376 17323
rect 10324 17280 10376 17289
rect 12164 17280 12216 17332
rect 13268 17280 13320 17332
rect 13820 17323 13872 17332
rect 13820 17289 13829 17323
rect 13829 17289 13863 17323
rect 13863 17289 13872 17323
rect 13820 17280 13872 17289
rect 14464 17323 14516 17332
rect 14464 17289 14473 17323
rect 14473 17289 14507 17323
rect 14507 17289 14516 17323
rect 14464 17280 14516 17289
rect 15568 17323 15620 17332
rect 15568 17289 15577 17323
rect 15577 17289 15611 17323
rect 15611 17289 15620 17323
rect 15568 17280 15620 17289
rect 17684 17323 17736 17332
rect 17684 17289 17693 17323
rect 17693 17289 17727 17323
rect 17727 17289 17736 17323
rect 17684 17280 17736 17289
rect 17776 17280 17828 17332
rect 19064 17280 19116 17332
rect 20628 17280 20680 17332
rect 4068 17212 4120 17264
rect 13636 17212 13688 17264
rect 14280 17212 14332 17264
rect 14556 17212 14608 17264
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 3240 16940 3292 16992
rect 3884 17144 3936 17196
rect 4160 17076 4212 17128
rect 4988 17119 5040 17128
rect 4988 17085 4997 17119
rect 4997 17085 5031 17119
rect 5031 17085 5040 17119
rect 4988 17076 5040 17085
rect 6000 17076 6052 17128
rect 7012 17144 7064 17196
rect 7472 17144 7524 17196
rect 9496 17144 9548 17196
rect 14464 17144 14516 17196
rect 14832 17187 14884 17196
rect 14832 17153 14841 17187
rect 14841 17153 14875 17187
rect 14875 17153 14884 17187
rect 14832 17144 14884 17153
rect 7196 17076 7248 17128
rect 8024 17119 8076 17128
rect 8024 17085 8033 17119
rect 8033 17085 8067 17119
rect 8067 17085 8076 17119
rect 8024 17076 8076 17085
rect 8576 17076 8628 17128
rect 8668 17076 8720 17128
rect 10140 17119 10192 17128
rect 9864 17008 9916 17060
rect 10140 17085 10149 17119
rect 10149 17085 10183 17119
rect 10183 17085 10192 17119
rect 10140 17076 10192 17085
rect 11520 17119 11572 17128
rect 11520 17085 11529 17119
rect 11529 17085 11563 17119
rect 11563 17085 11572 17119
rect 11520 17076 11572 17085
rect 12532 17008 12584 17060
rect 14372 17076 14424 17128
rect 15200 17212 15252 17264
rect 15936 17187 15988 17196
rect 15936 17153 15945 17187
rect 15945 17153 15979 17187
rect 15979 17153 15988 17187
rect 15936 17144 15988 17153
rect 17684 17144 17736 17196
rect 18144 17144 18196 17196
rect 18420 17144 18472 17196
rect 18880 17187 18932 17196
rect 18880 17153 18889 17187
rect 18889 17153 18923 17187
rect 18923 17153 18932 17187
rect 18880 17144 18932 17153
rect 19800 17144 19852 17196
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 16212 17119 16264 17128
rect 13820 17008 13872 17060
rect 15568 17008 15620 17060
rect 16212 17085 16221 17119
rect 16221 17085 16255 17119
rect 16255 17085 16264 17119
rect 16212 17076 16264 17085
rect 18696 17119 18748 17128
rect 17408 17008 17460 17060
rect 4528 16940 4580 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5448 16940 5500 16992
rect 8760 16940 8812 16992
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 15752 16940 15804 16992
rect 18696 17085 18705 17119
rect 18705 17085 18739 17119
rect 18739 17085 18748 17119
rect 18696 17076 18748 17085
rect 19616 17076 19668 17128
rect 19708 17076 19760 17128
rect 17960 16940 18012 16992
rect 18512 16940 18564 16992
rect 18604 16940 18656 16992
rect 20720 16983 20772 16992
rect 20720 16949 20729 16983
rect 20729 16949 20763 16983
rect 20763 16949 20772 16983
rect 20720 16940 20772 16949
rect 21272 16983 21324 16992
rect 21272 16949 21281 16983
rect 21281 16949 21315 16983
rect 21315 16949 21324 16983
rect 21272 16940 21324 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1584 16668 1636 16720
rect 5080 16736 5132 16788
rect 7196 16736 7248 16788
rect 10048 16736 10100 16788
rect 4160 16643 4212 16652
rect 4160 16609 4169 16643
rect 4169 16609 4203 16643
rect 4203 16609 4212 16643
rect 6828 16668 6880 16720
rect 7104 16668 7156 16720
rect 7932 16668 7984 16720
rect 9956 16711 10008 16720
rect 9956 16677 9965 16711
rect 9965 16677 9999 16711
rect 9999 16677 10008 16711
rect 9956 16668 10008 16677
rect 11152 16736 11204 16788
rect 12164 16736 12216 16788
rect 12348 16736 12400 16788
rect 15292 16736 15344 16788
rect 16028 16736 16080 16788
rect 17316 16736 17368 16788
rect 17776 16736 17828 16788
rect 18880 16736 18932 16788
rect 19616 16779 19668 16788
rect 19616 16745 19625 16779
rect 19625 16745 19659 16779
rect 19659 16745 19668 16779
rect 19616 16736 19668 16745
rect 10692 16668 10744 16720
rect 4160 16600 4212 16609
rect 9220 16600 9272 16652
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 10324 16643 10376 16652
rect 10324 16609 10333 16643
rect 10333 16609 10367 16643
rect 10367 16609 10376 16643
rect 10324 16600 10376 16609
rect 10600 16600 10652 16652
rect 11060 16643 11112 16652
rect 11060 16609 11069 16643
rect 11069 16609 11103 16643
rect 11103 16609 11112 16643
rect 11060 16600 11112 16609
rect 13544 16668 13596 16720
rect 17500 16668 17552 16720
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 13636 16643 13688 16652
rect 13636 16609 13645 16643
rect 13645 16609 13679 16643
rect 13679 16609 13688 16643
rect 13636 16600 13688 16609
rect 14832 16600 14884 16652
rect 15476 16600 15528 16652
rect 1676 16575 1728 16584
rect 1676 16541 1685 16575
rect 1685 16541 1719 16575
rect 1719 16541 1728 16575
rect 1676 16532 1728 16541
rect 112 16464 164 16516
rect 1400 16464 1452 16516
rect 3240 16532 3292 16584
rect 3332 16532 3384 16584
rect 4988 16532 5040 16584
rect 7932 16532 7984 16584
rect 9312 16575 9364 16584
rect 9312 16541 9321 16575
rect 9321 16541 9355 16575
rect 9355 16541 9364 16575
rect 9312 16532 9364 16541
rect 13176 16532 13228 16584
rect 13728 16532 13780 16584
rect 5264 16464 5316 16516
rect 7748 16464 7800 16516
rect 12624 16464 12676 16516
rect 14924 16464 14976 16516
rect 17224 16600 17276 16652
rect 17776 16643 17828 16652
rect 17776 16609 17785 16643
rect 17785 16609 17819 16643
rect 17819 16609 17828 16643
rect 17776 16600 17828 16609
rect 18788 16600 18840 16652
rect 20904 16600 20956 16652
rect 21180 16643 21232 16652
rect 18512 16575 18564 16584
rect 18512 16541 18521 16575
rect 18521 16541 18555 16575
rect 18555 16541 18564 16575
rect 18512 16532 18564 16541
rect 17776 16464 17828 16516
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 2136 16439 2188 16448
rect 2136 16405 2145 16439
rect 2145 16405 2179 16439
rect 2179 16405 2188 16439
rect 2136 16396 2188 16405
rect 2596 16396 2648 16448
rect 2964 16396 3016 16448
rect 5080 16439 5132 16448
rect 5080 16405 5089 16439
rect 5089 16405 5123 16439
rect 5123 16405 5132 16439
rect 5080 16396 5132 16405
rect 5540 16439 5592 16448
rect 5540 16405 5549 16439
rect 5549 16405 5583 16439
rect 5583 16405 5592 16439
rect 5540 16396 5592 16405
rect 7196 16439 7248 16448
rect 7196 16405 7205 16439
rect 7205 16405 7239 16439
rect 7239 16405 7248 16439
rect 7196 16396 7248 16405
rect 8208 16439 8260 16448
rect 8208 16405 8217 16439
rect 8217 16405 8251 16439
rect 8251 16405 8260 16439
rect 8208 16396 8260 16405
rect 8392 16396 8444 16448
rect 9404 16439 9456 16448
rect 9404 16405 9413 16439
rect 9413 16405 9447 16439
rect 9447 16405 9456 16439
rect 9404 16396 9456 16405
rect 14648 16396 14700 16448
rect 15660 16439 15712 16448
rect 15660 16405 15669 16439
rect 15669 16405 15703 16439
rect 15703 16405 15712 16439
rect 15660 16396 15712 16405
rect 18512 16396 18564 16448
rect 20812 16532 20864 16584
rect 21180 16609 21189 16643
rect 21189 16609 21223 16643
rect 21223 16609 21232 16643
rect 21180 16600 21232 16609
rect 19064 16396 19116 16448
rect 19616 16396 19668 16448
rect 20168 16396 20220 16448
rect 20628 16439 20680 16448
rect 20628 16405 20637 16439
rect 20637 16405 20671 16439
rect 20671 16405 20680 16439
rect 20628 16396 20680 16405
rect 21088 16396 21140 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 2504 16235 2556 16244
rect 2504 16201 2513 16235
rect 2513 16201 2547 16235
rect 2547 16201 2556 16235
rect 2504 16192 2556 16201
rect 3332 16235 3384 16244
rect 3332 16201 3341 16235
rect 3341 16201 3375 16235
rect 3375 16201 3384 16235
rect 3332 16192 3384 16201
rect 2596 16056 2648 16108
rect 3884 16124 3936 16176
rect 5356 16192 5408 16244
rect 9404 16192 9456 16244
rect 10876 16192 10928 16244
rect 12624 16235 12676 16244
rect 7012 16124 7064 16176
rect 8116 16124 8168 16176
rect 4068 16056 4120 16108
rect 11428 16124 11480 16176
rect 12624 16201 12633 16235
rect 12633 16201 12667 16235
rect 12667 16201 12676 16235
rect 12624 16192 12676 16201
rect 15476 16235 15528 16244
rect 15476 16201 15485 16235
rect 15485 16201 15519 16235
rect 15519 16201 15528 16235
rect 15476 16192 15528 16201
rect 15936 16192 15988 16244
rect 18052 16192 18104 16244
rect 13176 16124 13228 16176
rect 15292 16124 15344 16176
rect 17500 16167 17552 16176
rect 17500 16133 17509 16167
rect 17509 16133 17543 16167
rect 17543 16133 17552 16167
rect 17500 16124 17552 16133
rect 2504 15988 2556 16040
rect 3700 15988 3752 16040
rect 6736 15988 6788 16040
rect 7104 16031 7156 16040
rect 7104 15997 7113 16031
rect 7113 15997 7147 16031
rect 7147 15997 7156 16031
rect 7104 15988 7156 15997
rect 8208 15988 8260 16040
rect 2044 15963 2096 15972
rect 2044 15929 2053 15963
rect 2053 15929 2087 15963
rect 2087 15929 2096 15963
rect 2044 15920 2096 15929
rect 2780 15920 2832 15972
rect 7564 15920 7616 15972
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 2872 15852 2924 15904
rect 4804 15852 4856 15904
rect 5172 15852 5224 15904
rect 7932 15852 7984 15904
rect 8208 15852 8260 15904
rect 10048 16056 10100 16108
rect 10876 16056 10928 16108
rect 14924 16099 14976 16108
rect 14924 16065 14933 16099
rect 14933 16065 14967 16099
rect 14967 16065 14976 16099
rect 14924 16056 14976 16065
rect 15568 16056 15620 16108
rect 14556 15988 14608 16040
rect 10324 15920 10376 15972
rect 10968 15920 11020 15972
rect 16948 15920 17000 15972
rect 18144 15963 18196 15972
rect 18144 15929 18153 15963
rect 18153 15929 18187 15963
rect 18187 15929 18196 15963
rect 18880 16056 18932 16108
rect 20628 16192 20680 16244
rect 19524 15988 19576 16040
rect 18144 15920 18196 15929
rect 18512 15920 18564 15972
rect 9404 15895 9456 15904
rect 9404 15861 9413 15895
rect 9413 15861 9447 15895
rect 9447 15861 9456 15895
rect 9404 15852 9456 15861
rect 10048 15895 10100 15904
rect 10048 15861 10057 15895
rect 10057 15861 10091 15895
rect 10091 15861 10100 15895
rect 10048 15852 10100 15861
rect 10876 15895 10928 15904
rect 10876 15861 10885 15895
rect 10885 15861 10919 15895
rect 10919 15861 10928 15895
rect 10876 15852 10928 15861
rect 12348 15895 12400 15904
rect 12348 15861 12357 15895
rect 12357 15861 12391 15895
rect 12391 15861 12400 15895
rect 12348 15852 12400 15861
rect 13360 15895 13412 15904
rect 13360 15861 13369 15895
rect 13369 15861 13403 15895
rect 13403 15861 13412 15895
rect 13360 15852 13412 15861
rect 14648 15895 14700 15904
rect 14648 15861 14657 15895
rect 14657 15861 14691 15895
rect 14691 15861 14700 15895
rect 14648 15852 14700 15861
rect 19892 15895 19944 15904
rect 19892 15861 19901 15895
rect 19901 15861 19935 15895
rect 19935 15861 19944 15895
rect 19892 15852 19944 15861
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 2504 15648 2556 15700
rect 5908 15648 5960 15700
rect 8668 15648 8720 15700
rect 1400 15580 1452 15632
rect 8208 15580 8260 15632
rect 8300 15580 8352 15632
rect 11152 15648 11204 15700
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 11704 15691 11756 15700
rect 11704 15657 11713 15691
rect 11713 15657 11747 15691
rect 11747 15657 11756 15691
rect 11704 15648 11756 15657
rect 17500 15648 17552 15700
rect 17684 15691 17736 15700
rect 17684 15657 17693 15691
rect 17693 15657 17727 15691
rect 17727 15657 17736 15691
rect 17684 15648 17736 15657
rect 4804 15512 4856 15564
rect 5080 15512 5132 15564
rect 5356 15512 5408 15564
rect 6368 15512 6420 15564
rect 7012 15512 7064 15564
rect 7564 15555 7616 15564
rect 7564 15521 7573 15555
rect 7573 15521 7607 15555
rect 7607 15521 7616 15555
rect 7564 15512 7616 15521
rect 8116 15512 8168 15564
rect 848 15444 900 15496
rect 1492 15444 1544 15496
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 2780 15444 2832 15496
rect 3976 15444 4028 15496
rect 6552 15444 6604 15496
rect 8760 15512 8812 15564
rect 8300 15444 8352 15496
rect 8484 15444 8536 15496
rect 9680 15444 9732 15496
rect 11244 15444 11296 15496
rect 3332 15376 3384 15428
rect 7564 15376 7616 15428
rect 10416 15419 10468 15428
rect 10416 15385 10434 15419
rect 10434 15385 10468 15419
rect 17408 15580 17460 15632
rect 17868 15580 17920 15632
rect 11428 15512 11480 15564
rect 11704 15444 11756 15496
rect 12164 15444 12216 15496
rect 15476 15512 15528 15564
rect 17040 15512 17092 15564
rect 19616 15512 19668 15564
rect 20076 15512 20128 15564
rect 13452 15444 13504 15496
rect 10416 15376 10468 15385
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 3240 15351 3292 15360
rect 3240 15317 3249 15351
rect 3249 15317 3283 15351
rect 3283 15317 3292 15351
rect 3240 15308 3292 15317
rect 4160 15308 4212 15360
rect 4528 15351 4580 15360
rect 4528 15317 4537 15351
rect 4537 15317 4571 15351
rect 4571 15317 4580 15351
rect 4528 15308 4580 15317
rect 4988 15351 5040 15360
rect 4988 15317 4997 15351
rect 4997 15317 5031 15351
rect 5031 15317 5040 15351
rect 4988 15308 5040 15317
rect 5356 15351 5408 15360
rect 5356 15317 5365 15351
rect 5365 15317 5399 15351
rect 5399 15317 5408 15351
rect 5356 15308 5408 15317
rect 7932 15308 7984 15360
rect 12348 15376 12400 15428
rect 14280 15376 14332 15428
rect 11980 15308 12032 15360
rect 12440 15351 12492 15360
rect 12440 15317 12449 15351
rect 12449 15317 12483 15351
rect 12483 15317 12492 15351
rect 12440 15308 12492 15317
rect 12624 15308 12676 15360
rect 12900 15308 12952 15360
rect 15108 15308 15160 15360
rect 15384 15308 15436 15360
rect 17500 15444 17552 15496
rect 18972 15444 19024 15496
rect 19984 15487 20036 15496
rect 19984 15453 19993 15487
rect 19993 15453 20027 15487
rect 20027 15453 20036 15487
rect 19984 15444 20036 15453
rect 20536 15487 20588 15496
rect 20536 15453 20545 15487
rect 20545 15453 20579 15487
rect 20579 15453 20588 15487
rect 20536 15444 20588 15453
rect 20996 15444 21048 15496
rect 17408 15308 17460 15360
rect 18052 15351 18104 15360
rect 18052 15317 18061 15351
rect 18061 15317 18095 15351
rect 18095 15317 18104 15351
rect 18052 15308 18104 15317
rect 19616 15351 19668 15360
rect 19616 15317 19625 15351
rect 19625 15317 19659 15351
rect 19659 15317 19668 15351
rect 19616 15308 19668 15317
rect 20168 15351 20220 15360
rect 20168 15317 20177 15351
rect 20177 15317 20211 15351
rect 20211 15317 20220 15351
rect 20168 15308 20220 15317
rect 20720 15351 20772 15360
rect 20720 15317 20729 15351
rect 20729 15317 20763 15351
rect 20763 15317 20772 15351
rect 20720 15308 20772 15317
rect 21364 15308 21416 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 3332 15104 3384 15156
rect 3424 15104 3476 15156
rect 4988 15104 5040 15156
rect 2412 15036 2464 15088
rect 5448 15036 5500 15088
rect 6000 15036 6052 15088
rect 11152 15104 11204 15156
rect 11244 15104 11296 15156
rect 12348 15104 12400 15156
rect 13452 15104 13504 15156
rect 15108 15104 15160 15156
rect 17224 15104 17276 15156
rect 20628 15104 20680 15156
rect 7104 15036 7156 15088
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 6920 14968 6972 15020
rect 7932 14968 7984 15020
rect 9588 14968 9640 15020
rect 4712 14943 4764 14952
rect 4712 14909 4721 14943
rect 4721 14909 4755 14943
rect 4755 14909 4764 14943
rect 4712 14900 4764 14909
rect 4804 14900 4856 14952
rect 5448 14900 5500 14952
rect 2964 14832 3016 14884
rect 3516 14875 3568 14884
rect 3516 14841 3525 14875
rect 3525 14841 3559 14875
rect 3559 14841 3568 14875
rect 3516 14832 3568 14841
rect 4068 14832 4120 14884
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 3148 14807 3200 14816
rect 3148 14773 3157 14807
rect 3157 14773 3191 14807
rect 3191 14773 3200 14807
rect 3148 14764 3200 14773
rect 4252 14807 4304 14816
rect 4252 14773 4261 14807
rect 4261 14773 4295 14807
rect 4295 14773 4304 14807
rect 4252 14764 4304 14773
rect 6000 14900 6052 14952
rect 7012 14900 7064 14952
rect 7472 14943 7524 14952
rect 7472 14909 7481 14943
rect 7481 14909 7515 14943
rect 7515 14909 7524 14943
rect 7472 14900 7524 14909
rect 7564 14943 7616 14952
rect 7564 14909 7573 14943
rect 7573 14909 7607 14943
rect 7607 14909 7616 14943
rect 10784 15036 10836 15088
rect 14004 15011 14056 15020
rect 14004 14977 14022 15011
rect 14022 14977 14056 15011
rect 14280 15011 14332 15020
rect 14004 14968 14056 14977
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 15568 15036 15620 15088
rect 19064 15036 19116 15088
rect 17224 14968 17276 15020
rect 17408 14968 17460 15020
rect 18328 14968 18380 15020
rect 18880 15011 18932 15020
rect 18880 14977 18898 15011
rect 18898 14977 18932 15011
rect 18880 14968 18932 14977
rect 7564 14900 7616 14909
rect 8116 14832 8168 14884
rect 7472 14764 7524 14816
rect 8208 14764 8260 14816
rect 8484 14764 8536 14816
rect 9036 14764 9088 14816
rect 9680 14832 9732 14884
rect 11152 14832 11204 14884
rect 12716 14832 12768 14884
rect 11336 14764 11388 14816
rect 12164 14764 12216 14816
rect 16028 14764 16080 14816
rect 17776 14807 17828 14816
rect 17776 14773 17785 14807
rect 17785 14773 17819 14807
rect 17819 14773 17828 14807
rect 17776 14764 17828 14773
rect 21548 15036 21600 15088
rect 20904 14968 20956 15020
rect 21272 15011 21324 15020
rect 21272 14977 21281 15011
rect 21281 14977 21315 15011
rect 21315 14977 21324 15011
rect 21272 14968 21324 14977
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 7104 14560 7156 14612
rect 7472 14560 7524 14612
rect 10416 14603 10468 14612
rect 4068 14492 4120 14544
rect 10416 14569 10425 14603
rect 10425 14569 10459 14603
rect 10459 14569 10468 14603
rect 10416 14560 10468 14569
rect 10784 14560 10836 14612
rect 11152 14560 11204 14612
rect 11888 14560 11940 14612
rect 10600 14492 10652 14544
rect 4252 14467 4304 14476
rect 1952 14356 2004 14408
rect 4252 14433 4261 14467
rect 4261 14433 4295 14467
rect 4295 14433 4304 14467
rect 4252 14424 4304 14433
rect 6092 14467 6144 14476
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2044 14263 2096 14272
rect 2044 14229 2053 14263
rect 2053 14229 2087 14263
rect 2087 14229 2096 14263
rect 2044 14220 2096 14229
rect 3792 14356 3844 14408
rect 4528 14356 4580 14408
rect 4896 14399 4948 14408
rect 4896 14365 4905 14399
rect 4905 14365 4939 14399
rect 4939 14365 4948 14399
rect 4896 14356 4948 14365
rect 2688 14220 2740 14272
rect 4804 14288 4856 14340
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 5172 14356 5224 14408
rect 7196 14424 7248 14476
rect 12348 14467 12400 14476
rect 12348 14433 12357 14467
rect 12357 14433 12391 14467
rect 12391 14433 12400 14467
rect 12348 14424 12400 14433
rect 5540 14288 5592 14340
rect 8484 14356 8536 14408
rect 11244 14356 11296 14408
rect 12900 14356 12952 14408
rect 13912 14560 13964 14612
rect 16212 14560 16264 14612
rect 15752 14492 15804 14544
rect 15568 14356 15620 14408
rect 17224 14399 17276 14408
rect 9312 14331 9364 14340
rect 5264 14263 5316 14272
rect 5264 14229 5273 14263
rect 5273 14229 5307 14263
rect 5307 14229 5316 14263
rect 5264 14220 5316 14229
rect 5448 14220 5500 14272
rect 5908 14220 5960 14272
rect 9312 14297 9346 14331
rect 9346 14297 9364 14331
rect 9312 14288 9364 14297
rect 7564 14263 7616 14272
rect 7564 14229 7573 14263
rect 7573 14229 7607 14263
rect 7607 14229 7616 14263
rect 7564 14220 7616 14229
rect 8576 14220 8628 14272
rect 9404 14220 9456 14272
rect 11060 14288 11112 14340
rect 11336 14288 11388 14340
rect 12072 14288 12124 14340
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 17408 14356 17460 14408
rect 17592 14356 17644 14408
rect 18144 14356 18196 14408
rect 18880 14560 18932 14612
rect 20168 14356 20220 14408
rect 20812 14399 20864 14408
rect 20812 14365 20821 14399
rect 20821 14365 20855 14399
rect 20855 14365 20864 14399
rect 20812 14356 20864 14365
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 13728 14263 13780 14272
rect 13728 14229 13737 14263
rect 13737 14229 13771 14263
rect 13771 14229 13780 14263
rect 13728 14220 13780 14229
rect 14004 14220 14056 14272
rect 17040 14288 17092 14340
rect 20444 14288 20496 14340
rect 17224 14220 17276 14272
rect 17316 14220 17368 14272
rect 17592 14220 17644 14272
rect 17960 14220 18012 14272
rect 18880 14263 18932 14272
rect 18880 14229 18889 14263
rect 18889 14229 18923 14263
rect 18923 14229 18932 14263
rect 18880 14220 18932 14229
rect 21272 14263 21324 14272
rect 21272 14229 21281 14263
rect 21281 14229 21315 14263
rect 21315 14229 21324 14263
rect 21272 14220 21324 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 3884 14016 3936 14068
rect 5448 14016 5500 14068
rect 7104 14059 7156 14068
rect 7104 14025 7113 14059
rect 7113 14025 7147 14059
rect 7147 14025 7156 14059
rect 7104 14016 7156 14025
rect 2780 13948 2832 14000
rect 4068 13948 4120 14000
rect 5908 13948 5960 14000
rect 9404 14016 9456 14068
rect 9772 14016 9824 14068
rect 10600 14016 10652 14068
rect 11152 14059 11204 14068
rect 11152 14025 11161 14059
rect 11161 14025 11195 14059
rect 11195 14025 11204 14059
rect 11152 14016 11204 14025
rect 12072 14016 12124 14068
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 19064 14016 19116 14068
rect 20444 14016 20496 14068
rect 7840 13948 7892 14000
rect 8852 13948 8904 14000
rect 10140 13948 10192 14000
rect 12348 13948 12400 14000
rect 2596 13923 2648 13932
rect 2596 13889 2605 13923
rect 2605 13889 2639 13923
rect 2639 13889 2648 13923
rect 2596 13880 2648 13889
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 4344 13923 4396 13932
rect 4344 13889 4353 13923
rect 4353 13889 4387 13923
rect 4387 13889 4396 13923
rect 4344 13880 4396 13889
rect 4620 13880 4672 13932
rect 5356 13880 5408 13932
rect 5724 13880 5776 13932
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 3332 13676 3384 13728
rect 5908 13812 5960 13864
rect 7196 13880 7248 13932
rect 7748 13880 7800 13932
rect 9312 13880 9364 13932
rect 7472 13812 7524 13864
rect 6000 13676 6052 13728
rect 9128 13744 9180 13796
rect 9312 13744 9364 13796
rect 8484 13676 8536 13728
rect 11060 13812 11112 13864
rect 12348 13812 12400 13864
rect 12716 13880 12768 13932
rect 13820 13880 13872 13932
rect 14004 13948 14056 14000
rect 17316 13948 17368 14000
rect 18052 13948 18104 14000
rect 20628 13991 20680 14000
rect 20628 13957 20646 13991
rect 20646 13957 20680 13991
rect 20628 13948 20680 13957
rect 15292 13923 15344 13932
rect 15292 13889 15310 13923
rect 15310 13889 15344 13923
rect 15292 13880 15344 13889
rect 16120 13880 16172 13932
rect 15568 13855 15620 13864
rect 15568 13821 15577 13855
rect 15577 13821 15611 13855
rect 15611 13821 15620 13855
rect 15568 13812 15620 13821
rect 19892 13812 19944 13864
rect 20904 13923 20956 13932
rect 20904 13889 20913 13923
rect 20913 13889 20947 13923
rect 20947 13889 20956 13923
rect 20904 13880 20956 13889
rect 21548 13880 21600 13932
rect 17868 13744 17920 13796
rect 19616 13744 19668 13796
rect 20904 13744 20956 13796
rect 21640 13744 21692 13796
rect 9496 13676 9548 13728
rect 11888 13676 11940 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 2504 13472 2556 13524
rect 2412 13404 2464 13456
rect 2688 13404 2740 13456
rect 3056 13472 3108 13524
rect 4344 13472 4396 13524
rect 6000 13472 6052 13524
rect 5632 13404 5684 13456
rect 10140 13472 10192 13524
rect 13820 13472 13872 13524
rect 15568 13472 15620 13524
rect 15844 13515 15896 13524
rect 15844 13481 15853 13515
rect 15853 13481 15887 13515
rect 15887 13481 15896 13515
rect 15844 13472 15896 13481
rect 18144 13472 18196 13524
rect 18420 13472 18472 13524
rect 18788 13472 18840 13524
rect 19064 13472 19116 13524
rect 19432 13472 19484 13524
rect 20812 13472 20864 13524
rect 20996 13472 21048 13524
rect 11704 13404 11756 13456
rect 11888 13404 11940 13456
rect 15292 13404 15344 13456
rect 20352 13447 20404 13456
rect 20352 13413 20361 13447
rect 20361 13413 20395 13447
rect 20395 13413 20404 13447
rect 20352 13404 20404 13413
rect 5724 13336 5776 13388
rect 6644 13336 6696 13388
rect 7012 13336 7064 13388
rect 3424 13268 3476 13320
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 3608 13200 3660 13252
rect 5264 13268 5316 13320
rect 7104 13268 7156 13320
rect 7656 13268 7708 13320
rect 8484 13336 8536 13388
rect 9956 13336 10008 13388
rect 15476 13336 15528 13388
rect 19616 13336 19668 13388
rect 20628 13336 20680 13388
rect 9036 13268 9088 13320
rect 10784 13268 10836 13320
rect 6000 13200 6052 13252
rect 7840 13200 7892 13252
rect 8208 13243 8260 13252
rect 8208 13209 8217 13243
rect 8217 13209 8251 13243
rect 8251 13209 8260 13243
rect 8208 13200 8260 13209
rect 8484 13200 8536 13252
rect 12624 13268 12676 13320
rect 16212 13268 16264 13320
rect 11152 13200 11204 13252
rect 17408 13268 17460 13320
rect 20260 13268 20312 13320
rect 2780 13132 2832 13184
rect 3792 13132 3844 13184
rect 4068 13132 4120 13184
rect 4896 13132 4948 13184
rect 5724 13132 5776 13184
rect 7656 13175 7708 13184
rect 7656 13141 7665 13175
rect 7665 13141 7699 13175
rect 7699 13141 7708 13175
rect 7656 13132 7708 13141
rect 9956 13132 10008 13184
rect 11060 13132 11112 13184
rect 11888 13132 11940 13184
rect 12440 13132 12492 13184
rect 12716 13132 12768 13184
rect 13084 13132 13136 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 18420 13200 18472 13252
rect 19524 13200 19576 13252
rect 18328 13132 18380 13184
rect 19892 13175 19944 13184
rect 19892 13141 19901 13175
rect 19901 13141 19935 13175
rect 19935 13141 19944 13175
rect 19892 13132 19944 13141
rect 20628 13132 20680 13184
rect 20812 13175 20864 13184
rect 20812 13141 20821 13175
rect 20821 13141 20855 13175
rect 20855 13141 20864 13175
rect 20812 13132 20864 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 2596 12928 2648 12980
rect 3424 12928 3476 12980
rect 3608 12971 3660 12980
rect 3608 12937 3617 12971
rect 3617 12937 3651 12971
rect 3651 12937 3660 12971
rect 3608 12928 3660 12937
rect 4528 12971 4580 12980
rect 4528 12937 4537 12971
rect 4537 12937 4571 12971
rect 4571 12937 4580 12971
rect 4528 12928 4580 12937
rect 4712 12928 4764 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 10784 12971 10836 12980
rect 1952 12835 2004 12844
rect 1952 12801 1961 12835
rect 1961 12801 1995 12835
rect 1995 12801 2004 12835
rect 1952 12792 2004 12801
rect 2044 12792 2096 12844
rect 7656 12860 7708 12912
rect 9772 12860 9824 12912
rect 10232 12903 10284 12912
rect 10232 12869 10250 12903
rect 10250 12869 10284 12903
rect 10232 12860 10284 12869
rect 3056 12792 3108 12844
rect 3516 12792 3568 12844
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 5080 12792 5132 12844
rect 5724 12792 5776 12844
rect 7840 12792 7892 12844
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 2872 12724 2924 12776
rect 3332 12724 3384 12776
rect 4344 12724 4396 12776
rect 5448 12724 5500 12776
rect 5540 12656 5592 12708
rect 3332 12631 3384 12640
rect 3332 12597 3341 12631
rect 3341 12597 3375 12631
rect 3375 12597 3384 12631
rect 3332 12588 3384 12597
rect 7288 12724 7340 12776
rect 6000 12656 6052 12708
rect 9312 12724 9364 12776
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 12624 12928 12676 12980
rect 13820 12903 13872 12912
rect 13820 12869 13829 12903
rect 13829 12869 13863 12903
rect 13863 12869 13872 12903
rect 13820 12860 13872 12869
rect 11152 12724 11204 12776
rect 11244 12724 11296 12776
rect 12348 12792 12400 12844
rect 15476 12928 15528 12980
rect 18512 12928 18564 12980
rect 18696 12928 18748 12980
rect 19432 12971 19484 12980
rect 17040 12860 17092 12912
rect 17224 12860 17276 12912
rect 18788 12860 18840 12912
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 20536 12928 20588 12980
rect 19616 12860 19668 12912
rect 14648 12767 14700 12776
rect 14648 12733 14657 12767
rect 14657 12733 14691 12767
rect 14691 12733 14700 12767
rect 17500 12792 17552 12844
rect 19984 12792 20036 12844
rect 14648 12724 14700 12733
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 6644 12588 6696 12597
rect 7104 12631 7156 12640
rect 7104 12597 7113 12631
rect 7113 12597 7147 12631
rect 7147 12597 7156 12631
rect 7104 12588 7156 12597
rect 8668 12588 8720 12640
rect 9496 12588 9548 12640
rect 13728 12656 13780 12708
rect 14280 12656 14332 12708
rect 18788 12724 18840 12776
rect 20536 12767 20588 12776
rect 20536 12733 20545 12767
rect 20545 12733 20579 12767
rect 20579 12733 20588 12767
rect 20536 12724 20588 12733
rect 19524 12656 19576 12708
rect 19984 12656 20036 12708
rect 16488 12588 16540 12640
rect 16580 12588 16632 12640
rect 17408 12588 17460 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 1676 12384 1728 12436
rect 4528 12384 4580 12436
rect 6828 12384 6880 12436
rect 8116 12384 8168 12436
rect 2872 12316 2924 12368
rect 8300 12316 8352 12368
rect 2136 12248 2188 12300
rect 2412 12248 2464 12300
rect 3148 12248 3200 12300
rect 2964 12180 3016 12232
rect 6000 12248 6052 12300
rect 4804 12180 4856 12232
rect 7104 12248 7156 12300
rect 10876 12384 10928 12436
rect 11612 12384 11664 12436
rect 11888 12384 11940 12436
rect 14464 12384 14516 12436
rect 16580 12427 16632 12436
rect 12164 12316 12216 12368
rect 13820 12316 13872 12368
rect 14648 12316 14700 12368
rect 13452 12248 13504 12300
rect 13728 12248 13780 12300
rect 16580 12393 16589 12427
rect 16589 12393 16623 12427
rect 16623 12393 16632 12427
rect 16580 12384 16632 12393
rect 17408 12384 17460 12436
rect 18144 12384 18196 12436
rect 19064 12384 19116 12436
rect 19800 12384 19852 12436
rect 20076 12384 20128 12436
rect 20352 12384 20404 12436
rect 20996 12384 21048 12436
rect 21180 12427 21232 12436
rect 21180 12393 21189 12427
rect 21189 12393 21223 12427
rect 21223 12393 21232 12427
rect 21180 12384 21232 12393
rect 16948 12316 17000 12368
rect 9128 12223 9180 12232
rect 2596 12044 2648 12096
rect 3240 12087 3292 12096
rect 3240 12053 3249 12087
rect 3249 12053 3283 12087
rect 3283 12053 3292 12087
rect 3240 12044 3292 12053
rect 4068 12044 4120 12096
rect 4344 12044 4396 12096
rect 5356 12087 5408 12096
rect 5356 12053 5365 12087
rect 5365 12053 5399 12087
rect 5399 12053 5408 12087
rect 5356 12044 5408 12053
rect 7196 12112 7248 12164
rect 7564 12112 7616 12164
rect 7932 12044 7984 12096
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9036 12112 9088 12164
rect 13268 12180 13320 12232
rect 13636 12180 13688 12232
rect 15384 12180 15436 12232
rect 21088 12316 21140 12368
rect 18788 12248 18840 12300
rect 9864 12112 9916 12164
rect 11612 12112 11664 12164
rect 12072 12112 12124 12164
rect 19892 12180 19944 12232
rect 20444 12248 20496 12300
rect 21272 12223 21324 12232
rect 21272 12189 21281 12223
rect 21281 12189 21315 12223
rect 21315 12189 21324 12223
rect 21272 12180 21324 12189
rect 10048 12044 10100 12096
rect 11060 12044 11112 12096
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 13360 12087 13412 12096
rect 13360 12053 13369 12087
rect 13369 12053 13403 12087
rect 13403 12053 13412 12087
rect 13360 12044 13412 12053
rect 15936 12112 15988 12164
rect 17224 12112 17276 12164
rect 17868 12112 17920 12164
rect 16028 12044 16080 12096
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 20168 12087 20220 12096
rect 20168 12053 20177 12087
rect 20177 12053 20211 12087
rect 20211 12053 20220 12087
rect 20168 12044 20220 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 1860 11840 1912 11892
rect 4068 11840 4120 11892
rect 4436 11840 4488 11892
rect 5080 11840 5132 11892
rect 6920 11883 6972 11892
rect 6920 11849 6929 11883
rect 6929 11849 6963 11883
rect 6963 11849 6972 11883
rect 6920 11840 6972 11849
rect 9772 11840 9824 11892
rect 2320 11772 2372 11824
rect 3240 11772 3292 11824
rect 4620 11772 4672 11824
rect 5356 11772 5408 11824
rect 5540 11772 5592 11824
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 5080 11704 5132 11756
rect 2228 11636 2280 11645
rect 2872 11636 2924 11688
rect 2412 11568 2464 11620
rect 3884 11568 3936 11620
rect 4620 11636 4672 11688
rect 5448 11636 5500 11688
rect 6736 11636 6788 11688
rect 7840 11704 7892 11756
rect 10876 11772 10928 11824
rect 17316 11840 17368 11892
rect 18052 11883 18104 11892
rect 18052 11849 18061 11883
rect 18061 11849 18095 11883
rect 18095 11849 18104 11883
rect 18052 11840 18104 11849
rect 18972 11840 19024 11892
rect 19800 11883 19852 11892
rect 19800 11849 19809 11883
rect 19809 11849 19843 11883
rect 19843 11849 19852 11883
rect 19800 11840 19852 11849
rect 20168 11883 20220 11892
rect 20168 11849 20177 11883
rect 20177 11849 20211 11883
rect 20211 11849 20220 11883
rect 20168 11840 20220 11849
rect 20812 11840 20864 11892
rect 12164 11772 12216 11824
rect 15844 11772 15896 11824
rect 16580 11704 16632 11756
rect 17776 11772 17828 11824
rect 7380 11679 7432 11688
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 7472 11636 7524 11688
rect 9036 11636 9088 11688
rect 10876 11679 10928 11688
rect 10876 11645 10878 11679
rect 10878 11645 10912 11679
rect 10912 11645 10928 11679
rect 10876 11636 10928 11645
rect 13636 11636 13688 11688
rect 14924 11679 14976 11688
rect 14924 11645 14933 11679
rect 14933 11645 14967 11679
rect 14967 11645 14976 11679
rect 14924 11636 14976 11645
rect 18236 11772 18288 11824
rect 17960 11704 18012 11756
rect 20260 11772 20312 11824
rect 20628 11772 20680 11824
rect 9864 11568 9916 11620
rect 6828 11500 6880 11552
rect 8116 11500 8168 11552
rect 8300 11543 8352 11552
rect 8300 11509 8309 11543
rect 8309 11509 8343 11543
rect 8343 11509 8352 11543
rect 8300 11500 8352 11509
rect 9496 11500 9548 11552
rect 13084 11568 13136 11620
rect 13268 11611 13320 11620
rect 13268 11577 13277 11611
rect 13277 11577 13311 11611
rect 13311 11577 13320 11611
rect 13268 11568 13320 11577
rect 21548 11704 21600 11756
rect 14648 11500 14700 11552
rect 14832 11500 14884 11552
rect 16212 11500 16264 11552
rect 16580 11500 16632 11552
rect 17408 11500 17460 11552
rect 17868 11500 17920 11552
rect 19064 11500 19116 11552
rect 20444 11636 20496 11688
rect 20720 11636 20772 11688
rect 20904 11679 20956 11688
rect 20904 11645 20913 11679
rect 20913 11645 20947 11679
rect 20947 11645 20956 11679
rect 20904 11636 20956 11645
rect 20536 11568 20588 11620
rect 21180 11500 21232 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1952 11296 2004 11348
rect 3332 11339 3384 11348
rect 3332 11305 3341 11339
rect 3341 11305 3375 11339
rect 3375 11305 3384 11339
rect 3332 11296 3384 11305
rect 3976 11339 4028 11348
rect 3976 11305 3985 11339
rect 3985 11305 4019 11339
rect 4019 11305 4028 11339
rect 3976 11296 4028 11305
rect 4160 11296 4212 11348
rect 6828 11296 6880 11348
rect 1676 11092 1728 11144
rect 2872 11160 2924 11212
rect 4344 11160 4396 11212
rect 5264 11160 5316 11212
rect 5724 11228 5776 11280
rect 8484 11296 8536 11348
rect 10416 11296 10468 11348
rect 10876 11339 10928 11348
rect 10876 11305 10885 11339
rect 10885 11305 10919 11339
rect 10919 11305 10928 11339
rect 10876 11296 10928 11305
rect 11888 11296 11940 11348
rect 12072 11296 12124 11348
rect 17040 11296 17092 11348
rect 17592 11339 17644 11348
rect 17592 11305 17601 11339
rect 17601 11305 17635 11339
rect 17635 11305 17644 11339
rect 17592 11296 17644 11305
rect 9128 11203 9180 11212
rect 9128 11169 9137 11203
rect 9137 11169 9171 11203
rect 9171 11169 9180 11203
rect 9128 11160 9180 11169
rect 2044 11067 2096 11076
rect 2044 11033 2053 11067
rect 2053 11033 2087 11067
rect 2087 11033 2096 11067
rect 2044 11024 2096 11033
rect 3332 11092 3384 11144
rect 7472 11092 7524 11144
rect 8208 11092 8260 11144
rect 9220 11092 9272 11144
rect 13820 11228 13872 11280
rect 18788 11296 18840 11348
rect 19984 11296 20036 11348
rect 22100 11296 22152 11348
rect 17960 11271 18012 11280
rect 17960 11237 17969 11271
rect 17969 11237 18003 11271
rect 18003 11237 18012 11271
rect 17960 11228 18012 11237
rect 18236 11228 18288 11280
rect 19524 11228 19576 11280
rect 10876 11160 10928 11212
rect 11244 11092 11296 11144
rect 19248 11160 19300 11212
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 19156 11092 19208 11144
rect 20996 11160 21048 11212
rect 3884 11067 3936 11076
rect 3884 11033 3893 11067
rect 3893 11033 3927 11067
rect 3927 11033 3936 11067
rect 3884 11024 3936 11033
rect 4896 11067 4948 11076
rect 4896 11033 4905 11067
rect 4905 11033 4939 11067
rect 4939 11033 4948 11067
rect 4896 11024 4948 11033
rect 1952 10999 2004 11008
rect 1952 10965 1961 10999
rect 1961 10965 1995 10999
rect 1995 10965 2004 10999
rect 1952 10956 2004 10965
rect 2964 10999 3016 11008
rect 2964 10965 2973 10999
rect 2973 10965 3007 10999
rect 3007 10965 3016 10999
rect 2964 10956 3016 10965
rect 4160 10956 4212 11008
rect 4436 10956 4488 11008
rect 6920 11024 6972 11076
rect 9588 11024 9640 11076
rect 5080 10956 5132 11008
rect 5632 10999 5684 11008
rect 5632 10965 5641 10999
rect 5641 10965 5675 10999
rect 5675 10965 5684 10999
rect 5632 10956 5684 10965
rect 7104 10956 7156 11008
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 10232 10956 10284 11008
rect 12072 10956 12124 11008
rect 14924 10956 14976 11008
rect 17040 10956 17092 11008
rect 20536 11024 20588 11076
rect 21272 11067 21324 11076
rect 21272 11033 21281 11067
rect 21281 11033 21315 11067
rect 21315 11033 21324 11067
rect 21272 11024 21324 11033
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 1400 10752 1452 10804
rect 4068 10752 4120 10804
rect 5448 10752 5500 10804
rect 6000 10752 6052 10804
rect 6276 10752 6328 10804
rect 10876 10795 10928 10804
rect 3148 10684 3200 10736
rect 3884 10684 3936 10736
rect 6460 10684 6512 10736
rect 6644 10684 6696 10736
rect 7288 10684 7340 10736
rect 7472 10684 7524 10736
rect 8300 10684 8352 10736
rect 10140 10684 10192 10736
rect 10600 10684 10652 10736
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 11060 10684 11112 10736
rect 1584 10616 1636 10668
rect 2964 10591 3016 10600
rect 2964 10557 2973 10591
rect 2973 10557 3007 10591
rect 3007 10557 3016 10591
rect 2964 10548 3016 10557
rect 3056 10591 3108 10600
rect 3056 10557 3065 10591
rect 3065 10557 3099 10591
rect 3099 10557 3108 10591
rect 5540 10616 5592 10668
rect 6000 10616 6052 10668
rect 8024 10616 8076 10668
rect 9864 10616 9916 10668
rect 3056 10548 3108 10557
rect 4896 10548 4948 10600
rect 5264 10548 5316 10600
rect 10876 10616 10928 10668
rect 2780 10480 2832 10532
rect 8484 10480 8536 10532
rect 2136 10412 2188 10464
rect 5172 10412 5224 10464
rect 7104 10412 7156 10464
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 10784 10548 10836 10600
rect 13820 10684 13872 10736
rect 14372 10752 14424 10804
rect 17408 10795 17460 10804
rect 17408 10761 17417 10795
rect 17417 10761 17451 10795
rect 17451 10761 17460 10795
rect 17408 10752 17460 10761
rect 18604 10752 18656 10804
rect 20536 10795 20588 10804
rect 14556 10684 14608 10736
rect 15016 10684 15068 10736
rect 17040 10684 17092 10736
rect 19616 10684 19668 10736
rect 20536 10761 20545 10795
rect 20545 10761 20579 10795
rect 20579 10761 20588 10795
rect 20536 10752 20588 10761
rect 18236 10616 18288 10668
rect 19156 10659 19208 10668
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 19248 10616 19300 10668
rect 21272 10659 21324 10668
rect 21272 10625 21281 10659
rect 21281 10625 21315 10659
rect 21315 10625 21324 10659
rect 21272 10616 21324 10625
rect 13176 10523 13228 10532
rect 13176 10489 13185 10523
rect 13185 10489 13219 10523
rect 13219 10489 13228 10523
rect 13176 10480 13228 10489
rect 15844 10548 15896 10600
rect 16304 10548 16356 10600
rect 12440 10455 12492 10464
rect 12440 10421 12449 10455
rect 12449 10421 12483 10455
rect 12483 10421 12492 10455
rect 14924 10455 14976 10464
rect 12440 10412 12492 10421
rect 14924 10421 14933 10455
rect 14933 10421 14967 10455
rect 14967 10421 14976 10455
rect 14924 10412 14976 10421
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 1952 10208 2004 10260
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 4896 10251 4948 10260
rect 4896 10217 4905 10251
rect 4905 10217 4939 10251
rect 4939 10217 4948 10251
rect 4896 10208 4948 10217
rect 6552 10208 6604 10260
rect 6736 10208 6788 10260
rect 7288 10208 7340 10260
rect 9220 10208 9272 10260
rect 1584 10140 1636 10192
rect 2136 10115 2188 10124
rect 2136 10081 2145 10115
rect 2145 10081 2179 10115
rect 2179 10081 2188 10115
rect 2136 10072 2188 10081
rect 5356 10140 5408 10192
rect 5540 10140 5592 10192
rect 2412 10072 2464 10124
rect 3424 10072 3476 10124
rect 4160 10072 4212 10124
rect 4344 10115 4396 10124
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 5724 10115 5776 10124
rect 5724 10081 5733 10115
rect 5733 10081 5767 10115
rect 5767 10081 5776 10115
rect 5724 10072 5776 10081
rect 7472 10140 7524 10192
rect 6828 10115 6880 10124
rect 3148 10004 3200 10056
rect 3240 10047 3292 10056
rect 3240 10013 3249 10047
rect 3249 10013 3283 10047
rect 3283 10013 3292 10047
rect 3240 10004 3292 10013
rect 3976 10004 4028 10056
rect 5448 10004 5500 10056
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 8024 10072 8076 10081
rect 8484 10004 8536 10056
rect 10876 10208 10928 10260
rect 13820 10208 13872 10260
rect 14280 10208 14332 10260
rect 14832 10251 14884 10260
rect 14832 10217 14841 10251
rect 14841 10217 14875 10251
rect 14875 10217 14884 10251
rect 14832 10208 14884 10217
rect 11244 10004 11296 10056
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 14372 10072 14424 10124
rect 17132 10208 17184 10260
rect 16948 10140 17000 10192
rect 17868 10208 17920 10260
rect 18236 10208 18288 10260
rect 18512 10208 18564 10260
rect 17224 10072 17276 10124
rect 19064 10072 19116 10124
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 20536 10115 20588 10124
rect 20536 10081 20545 10115
rect 20545 10081 20579 10115
rect 20579 10081 20588 10115
rect 20536 10072 20588 10081
rect 13820 10004 13872 10056
rect 14924 10004 14976 10056
rect 2780 9979 2832 9988
rect 2780 9945 2789 9979
rect 2789 9945 2823 9979
rect 2823 9945 2832 9979
rect 2780 9936 2832 9945
rect 5908 9936 5960 9988
rect 6276 9936 6328 9988
rect 7472 9979 7524 9988
rect 7472 9945 7481 9979
rect 7481 9945 7515 9979
rect 7515 9945 7524 9979
rect 8208 9979 8260 9988
rect 7472 9936 7524 9945
rect 8208 9945 8217 9979
rect 8217 9945 8251 9979
rect 8251 9945 8260 9979
rect 8208 9936 8260 9945
rect 10048 9979 10100 9988
rect 10048 9945 10066 9979
rect 10066 9945 10100 9979
rect 10048 9936 10100 9945
rect 2872 9868 2924 9920
rect 4160 9868 4212 9920
rect 4252 9868 4304 9920
rect 4896 9868 4948 9920
rect 5264 9911 5316 9920
rect 5264 9877 5273 9911
rect 5273 9877 5307 9911
rect 5307 9877 5316 9911
rect 5264 9868 5316 9877
rect 8300 9868 8352 9920
rect 11704 9868 11756 9920
rect 11980 9868 12032 9920
rect 13268 9936 13320 9988
rect 14464 9936 14516 9988
rect 13820 9868 13872 9920
rect 14832 9868 14884 9920
rect 15844 9936 15896 9988
rect 20076 10004 20128 10056
rect 20168 9979 20220 9988
rect 17316 9868 17368 9920
rect 18144 9868 18196 9920
rect 20168 9945 20177 9979
rect 20177 9945 20211 9979
rect 20211 9945 20220 9979
rect 20168 9936 20220 9945
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 4160 9664 4212 9716
rect 9496 9664 9548 9716
rect 10876 9707 10928 9716
rect 10876 9673 10885 9707
rect 10885 9673 10919 9707
rect 10919 9673 10928 9707
rect 10876 9664 10928 9673
rect 11060 9664 11112 9716
rect 11796 9664 11848 9716
rect 12440 9664 12492 9716
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 2320 9460 2372 9512
rect 2964 9596 3016 9648
rect 4068 9596 4120 9648
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3884 9571 3936 9580
rect 1860 9392 1912 9444
rect 3884 9537 3893 9571
rect 3893 9537 3927 9571
rect 3927 9537 3936 9571
rect 3884 9528 3936 9537
rect 3700 9460 3752 9512
rect 5080 9596 5132 9648
rect 5724 9596 5776 9648
rect 8576 9596 8628 9648
rect 9128 9596 9180 9648
rect 9220 9596 9272 9648
rect 4436 9528 4488 9580
rect 5356 9528 5408 9580
rect 5448 9528 5500 9580
rect 6000 9528 6052 9580
rect 6828 9528 6880 9580
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 5632 9460 5684 9512
rect 4528 9392 4580 9444
rect 8300 9460 8352 9512
rect 10784 9596 10836 9648
rect 9128 9460 9180 9512
rect 12348 9528 12400 9580
rect 13084 9528 13136 9580
rect 17500 9596 17552 9648
rect 20168 9664 20220 9716
rect 20444 9664 20496 9716
rect 17868 9528 17920 9580
rect 18236 9528 18288 9580
rect 19616 9528 19668 9580
rect 20536 9571 20588 9580
rect 20536 9537 20545 9571
rect 20545 9537 20579 9571
rect 20579 9537 20588 9571
rect 20536 9528 20588 9537
rect 2596 9324 2648 9376
rect 2780 9367 2832 9376
rect 2780 9333 2789 9367
rect 2789 9333 2823 9367
rect 2823 9333 2832 9367
rect 2780 9324 2832 9333
rect 2964 9324 3016 9376
rect 3516 9324 3568 9376
rect 5540 9367 5592 9376
rect 5540 9333 5549 9367
rect 5549 9333 5583 9367
rect 5583 9333 5592 9367
rect 5540 9324 5592 9333
rect 6000 9324 6052 9376
rect 7288 9324 7340 9376
rect 7472 9324 7524 9376
rect 11704 9392 11756 9444
rect 12072 9392 12124 9444
rect 13820 9460 13872 9512
rect 17500 9503 17552 9512
rect 17500 9469 17509 9503
rect 17509 9469 17543 9503
rect 17543 9469 17552 9503
rect 17500 9460 17552 9469
rect 17592 9503 17644 9512
rect 17592 9469 17601 9503
rect 17601 9469 17635 9503
rect 17635 9469 17644 9503
rect 19708 9503 19760 9512
rect 17592 9460 17644 9469
rect 19708 9469 19717 9503
rect 19717 9469 19751 9503
rect 19751 9469 19760 9503
rect 19708 9460 19760 9469
rect 20812 9503 20864 9512
rect 20812 9469 20821 9503
rect 20821 9469 20855 9503
rect 20855 9469 20864 9503
rect 20812 9460 20864 9469
rect 13544 9435 13596 9444
rect 13544 9401 13553 9435
rect 13553 9401 13587 9435
rect 13587 9401 13596 9435
rect 13544 9392 13596 9401
rect 15476 9392 15528 9444
rect 17684 9392 17736 9444
rect 19892 9392 19944 9444
rect 9404 9324 9456 9376
rect 10600 9367 10652 9376
rect 10600 9333 10609 9367
rect 10609 9333 10643 9367
rect 10643 9333 10652 9367
rect 10600 9324 10652 9333
rect 12992 9324 13044 9376
rect 13452 9324 13504 9376
rect 15568 9367 15620 9376
rect 15568 9333 15577 9367
rect 15577 9333 15611 9367
rect 15611 9333 15620 9367
rect 15568 9324 15620 9333
rect 16212 9324 16264 9376
rect 19984 9324 20036 9376
rect 20628 9324 20680 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 1768 8984 1820 9036
rect 5724 9120 5776 9172
rect 7012 9120 7064 9172
rect 8024 9120 8076 9172
rect 9220 9120 9272 9172
rect 9588 9120 9640 9172
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 2412 8848 2464 8900
rect 3056 9052 3108 9104
rect 4528 9052 4580 9104
rect 5356 9052 5408 9104
rect 7564 9052 7616 9104
rect 8484 9052 8536 9104
rect 9036 9052 9088 9104
rect 10876 9120 10928 9172
rect 11244 9120 11296 9172
rect 16304 9120 16356 9172
rect 17224 9120 17276 9172
rect 19800 9163 19852 9172
rect 11152 9052 11204 9104
rect 11520 9095 11572 9104
rect 11520 9061 11529 9095
rect 11529 9061 11563 9095
rect 11563 9061 11572 9095
rect 11520 9052 11572 9061
rect 14280 9052 14332 9104
rect 17776 9052 17828 9104
rect 3148 9027 3200 9036
rect 3148 8993 3157 9027
rect 3157 8993 3191 9027
rect 3191 8993 3200 9027
rect 3148 8984 3200 8993
rect 4436 8984 4488 9036
rect 6828 8984 6880 9036
rect 4896 8916 4948 8968
rect 5540 8916 5592 8968
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 10876 8984 10928 9036
rect 15568 9027 15620 9036
rect 15568 8993 15577 9027
rect 15577 8993 15611 9027
rect 15611 8993 15620 9027
rect 15568 8984 15620 8993
rect 10600 8916 10652 8968
rect 11520 8916 11572 8968
rect 14556 8916 14608 8968
rect 15660 8916 15712 8968
rect 17960 8916 18012 8968
rect 3148 8848 3200 8900
rect 3792 8848 3844 8900
rect 4252 8780 4304 8832
rect 9680 8848 9732 8900
rect 10140 8848 10192 8900
rect 11980 8848 12032 8900
rect 12348 8848 12400 8900
rect 12808 8848 12860 8900
rect 13452 8848 13504 8900
rect 15292 8891 15344 8900
rect 15292 8857 15310 8891
rect 15310 8857 15344 8891
rect 15292 8848 15344 8857
rect 5080 8780 5132 8832
rect 5724 8780 5776 8832
rect 7288 8780 7340 8832
rect 9220 8780 9272 8832
rect 9496 8780 9548 8832
rect 17040 8848 17092 8900
rect 17224 8891 17276 8900
rect 17224 8857 17242 8891
rect 17242 8857 17276 8891
rect 17224 8848 17276 8857
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 19064 8916 19116 8968
rect 19800 9129 19809 9163
rect 19809 9129 19843 9163
rect 19843 9129 19852 9163
rect 19800 9120 19852 9129
rect 20168 8984 20220 9036
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 19340 8848 19392 8900
rect 21088 8891 21140 8900
rect 18696 8823 18748 8832
rect 16120 8780 16172 8789
rect 18696 8789 18705 8823
rect 18705 8789 18739 8823
rect 18739 8789 18748 8823
rect 18696 8780 18748 8789
rect 20168 8823 20220 8832
rect 20168 8789 20177 8823
rect 20177 8789 20211 8823
rect 20211 8789 20220 8823
rect 20168 8780 20220 8789
rect 20260 8823 20312 8832
rect 20260 8789 20269 8823
rect 20269 8789 20303 8823
rect 20303 8789 20312 8823
rect 21088 8857 21097 8891
rect 21097 8857 21131 8891
rect 21131 8857 21140 8891
rect 21088 8848 21140 8857
rect 20260 8780 20312 8789
rect 20536 8780 20588 8832
rect 21364 8780 21416 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 2136 8576 2188 8628
rect 3976 8576 4028 8628
rect 6644 8576 6696 8628
rect 8760 8619 8812 8628
rect 8760 8585 8769 8619
rect 8769 8585 8803 8619
rect 8803 8585 8812 8619
rect 8760 8576 8812 8585
rect 9128 8619 9180 8628
rect 5356 8508 5408 8560
rect 7196 8508 7248 8560
rect 8208 8551 8260 8560
rect 8208 8517 8217 8551
rect 8217 8517 8251 8551
rect 8251 8517 8260 8551
rect 8208 8508 8260 8517
rect 1492 8440 1544 8492
rect 4712 8440 4764 8492
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 3148 8415 3200 8424
rect 3148 8381 3157 8415
rect 3157 8381 3191 8415
rect 3191 8381 3200 8415
rect 3148 8372 3200 8381
rect 4160 8372 4212 8424
rect 4252 8372 4304 8424
rect 5448 8483 5500 8492
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 5632 8440 5684 8492
rect 5540 8372 5592 8424
rect 8300 8372 8352 8424
rect 2688 8304 2740 8356
rect 3792 8304 3844 8356
rect 3976 8304 4028 8356
rect 6644 8304 6696 8356
rect 7288 8304 7340 8356
rect 9128 8585 9137 8619
rect 9137 8585 9171 8619
rect 9171 8585 9180 8619
rect 9128 8576 9180 8585
rect 9496 8576 9548 8628
rect 9312 8508 9364 8560
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9772 8508 9824 8560
rect 10048 8576 10100 8628
rect 12256 8576 12308 8628
rect 13360 8576 13412 8628
rect 16120 8576 16172 8628
rect 16304 8576 16356 8628
rect 17500 8576 17552 8628
rect 20444 8619 20496 8628
rect 20444 8585 20453 8619
rect 20453 8585 20487 8619
rect 20487 8585 20496 8619
rect 20444 8576 20496 8585
rect 15200 8508 15252 8560
rect 15292 8508 15344 8560
rect 17224 8508 17276 8560
rect 17408 8508 17460 8560
rect 17684 8508 17736 8560
rect 18236 8508 18288 8560
rect 18328 8551 18380 8560
rect 18328 8517 18337 8551
rect 18337 8517 18371 8551
rect 18371 8517 18380 8551
rect 18696 8551 18748 8560
rect 18328 8508 18380 8517
rect 18696 8517 18705 8551
rect 18705 8517 18739 8551
rect 18739 8517 18748 8551
rect 18696 8508 18748 8517
rect 19340 8508 19392 8560
rect 19524 8508 19576 8560
rect 21364 8508 21416 8560
rect 9404 8440 9456 8449
rect 9404 8304 9456 8356
rect 13268 8440 13320 8492
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 19064 8440 19116 8492
rect 13544 8372 13596 8424
rect 6552 8236 6604 8288
rect 9128 8236 9180 8288
rect 10784 8236 10836 8288
rect 11152 8279 11204 8288
rect 11152 8245 11161 8279
rect 11161 8245 11195 8279
rect 11195 8245 11204 8279
rect 11152 8236 11204 8245
rect 18696 8372 18748 8424
rect 19892 8440 19944 8492
rect 20720 8440 20772 8492
rect 20628 8415 20680 8424
rect 20628 8381 20637 8415
rect 20637 8381 20671 8415
rect 20671 8381 20680 8415
rect 20628 8372 20680 8381
rect 15384 8347 15436 8356
rect 15384 8313 15393 8347
rect 15393 8313 15427 8347
rect 15427 8313 15436 8347
rect 15384 8304 15436 8313
rect 21088 8347 21140 8356
rect 21088 8313 21097 8347
rect 21097 8313 21131 8347
rect 21131 8313 21140 8347
rect 21088 8304 21140 8313
rect 16120 8236 16172 8288
rect 17040 8236 17092 8288
rect 19064 8236 19116 8288
rect 19708 8236 19760 8288
rect 20444 8236 20496 8288
rect 20628 8236 20680 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 2320 8032 2372 8084
rect 3884 8032 3936 8084
rect 5908 8075 5960 8084
rect 5908 8041 5917 8075
rect 5917 8041 5951 8075
rect 5951 8041 5960 8075
rect 5908 8032 5960 8041
rect 6828 8032 6880 8084
rect 8668 8032 8720 8084
rect 9680 8032 9732 8084
rect 18696 8032 18748 8084
rect 20996 8032 21048 8084
rect 21456 8032 21508 8084
rect 2964 7964 3016 8016
rect 3332 8007 3384 8016
rect 3332 7973 3341 8007
rect 3341 7973 3375 8007
rect 3375 7973 3384 8007
rect 3332 7964 3384 7973
rect 1676 7896 1728 7948
rect 2412 7896 2464 7948
rect 5172 7939 5224 7948
rect 2872 7828 2924 7880
rect 3240 7828 3292 7880
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 4620 7828 4672 7880
rect 5172 7905 5181 7939
rect 5181 7905 5215 7939
rect 5215 7905 5224 7939
rect 5172 7896 5224 7905
rect 5724 7896 5776 7948
rect 7012 7896 7064 7948
rect 7288 7896 7340 7948
rect 9772 7964 9824 8016
rect 15108 7964 15160 8016
rect 18788 7964 18840 8016
rect 19524 7964 19576 8016
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 6000 7828 6052 7880
rect 7380 7828 7432 7880
rect 12716 7939 12768 7948
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 8300 7828 8352 7880
rect 10048 7828 10100 7880
rect 10692 7828 10744 7880
rect 11152 7828 11204 7880
rect 7564 7760 7616 7812
rect 12716 7905 12725 7939
rect 12725 7905 12759 7939
rect 12759 7905 12768 7939
rect 12716 7896 12768 7905
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 1860 7692 1912 7744
rect 2136 7692 2188 7744
rect 4344 7692 4396 7744
rect 5816 7692 5868 7744
rect 6736 7692 6788 7744
rect 6828 7735 6880 7744
rect 6828 7701 6837 7735
rect 6837 7701 6871 7735
rect 6871 7701 6880 7735
rect 8208 7735 8260 7744
rect 6828 7692 6880 7701
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 9680 7692 9732 7744
rect 11152 7735 11204 7744
rect 11152 7701 11161 7735
rect 11161 7701 11195 7735
rect 11195 7701 11204 7735
rect 11152 7692 11204 7701
rect 14280 7760 14332 7812
rect 17132 7871 17184 7880
rect 17132 7837 17166 7871
rect 17166 7837 17184 7871
rect 16120 7803 16172 7812
rect 13636 7692 13688 7744
rect 16120 7769 16129 7803
rect 16129 7769 16163 7803
rect 16163 7769 16172 7803
rect 16120 7760 16172 7769
rect 17132 7828 17184 7837
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 20628 7828 20680 7880
rect 17040 7760 17092 7812
rect 17868 7760 17920 7812
rect 14924 7692 14976 7744
rect 15844 7692 15896 7744
rect 16028 7692 16080 7744
rect 17960 7692 18012 7744
rect 18328 7692 18380 7744
rect 19524 7692 19576 7744
rect 20536 7760 20588 7812
rect 21272 7803 21324 7812
rect 21272 7769 21281 7803
rect 21281 7769 21315 7803
rect 21315 7769 21324 7803
rect 21272 7760 21324 7769
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 664 7488 716 7540
rect 1124 7488 1176 7540
rect 1860 7531 1912 7540
rect 1860 7497 1869 7531
rect 1869 7497 1903 7531
rect 1903 7497 1912 7531
rect 1860 7488 1912 7497
rect 2044 7488 2096 7540
rect 2596 7488 2648 7540
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 5356 7488 5408 7540
rect 6552 7488 6604 7540
rect 9312 7531 9364 7540
rect 9312 7497 9321 7531
rect 9321 7497 9355 7531
rect 9355 7497 9364 7531
rect 9312 7488 9364 7497
rect 9404 7488 9456 7540
rect 12164 7488 12216 7540
rect 14648 7488 14700 7540
rect 940 7352 992 7404
rect 1124 7352 1176 7404
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 1584 7284 1636 7336
rect 2872 7284 2924 7336
rect 4436 7352 4488 7404
rect 4988 7352 5040 7404
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 7840 7420 7892 7472
rect 12348 7420 12400 7472
rect 6644 7284 6696 7336
rect 8392 7352 8444 7404
rect 10600 7352 10652 7404
rect 11980 7352 12032 7404
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 14648 7395 14700 7404
rect 14648 7361 14657 7395
rect 14657 7361 14691 7395
rect 14691 7361 14700 7395
rect 14648 7352 14700 7361
rect 8576 7284 8628 7336
rect 9312 7284 9364 7336
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 11152 7284 11204 7336
rect 15752 7352 15804 7404
rect 17040 7352 17092 7404
rect 17132 7352 17184 7404
rect 20260 7488 20312 7540
rect 20720 7488 20772 7540
rect 18880 7420 18932 7472
rect 2596 7216 2648 7268
rect 7196 7216 7248 7268
rect 8392 7216 8444 7268
rect 3424 7148 3476 7200
rect 6368 7191 6420 7200
rect 6368 7157 6377 7191
rect 6377 7157 6411 7191
rect 6411 7157 6420 7191
rect 6368 7148 6420 7157
rect 7012 7148 7064 7200
rect 9496 7216 9548 7268
rect 12624 7259 12676 7268
rect 10784 7148 10836 7200
rect 11152 7148 11204 7200
rect 12624 7225 12633 7259
rect 12633 7225 12667 7259
rect 12667 7225 12676 7259
rect 12624 7216 12676 7225
rect 17224 7284 17276 7336
rect 21180 7420 21232 7472
rect 18420 7327 18472 7336
rect 18420 7293 18429 7327
rect 18429 7293 18463 7327
rect 18463 7293 18472 7327
rect 18420 7284 18472 7293
rect 18972 7284 19024 7336
rect 20628 7284 20680 7336
rect 21272 7327 21324 7336
rect 21272 7293 21281 7327
rect 21281 7293 21315 7327
rect 21315 7293 21324 7327
rect 21272 7284 21324 7293
rect 12072 7148 12124 7200
rect 12440 7148 12492 7200
rect 13452 7148 13504 7200
rect 16120 7216 16172 7268
rect 17960 7216 18012 7268
rect 17868 7148 17920 7200
rect 18788 7148 18840 7200
rect 20536 7148 20588 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 1952 6944 2004 6996
rect 2688 6944 2740 6996
rect 7380 6987 7432 6996
rect 2320 6851 2372 6860
rect 2320 6817 2329 6851
rect 2329 6817 2363 6851
rect 2363 6817 2372 6851
rect 2320 6808 2372 6817
rect 5356 6876 5408 6928
rect 7380 6953 7389 6987
rect 7389 6953 7423 6987
rect 7423 6953 7432 6987
rect 7380 6944 7432 6953
rect 7564 6944 7616 6996
rect 2780 6740 2832 6792
rect 6736 6808 6788 6860
rect 6368 6740 6420 6792
rect 6644 6740 6696 6792
rect 9404 6876 9456 6928
rect 7288 6808 7340 6860
rect 8576 6808 8628 6860
rect 8668 6808 8720 6860
rect 10692 6808 10744 6860
rect 9772 6740 9824 6792
rect 12072 6944 12124 6996
rect 14464 6944 14516 6996
rect 14648 6944 14700 6996
rect 17040 6944 17092 6996
rect 17868 6944 17920 6996
rect 21272 6944 21324 6996
rect 12808 6808 12860 6860
rect 14280 6808 14332 6860
rect 15568 6808 15620 6860
rect 15844 6808 15896 6860
rect 16120 6851 16172 6860
rect 16120 6817 16129 6851
rect 16129 6817 16163 6851
rect 16163 6817 16172 6851
rect 16120 6808 16172 6817
rect 16304 6808 16356 6860
rect 17408 6851 17460 6860
rect 10968 6740 11020 6792
rect 11060 6740 11112 6792
rect 14832 6740 14884 6792
rect 15108 6740 15160 6792
rect 17408 6817 17417 6851
rect 17417 6817 17451 6851
rect 17451 6817 17460 6851
rect 17408 6808 17460 6817
rect 17592 6876 17644 6928
rect 18236 6808 18288 6860
rect 18420 6808 18472 6860
rect 20904 6808 20956 6860
rect 20628 6783 20680 6792
rect 3424 6672 3476 6724
rect 4620 6672 4672 6724
rect 4896 6672 4948 6724
rect 2136 6647 2188 6656
rect 2136 6613 2145 6647
rect 2145 6613 2179 6647
rect 2179 6613 2188 6647
rect 2136 6604 2188 6613
rect 2688 6647 2740 6656
rect 2688 6613 2697 6647
rect 2697 6613 2731 6647
rect 2731 6613 2740 6647
rect 2688 6604 2740 6613
rect 3148 6647 3200 6656
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3792 6647 3844 6656
rect 3148 6604 3200 6613
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 5080 6647 5132 6656
rect 4252 6604 4304 6613
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 7380 6672 7432 6724
rect 7748 6647 7800 6656
rect 7748 6613 7757 6647
rect 7757 6613 7791 6647
rect 7791 6613 7800 6647
rect 7748 6604 7800 6613
rect 8208 6604 8260 6656
rect 9864 6672 9916 6724
rect 10140 6604 10192 6656
rect 11980 6604 12032 6656
rect 12164 6715 12216 6724
rect 12164 6681 12182 6715
rect 12182 6681 12216 6715
rect 12164 6672 12216 6681
rect 12348 6672 12400 6724
rect 15384 6672 15436 6724
rect 20628 6749 20637 6783
rect 20637 6749 20671 6783
rect 20671 6749 20680 6783
rect 20628 6740 20680 6749
rect 17500 6672 17552 6724
rect 12532 6604 12584 6656
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 13084 6647 13136 6656
rect 13084 6613 13093 6647
rect 13093 6613 13127 6647
rect 13127 6613 13136 6647
rect 13084 6604 13136 6613
rect 13636 6647 13688 6656
rect 13636 6613 13645 6647
rect 13645 6613 13679 6647
rect 13679 6613 13688 6647
rect 13636 6604 13688 6613
rect 14832 6604 14884 6656
rect 15016 6647 15068 6656
rect 15016 6613 15025 6647
rect 15025 6613 15059 6647
rect 15059 6613 15068 6647
rect 15016 6604 15068 6613
rect 16212 6647 16264 6656
rect 16212 6613 16221 6647
rect 16221 6613 16255 6647
rect 16255 6613 16264 6647
rect 16212 6604 16264 6613
rect 16580 6647 16632 6656
rect 16580 6613 16589 6647
rect 16589 6613 16623 6647
rect 16623 6613 16632 6647
rect 16580 6604 16632 6613
rect 16948 6604 17000 6656
rect 17592 6647 17644 6656
rect 17592 6613 17601 6647
rect 17601 6613 17635 6647
rect 17635 6613 17644 6647
rect 19616 6672 19668 6724
rect 20536 6672 20588 6724
rect 17592 6604 17644 6613
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 19248 6647 19300 6656
rect 19248 6613 19257 6647
rect 19257 6613 19291 6647
rect 19291 6613 19300 6647
rect 19248 6604 19300 6613
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 2136 6400 2188 6452
rect 3148 6400 3200 6452
rect 3884 6400 3936 6452
rect 4988 6400 5040 6452
rect 5356 6400 5408 6452
rect 6552 6443 6604 6452
rect 1492 6375 1544 6384
rect 1492 6341 1501 6375
rect 1501 6341 1535 6375
rect 1535 6341 1544 6375
rect 1492 6332 1544 6341
rect 1676 6332 1728 6384
rect 6276 6332 6328 6384
rect 2136 6264 2188 6316
rect 2964 6264 3016 6316
rect 4436 6307 4488 6316
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 4804 6264 4856 6316
rect 4988 6307 5040 6316
rect 4988 6273 4997 6307
rect 4997 6273 5031 6307
rect 5031 6273 5040 6307
rect 4988 6264 5040 6273
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 6552 6409 6561 6443
rect 6561 6409 6595 6443
rect 6595 6409 6604 6443
rect 6552 6400 6604 6409
rect 7104 6443 7156 6452
rect 7104 6409 7113 6443
rect 7113 6409 7147 6443
rect 7147 6409 7156 6443
rect 7104 6400 7156 6409
rect 7564 6332 7616 6384
rect 8116 6375 8168 6384
rect 7288 6264 7340 6316
rect 1768 6128 1820 6180
rect 3056 6196 3108 6248
rect 4620 6239 4672 6248
rect 4620 6205 4629 6239
rect 4629 6205 4663 6239
rect 4663 6205 4672 6239
rect 4620 6196 4672 6205
rect 5172 6171 5224 6180
rect 5172 6137 5181 6171
rect 5181 6137 5215 6171
rect 5215 6137 5224 6171
rect 5172 6128 5224 6137
rect 7380 6196 7432 6248
rect 7564 6239 7616 6248
rect 7564 6205 7573 6239
rect 7573 6205 7607 6239
rect 7607 6205 7616 6239
rect 7564 6196 7616 6205
rect 8116 6341 8125 6375
rect 8125 6341 8159 6375
rect 8159 6341 8168 6375
rect 8116 6332 8168 6341
rect 9128 6332 9180 6384
rect 9404 6332 9456 6384
rect 9772 6400 9824 6452
rect 12072 6400 12124 6452
rect 12808 6400 12860 6452
rect 12992 6443 13044 6452
rect 12992 6409 13001 6443
rect 13001 6409 13035 6443
rect 13035 6409 13044 6443
rect 12992 6400 13044 6409
rect 14556 6400 14608 6452
rect 17224 6400 17276 6452
rect 20904 6400 20956 6452
rect 8576 6264 8628 6316
rect 11704 6332 11756 6384
rect 14280 6332 14332 6384
rect 15016 6332 15068 6384
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 12808 6264 12860 6316
rect 14464 6264 14516 6316
rect 16028 6307 16080 6316
rect 16028 6273 16046 6307
rect 16046 6273 16080 6307
rect 16028 6264 16080 6273
rect 11244 6196 11296 6248
rect 17040 6332 17092 6384
rect 17592 6264 17644 6316
rect 17868 6307 17920 6316
rect 17868 6273 17886 6307
rect 17886 6273 17920 6307
rect 17868 6264 17920 6273
rect 18052 6264 18104 6316
rect 20628 6332 20680 6384
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 18972 6264 19024 6316
rect 19984 6264 20036 6316
rect 19616 6239 19668 6248
rect 19616 6205 19625 6239
rect 19625 6205 19659 6239
rect 19659 6205 19668 6239
rect 19616 6196 19668 6205
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 3148 6060 3200 6112
rect 5356 6060 5408 6112
rect 6828 6128 6880 6180
rect 6736 6060 6788 6112
rect 8576 6103 8628 6112
rect 8576 6069 8585 6103
rect 8585 6069 8619 6103
rect 8619 6069 8628 6103
rect 8576 6060 8628 6069
rect 18604 6128 18656 6180
rect 10692 6060 10744 6112
rect 11060 6060 11112 6112
rect 11244 6060 11296 6112
rect 12256 6103 12308 6112
rect 12256 6069 12265 6103
rect 12265 6069 12299 6103
rect 12299 6069 12308 6103
rect 12256 6060 12308 6069
rect 12992 6060 13044 6112
rect 18972 6060 19024 6112
rect 19248 6060 19300 6112
rect 20720 6196 20772 6248
rect 19892 6060 19944 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 2504 5856 2556 5908
rect 4160 5856 4212 5908
rect 5540 5856 5592 5908
rect 20 5788 72 5840
rect 940 5788 992 5840
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 5080 5788 5132 5840
rect 5172 5788 5224 5840
rect 5632 5788 5684 5840
rect 8576 5856 8628 5908
rect 9128 5856 9180 5908
rect 9680 5856 9732 5908
rect 12532 5856 12584 5908
rect 13268 5856 13320 5908
rect 14280 5856 14332 5908
rect 17224 5856 17276 5908
rect 17408 5856 17460 5908
rect 19340 5856 19392 5908
rect 19524 5856 19576 5908
rect 2780 5763 2832 5772
rect 2780 5729 2789 5763
rect 2789 5729 2823 5763
rect 2823 5729 2832 5763
rect 2780 5720 2832 5729
rect 2964 5763 3016 5772
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 4804 5763 4856 5772
rect 2964 5720 3016 5729
rect 2688 5652 2740 5704
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 3424 5652 3476 5704
rect 2504 5584 2556 5636
rect 4344 5652 4396 5704
rect 4804 5729 4813 5763
rect 4813 5729 4847 5763
rect 4847 5729 4856 5763
rect 4804 5720 4856 5729
rect 15660 5788 15712 5840
rect 8208 5720 8260 5772
rect 8576 5720 8628 5772
rect 10508 5720 10560 5772
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 12808 5763 12860 5772
rect 12808 5729 12817 5763
rect 12817 5729 12851 5763
rect 12851 5729 12860 5763
rect 12808 5720 12860 5729
rect 14464 5763 14516 5772
rect 14464 5729 14473 5763
rect 14473 5729 14507 5763
rect 14507 5729 14516 5763
rect 14464 5720 14516 5729
rect 5448 5652 5500 5704
rect 5908 5695 5960 5704
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 6368 5695 6420 5704
rect 5908 5652 5960 5661
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 6644 5652 6696 5704
rect 6920 5652 6972 5704
rect 7196 5652 7248 5704
rect 7840 5652 7892 5704
rect 9036 5652 9088 5704
rect 5816 5584 5868 5636
rect 4068 5516 4120 5568
rect 5264 5516 5316 5568
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 6276 5516 6328 5568
rect 9864 5584 9916 5636
rect 10048 5584 10100 5636
rect 11060 5584 11112 5636
rect 11704 5584 11756 5636
rect 16856 5720 16908 5772
rect 19156 5788 19208 5840
rect 19800 5788 19852 5840
rect 17040 5763 17092 5772
rect 17040 5729 17049 5763
rect 17049 5729 17083 5763
rect 17083 5729 17092 5763
rect 17040 5720 17092 5729
rect 18144 5720 18196 5772
rect 20168 5856 20220 5908
rect 20352 5788 20404 5840
rect 20536 5720 20588 5772
rect 21272 5720 21324 5772
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 16948 5652 17000 5704
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 19892 5695 19944 5704
rect 18880 5652 18932 5661
rect 19892 5661 19901 5695
rect 19901 5661 19935 5695
rect 19935 5661 19944 5695
rect 19892 5652 19944 5661
rect 21548 5652 21600 5704
rect 11980 5516 12032 5568
rect 12716 5516 12768 5568
rect 13728 5559 13780 5568
rect 13728 5525 13737 5559
rect 13737 5525 13771 5559
rect 13771 5525 13780 5559
rect 13728 5516 13780 5525
rect 15568 5516 15620 5568
rect 15936 5516 15988 5568
rect 17868 5516 17920 5568
rect 17960 5516 18012 5568
rect 19248 5584 19300 5636
rect 19984 5584 20036 5636
rect 20904 5627 20956 5636
rect 20904 5593 20913 5627
rect 20913 5593 20947 5627
rect 20947 5593 20956 5627
rect 20904 5584 20956 5593
rect 19800 5559 19852 5568
rect 19800 5525 19809 5559
rect 19809 5525 19843 5559
rect 19843 5525 19852 5559
rect 19800 5516 19852 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 4988 5312 5040 5364
rect 8024 5312 8076 5364
rect 9036 5312 9088 5364
rect 9588 5312 9640 5364
rect 10968 5312 11020 5364
rect 940 5244 992 5296
rect 1676 5287 1728 5296
rect 1676 5253 1685 5287
rect 1685 5253 1719 5287
rect 1719 5253 1728 5287
rect 1676 5244 1728 5253
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 3424 5176 3476 5228
rect 4344 5244 4396 5296
rect 4436 5176 4488 5228
rect 2688 5151 2740 5160
rect 2688 5117 2697 5151
rect 2697 5117 2731 5151
rect 2731 5117 2740 5151
rect 2688 5108 2740 5117
rect 3240 5108 3292 5160
rect 5908 5176 5960 5228
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 9496 5176 9548 5228
rect 11796 5244 11848 5296
rect 12348 5244 12400 5296
rect 5816 5151 5868 5160
rect 848 5040 900 5092
rect 3332 5040 3384 5092
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 3884 5040 3936 5092
rect 112 4972 164 5024
rect 940 4972 992 5024
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 3792 4972 3844 5024
rect 3976 4972 4028 5024
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 4896 5040 4948 5092
rect 7656 5108 7708 5160
rect 8116 5151 8168 5160
rect 8116 5117 8125 5151
rect 8125 5117 8159 5151
rect 8159 5117 8168 5151
rect 8116 5108 8168 5117
rect 10508 5219 10560 5228
rect 10508 5185 10517 5219
rect 10517 5185 10551 5219
rect 10551 5185 10560 5219
rect 10508 5176 10560 5185
rect 12072 5176 12124 5228
rect 11796 5151 11848 5160
rect 11796 5117 11805 5151
rect 11805 5117 11839 5151
rect 11839 5117 11848 5151
rect 11796 5108 11848 5117
rect 14464 5312 14516 5364
rect 16304 5312 16356 5364
rect 17132 5312 17184 5364
rect 17408 5312 17460 5364
rect 17592 5355 17644 5364
rect 17592 5321 17601 5355
rect 17601 5321 17635 5355
rect 17635 5321 17644 5355
rect 17592 5312 17644 5321
rect 17960 5312 18012 5364
rect 19156 5312 19208 5364
rect 19340 5355 19392 5364
rect 19340 5321 19349 5355
rect 19349 5321 19383 5355
rect 19383 5321 19392 5355
rect 19340 5312 19392 5321
rect 19708 5312 19760 5364
rect 20536 5312 20588 5364
rect 16212 5244 16264 5296
rect 14924 5219 14976 5228
rect 14924 5185 14933 5219
rect 14933 5185 14967 5219
rect 14967 5185 14976 5219
rect 14924 5176 14976 5185
rect 5540 4972 5592 5024
rect 6920 4972 6972 5024
rect 8024 4972 8076 5024
rect 8668 5015 8720 5024
rect 8668 4981 8677 5015
rect 8677 4981 8711 5015
rect 8711 4981 8720 5015
rect 8668 4972 8720 4981
rect 9312 5040 9364 5092
rect 9496 5040 9548 5092
rect 12164 5083 12216 5092
rect 12164 5049 12173 5083
rect 12173 5049 12207 5083
rect 12207 5049 12216 5083
rect 12164 5040 12216 5049
rect 13636 5040 13688 5092
rect 14464 5083 14516 5092
rect 14464 5049 14473 5083
rect 14473 5049 14507 5083
rect 14507 5049 14516 5083
rect 14464 5040 14516 5049
rect 11060 4972 11112 5024
rect 14556 4972 14608 5024
rect 15752 5176 15804 5228
rect 16304 5176 16356 5228
rect 20168 5244 20220 5296
rect 20260 5244 20312 5296
rect 20628 5244 20680 5296
rect 17132 5219 17184 5228
rect 17132 5185 17141 5219
rect 17141 5185 17175 5219
rect 17175 5185 17184 5219
rect 17132 5176 17184 5185
rect 17316 5176 17368 5228
rect 17776 5176 17828 5228
rect 18144 5176 18196 5228
rect 19064 5219 19116 5228
rect 19064 5185 19073 5219
rect 19073 5185 19107 5219
rect 19107 5185 19116 5219
rect 19064 5176 19116 5185
rect 19892 5176 19944 5228
rect 19984 5176 20036 5228
rect 21364 5244 21416 5296
rect 19708 5108 19760 5160
rect 21088 5083 21140 5092
rect 21088 5049 21097 5083
rect 21097 5049 21131 5083
rect 21131 5049 21140 5083
rect 21088 5040 21140 5049
rect 15200 4972 15252 5024
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 15384 4972 15436 4981
rect 17960 4972 18012 5024
rect 18512 4972 18564 5024
rect 20076 4972 20128 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 2780 4768 2832 4820
rect 4896 4811 4948 4820
rect 1400 4632 1452 4684
rect 3792 4700 3844 4752
rect 4896 4777 4905 4811
rect 4905 4777 4939 4811
rect 4939 4777 4948 4811
rect 4896 4768 4948 4777
rect 5908 4811 5960 4820
rect 5908 4777 5917 4811
rect 5917 4777 5951 4811
rect 5951 4777 5960 4811
rect 5908 4768 5960 4777
rect 4988 4700 5040 4752
rect 2320 4632 2372 4684
rect 2688 4632 2740 4684
rect 4804 4632 4856 4684
rect 5540 4700 5592 4752
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 5448 4632 5500 4641
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 4344 4564 4396 4616
rect 4620 4564 4672 4616
rect 4712 4564 4764 4616
rect 7656 4768 7708 4820
rect 7748 4768 7800 4820
rect 8116 4768 8168 4820
rect 8484 4768 8536 4820
rect 9864 4768 9916 4820
rect 10508 4811 10560 4820
rect 10508 4777 10517 4811
rect 10517 4777 10551 4811
rect 10551 4777 10560 4811
rect 10508 4768 10560 4777
rect 10600 4768 10652 4820
rect 11244 4811 11296 4820
rect 11244 4777 11253 4811
rect 11253 4777 11287 4811
rect 11287 4777 11296 4811
rect 11244 4768 11296 4777
rect 12808 4768 12860 4820
rect 17132 4768 17184 4820
rect 6460 4632 6512 4684
rect 7380 4632 7432 4684
rect 8024 4632 8076 4684
rect 9128 4675 9180 4684
rect 7472 4564 7524 4616
rect 7748 4607 7800 4616
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 9128 4641 9137 4675
rect 9137 4641 9171 4675
rect 9171 4641 9180 4675
rect 9128 4632 9180 4641
rect 10968 4700 11020 4752
rect 10416 4632 10468 4684
rect 10600 4632 10652 4684
rect 2780 4539 2832 4548
rect 2780 4505 2789 4539
rect 2789 4505 2823 4539
rect 2823 4505 2832 4539
rect 2780 4496 2832 4505
rect 3424 4496 3476 4548
rect 3148 4428 3200 4480
rect 8116 4496 8168 4548
rect 11152 4564 11204 4616
rect 13268 4632 13320 4684
rect 17776 4700 17828 4752
rect 19616 4700 19668 4752
rect 19892 4700 19944 4752
rect 20168 4700 20220 4752
rect 11796 4564 11848 4616
rect 13176 4564 13228 4616
rect 13728 4564 13780 4616
rect 17132 4632 17184 4684
rect 20260 4632 20312 4684
rect 20812 4675 20864 4684
rect 20812 4641 20821 4675
rect 20821 4641 20855 4675
rect 20855 4641 20864 4675
rect 20812 4632 20864 4641
rect 14740 4564 14792 4616
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 16856 4564 16908 4616
rect 17224 4564 17276 4616
rect 18144 4564 18196 4616
rect 18788 4564 18840 4616
rect 19156 4564 19208 4616
rect 20076 4564 20128 4616
rect 15384 4496 15436 4548
rect 18880 4496 18932 4548
rect 19064 4496 19116 4548
rect 19708 4496 19760 4548
rect 3976 4428 4028 4480
rect 4620 4428 4672 4480
rect 5540 4471 5592 4480
rect 5540 4437 5549 4471
rect 5549 4437 5583 4471
rect 5583 4437 5592 4471
rect 5540 4428 5592 4437
rect 7564 4428 7616 4480
rect 8208 4471 8260 4480
rect 8208 4437 8217 4471
rect 8217 4437 8251 4471
rect 8251 4437 8260 4471
rect 8208 4428 8260 4437
rect 9128 4428 9180 4480
rect 13176 4428 13228 4480
rect 14924 4428 14976 4480
rect 15108 4428 15160 4480
rect 17224 4428 17276 4480
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 17684 4428 17736 4480
rect 19156 4428 19208 4480
rect 19524 4428 19576 4480
rect 20628 4471 20680 4480
rect 20628 4437 20637 4471
rect 20637 4437 20671 4471
rect 20671 4437 20680 4471
rect 20628 4428 20680 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 1676 4224 1728 4276
rect 3240 4224 3292 4276
rect 6000 4267 6052 4276
rect 6000 4233 6009 4267
rect 6009 4233 6043 4267
rect 6043 4233 6052 4267
rect 6000 4224 6052 4233
rect 7472 4224 7524 4276
rect 8116 4267 8168 4276
rect 8116 4233 8125 4267
rect 8125 4233 8159 4267
rect 8159 4233 8168 4267
rect 8116 4224 8168 4233
rect 7564 4156 7616 4208
rect 9772 4224 9824 4276
rect 10600 4224 10652 4276
rect 11060 4224 11112 4276
rect 15936 4224 15988 4276
rect 18880 4224 18932 4276
rect 19064 4224 19116 4276
rect 2320 4088 2372 4140
rect 2872 4131 2924 4140
rect 2872 4097 2881 4131
rect 2881 4097 2915 4131
rect 2915 4097 2924 4131
rect 2872 4088 2924 4097
rect 2688 4020 2740 4072
rect 3056 3952 3108 4004
rect 4620 4088 4672 4140
rect 5632 4088 5684 4140
rect 5724 4020 5776 4072
rect 5908 4088 5960 4140
rect 7472 4131 7524 4140
rect 7472 4097 7481 4131
rect 7481 4097 7515 4131
rect 7515 4097 7524 4131
rect 7472 4088 7524 4097
rect 7932 4131 7984 4140
rect 7932 4097 7941 4131
rect 7941 4097 7975 4131
rect 7975 4097 7984 4131
rect 7932 4088 7984 4097
rect 6000 4020 6052 4072
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 8668 4088 8720 4140
rect 10508 4156 10560 4208
rect 13544 4156 13596 4208
rect 15200 4156 15252 4208
rect 18604 4156 18656 4208
rect 20812 4199 20864 4208
rect 9588 4131 9640 4140
rect 9588 4097 9622 4131
rect 9622 4097 9640 4131
rect 9588 4088 9640 4097
rect 9864 4088 9916 4140
rect 12992 4088 13044 4140
rect 13268 4088 13320 4140
rect 14372 4088 14424 4140
rect 15476 4131 15528 4140
rect 15476 4097 15485 4131
rect 15485 4097 15519 4131
rect 15519 4097 15528 4131
rect 15476 4088 15528 4097
rect 15936 4131 15988 4140
rect 15936 4097 15945 4131
rect 15945 4097 15979 4131
rect 15979 4097 15988 4131
rect 15936 4088 15988 4097
rect 17040 4131 17092 4140
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 18696 4088 18748 4140
rect 18972 4088 19024 4140
rect 19432 4131 19484 4140
rect 19432 4097 19450 4131
rect 19450 4097 19484 4131
rect 20812 4165 20821 4199
rect 20821 4165 20855 4199
rect 20855 4165 20864 4199
rect 20812 4156 20864 4165
rect 19432 4088 19484 4097
rect 20444 4088 20496 4140
rect 2044 3884 2096 3936
rect 4068 3927 4120 3936
rect 4068 3893 4077 3927
rect 4077 3893 4111 3927
rect 4111 3893 4120 3927
rect 4068 3884 4120 3893
rect 5080 3927 5132 3936
rect 5080 3893 5089 3927
rect 5089 3893 5123 3927
rect 5123 3893 5132 3927
rect 5080 3884 5132 3893
rect 6092 3952 6144 4004
rect 9128 4020 9180 4072
rect 7564 3952 7616 4004
rect 8300 3952 8352 4004
rect 10416 3952 10468 4004
rect 15844 4020 15896 4072
rect 7656 3927 7708 3936
rect 7656 3893 7665 3927
rect 7665 3893 7699 3927
rect 7699 3893 7708 3927
rect 7656 3884 7708 3893
rect 10600 3884 10652 3936
rect 11612 3884 11664 3936
rect 14832 3952 14884 4004
rect 17500 4020 17552 4072
rect 20260 4020 20312 4072
rect 20536 4020 20588 4072
rect 18696 3952 18748 4004
rect 20444 3995 20496 4004
rect 20444 3961 20453 3995
rect 20453 3961 20487 3995
rect 20487 3961 20496 3995
rect 20444 3952 20496 3961
rect 12716 3884 12768 3936
rect 15200 3927 15252 3936
rect 15200 3893 15209 3927
rect 15209 3893 15243 3927
rect 15243 3893 15252 3927
rect 15200 3884 15252 3893
rect 16580 3884 16632 3936
rect 18236 3884 18288 3936
rect 18420 3884 18472 3936
rect 18788 3884 18840 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 2688 3723 2740 3732
rect 2688 3689 2697 3723
rect 2697 3689 2731 3723
rect 2731 3689 2740 3723
rect 2688 3680 2740 3689
rect 3056 3680 3108 3732
rect 4160 3680 4212 3732
rect 4252 3680 4304 3732
rect 5540 3680 5592 3732
rect 2872 3612 2924 3664
rect 4804 3612 4856 3664
rect 6736 3680 6788 3732
rect 7656 3680 7708 3732
rect 10416 3680 10468 3732
rect 10600 3680 10652 3732
rect 2136 3544 2188 3596
rect 3148 3587 3200 3596
rect 3148 3553 3157 3587
rect 3157 3553 3191 3587
rect 3191 3553 3200 3587
rect 3148 3544 3200 3553
rect 4160 3544 4212 3596
rect 4344 3587 4396 3596
rect 4344 3553 4353 3587
rect 4353 3553 4387 3587
rect 4387 3553 4396 3587
rect 4344 3544 4396 3553
rect 4988 3544 5040 3596
rect 5540 3544 5592 3596
rect 6276 3544 6328 3596
rect 8484 3612 8536 3664
rect 9404 3612 9456 3664
rect 12072 3655 12124 3664
rect 12072 3621 12081 3655
rect 12081 3621 12115 3655
rect 12115 3621 12124 3655
rect 12072 3612 12124 3621
rect 7472 3544 7524 3596
rect 5172 3476 5224 3528
rect 5356 3476 5408 3528
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 8208 3476 8260 3528
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 10508 3544 10560 3596
rect 12900 3680 12952 3732
rect 13176 3680 13228 3732
rect 15752 3680 15804 3732
rect 16120 3723 16172 3732
rect 16120 3689 16129 3723
rect 16129 3689 16163 3723
rect 16163 3689 16172 3723
rect 16120 3680 16172 3689
rect 16948 3680 17000 3732
rect 17040 3680 17092 3732
rect 18236 3680 18288 3732
rect 14648 3612 14700 3664
rect 17868 3612 17920 3664
rect 14372 3544 14424 3596
rect 14740 3587 14792 3596
rect 14740 3553 14749 3587
rect 14749 3553 14783 3587
rect 14783 3553 14792 3587
rect 14740 3544 14792 3553
rect 18144 3587 18196 3596
rect 18144 3553 18153 3587
rect 18153 3553 18187 3587
rect 18187 3553 18196 3587
rect 18144 3544 18196 3553
rect 10140 3519 10192 3528
rect 10140 3485 10158 3519
rect 10158 3485 10192 3519
rect 10140 3476 10192 3485
rect 2044 3451 2096 3460
rect 2044 3417 2053 3451
rect 2053 3417 2087 3451
rect 2087 3417 2096 3451
rect 2044 3408 2096 3417
rect 2964 3340 3016 3392
rect 3424 3340 3476 3392
rect 4620 3408 4672 3460
rect 7656 3408 7708 3460
rect 11980 3476 12032 3528
rect 12256 3476 12308 3528
rect 14280 3519 14332 3528
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 4528 3340 4580 3392
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 5632 3340 5684 3392
rect 6000 3340 6052 3392
rect 10692 3408 10744 3460
rect 11612 3408 11664 3460
rect 11796 3408 11848 3460
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 9036 3340 9088 3392
rect 9496 3340 9548 3392
rect 9680 3340 9732 3392
rect 11704 3340 11756 3392
rect 12348 3383 12400 3392
rect 12348 3349 12357 3383
rect 12357 3349 12391 3383
rect 12391 3349 12400 3383
rect 12348 3340 12400 3349
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 16580 3476 16632 3528
rect 14832 3408 14884 3460
rect 15108 3408 15160 3460
rect 14188 3340 14240 3392
rect 17316 3476 17368 3528
rect 17960 3476 18012 3528
rect 18788 3519 18840 3528
rect 18788 3485 18797 3519
rect 18797 3485 18831 3519
rect 18831 3485 18840 3519
rect 18788 3476 18840 3485
rect 19800 3680 19852 3732
rect 19064 3612 19116 3664
rect 20168 3544 20220 3596
rect 20904 3544 20956 3596
rect 19708 3476 19760 3528
rect 21548 3476 21600 3528
rect 18328 3408 18380 3460
rect 18420 3408 18472 3460
rect 19156 3408 19208 3460
rect 17868 3340 17920 3392
rect 18788 3340 18840 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 1860 3136 1912 3188
rect 4160 3136 4212 3188
rect 5816 3136 5868 3188
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 7656 3179 7708 3188
rect 7656 3145 7665 3179
rect 7665 3145 7699 3179
rect 7699 3145 7708 3179
rect 7656 3136 7708 3145
rect 1216 3068 1268 3120
rect 3976 3068 4028 3120
rect 5080 3068 5132 3120
rect 7472 3068 7524 3120
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2412 3000 2464 3052
rect 2596 3000 2648 3052
rect 3884 3000 3936 3052
rect 4068 3043 4120 3052
rect 4068 3009 4077 3043
rect 4077 3009 4111 3043
rect 4111 3009 4120 3043
rect 4068 3000 4120 3009
rect 4436 3000 4488 3052
rect 6092 3000 6144 3052
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 6460 3000 6512 3052
rect 6644 3000 6696 3052
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 11704 3136 11756 3188
rect 8576 3068 8628 3120
rect 13452 3068 13504 3120
rect 4528 2932 4580 2984
rect 5908 2864 5960 2916
rect 9312 3000 9364 3052
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 9680 3000 9732 3052
rect 9864 3043 9916 3052
rect 9864 3009 9873 3043
rect 9873 3009 9907 3043
rect 9907 3009 9916 3043
rect 9864 3000 9916 3009
rect 10784 3000 10836 3052
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 11980 3043 12032 3052
rect 9772 2975 9824 2984
rect 9772 2941 9781 2975
rect 9781 2941 9815 2975
rect 9815 2941 9824 2975
rect 9772 2932 9824 2941
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 12532 3000 12584 3052
rect 12716 3043 12768 3052
rect 12716 3009 12725 3043
rect 12725 3009 12759 3043
rect 12759 3009 12768 3043
rect 12716 3000 12768 3009
rect 17960 3136 18012 3188
rect 18696 3136 18748 3188
rect 19248 3136 19300 3188
rect 14648 3068 14700 3120
rect 14372 3000 14424 3052
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 17592 3068 17644 3120
rect 18972 3068 19024 3120
rect 17132 3000 17184 3052
rect 18880 3000 18932 3052
rect 19984 3043 20036 3052
rect 19984 3009 19993 3043
rect 19993 3009 20027 3043
rect 20027 3009 20036 3043
rect 19984 3000 20036 3009
rect 20628 3000 20680 3052
rect 20996 3000 21048 3052
rect 13084 2932 13136 2984
rect 13360 2975 13412 2984
rect 13360 2941 13369 2975
rect 13369 2941 13403 2975
rect 13403 2941 13412 2975
rect 13360 2932 13412 2941
rect 15568 2932 15620 2984
rect 16580 2932 16632 2984
rect 18236 2932 18288 2984
rect 20260 2975 20312 2984
rect 1124 2796 1176 2848
rect 2780 2796 2832 2848
rect 3424 2796 3476 2848
rect 4344 2796 4396 2848
rect 8024 2839 8076 2848
rect 8024 2805 8033 2839
rect 8033 2805 8067 2839
rect 8067 2805 8076 2839
rect 8024 2796 8076 2805
rect 8576 2796 8628 2848
rect 10324 2796 10376 2848
rect 11612 2839 11664 2848
rect 11612 2805 11621 2839
rect 11621 2805 11655 2839
rect 11655 2805 11664 2839
rect 11612 2796 11664 2805
rect 11704 2796 11756 2848
rect 18144 2864 18196 2916
rect 20260 2941 20269 2975
rect 20269 2941 20303 2975
rect 20303 2941 20312 2975
rect 20260 2932 20312 2941
rect 14188 2796 14240 2848
rect 14280 2796 14332 2848
rect 14740 2796 14792 2848
rect 15844 2796 15896 2848
rect 16304 2839 16356 2848
rect 16304 2805 16313 2839
rect 16313 2805 16347 2839
rect 16347 2805 16356 2839
rect 16304 2796 16356 2805
rect 16948 2796 17000 2848
rect 20076 2796 20128 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 1860 2635 1912 2644
rect 1860 2601 1869 2635
rect 1869 2601 1903 2635
rect 1903 2601 1912 2635
rect 1860 2592 1912 2601
rect 4528 2592 4580 2644
rect 5356 2592 5408 2644
rect 2964 2524 3016 2576
rect 3976 2524 4028 2576
rect 6460 2524 6512 2576
rect 7288 2592 7340 2644
rect 9864 2592 9916 2644
rect 12256 2635 12308 2644
rect 12256 2601 12265 2635
rect 12265 2601 12299 2635
rect 12299 2601 12308 2635
rect 12256 2592 12308 2601
rect 1216 2388 1268 2440
rect 3700 2456 3752 2508
rect 4160 2456 4212 2508
rect 5172 2456 5224 2508
rect 664 2320 716 2372
rect 2228 2363 2280 2372
rect 2228 2329 2237 2363
rect 2237 2329 2271 2363
rect 2271 2329 2280 2363
rect 2228 2320 2280 2329
rect 2780 2431 2832 2440
rect 2780 2397 2789 2431
rect 2789 2397 2823 2431
rect 2823 2397 2832 2431
rect 3240 2431 3292 2440
rect 2780 2388 2832 2397
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 6736 2456 6788 2508
rect 4804 2320 4856 2372
rect 6828 2388 6880 2440
rect 7012 2524 7064 2576
rect 7656 2499 7708 2508
rect 7656 2465 7665 2499
rect 7665 2465 7699 2499
rect 7699 2465 7708 2499
rect 7656 2456 7708 2465
rect 8024 2456 8076 2508
rect 7012 2388 7064 2440
rect 8208 2388 8260 2440
rect 3424 2295 3476 2304
rect 3424 2261 3433 2295
rect 3433 2261 3467 2295
rect 3467 2261 3476 2295
rect 3424 2252 3476 2261
rect 3976 2252 4028 2304
rect 7104 2252 7156 2304
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 9312 2388 9364 2440
rect 10140 2456 10192 2508
rect 10600 2499 10652 2508
rect 10600 2465 10609 2499
rect 10609 2465 10643 2499
rect 10643 2465 10652 2499
rect 10600 2456 10652 2465
rect 12440 2456 12492 2508
rect 14924 2592 14976 2644
rect 18880 2592 18932 2644
rect 20812 2592 20864 2644
rect 13636 2524 13688 2576
rect 15108 2524 15160 2576
rect 17132 2524 17184 2576
rect 18052 2524 18104 2576
rect 20904 2524 20956 2576
rect 10048 2388 10100 2440
rect 11612 2388 11664 2440
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13176 2388 13228 2397
rect 18880 2456 18932 2508
rect 15200 2431 15252 2440
rect 12256 2320 12308 2372
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16580 2388 16632 2440
rect 17224 2431 17276 2440
rect 17224 2397 17233 2431
rect 17233 2397 17267 2431
rect 17267 2397 17276 2431
rect 17224 2388 17276 2397
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 18512 2388 18564 2440
rect 20076 2431 20128 2440
rect 20076 2397 20085 2431
rect 20085 2397 20119 2431
rect 20119 2397 20128 2431
rect 20076 2388 20128 2397
rect 14372 2320 14424 2372
rect 11244 2252 11296 2304
rect 11980 2252 12032 2304
rect 12072 2252 12124 2304
rect 12440 2252 12492 2304
rect 12532 2252 12584 2304
rect 12900 2252 12952 2304
rect 13544 2252 13596 2304
rect 16212 2320 16264 2372
rect 15476 2252 15528 2304
rect 17684 2320 17736 2372
rect 17592 2252 17644 2304
rect 21180 2320 21232 2372
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 756 2048 808 2100
rect 4804 2048 4856 2100
rect 6828 2048 6880 2100
rect 9956 2048 10008 2100
rect 10968 2048 11020 2100
rect 12440 2048 12492 2100
rect 13452 2048 13504 2100
rect 13728 2048 13780 2100
rect 19248 2048 19300 2100
rect 3240 1980 3292 2032
rect 6276 1980 6328 2032
rect 7564 1980 7616 2032
rect 13176 1980 13228 2032
rect 3424 1912 3476 1964
rect 9496 1912 9548 1964
rect 8392 1844 8444 1896
rect 12072 1844 12124 1896
rect 3516 1776 3568 1828
rect 12256 1776 12308 1828
rect 4344 1708 4396 1760
rect 12624 1708 12676 1760
<< metal2 >>
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 2962 21312 3018 21321
rect 2962 21247 3018 21256
rect 1950 20904 2006 20913
rect 1950 20839 2006 20848
rect 1676 20460 1728 20466
rect 1676 20402 1728 20408
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1504 20097 1532 20198
rect 1490 20088 1546 20097
rect 1688 20058 1716 20402
rect 1490 20023 1546 20032
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1964 19990 1992 20839
rect 2044 20596 2096 20602
rect 2044 20538 2096 20544
rect 2056 20505 2084 20538
rect 2042 20496 2098 20505
rect 2976 20466 3004 21247
rect 5736 20602 5764 22200
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 12072 20528 12124 20534
rect 12072 20470 12124 20476
rect 2042 20431 2098 20440
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2964 20460 3016 20466
rect 2964 20402 3016 20408
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 2228 20256 2280 20262
rect 2228 20198 2280 20204
rect 1952 19984 2004 19990
rect 1952 19926 2004 19932
rect 2240 19854 2268 20198
rect 2608 20058 2636 20402
rect 5172 20392 5224 20398
rect 5172 20334 5224 20340
rect 4712 20324 4764 20330
rect 4712 20266 4764 20272
rect 3424 20256 3476 20262
rect 3424 20198 3476 20204
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 2686 19952 2742 19961
rect 2686 19887 2742 19896
rect 2700 19854 2728 19887
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2688 19848 2740 19854
rect 2688 19790 2740 19796
rect 1492 19712 1544 19718
rect 1490 19680 1492 19689
rect 1544 19680 1546 19689
rect 1490 19615 1546 19624
rect 1214 19544 1270 19553
rect 1214 19479 1270 19488
rect 938 18728 994 18737
rect 938 18663 994 18672
rect 20 17876 72 17882
rect 20 17818 72 17824
rect 32 5846 60 17818
rect 112 16516 164 16522
rect 112 16458 164 16464
rect 20 5840 72 5846
rect 20 5782 72 5788
rect 124 5030 152 16458
rect 848 15496 900 15502
rect 848 15438 900 15444
rect 664 7540 716 7546
rect 664 7482 716 7488
rect 112 5024 164 5030
rect 112 4966 164 4972
rect 676 2378 704 7482
rect 860 5098 888 15438
rect 952 7410 980 18663
rect 1030 18592 1086 18601
rect 1030 18527 1086 18536
rect 1044 17882 1072 18527
rect 1032 17876 1084 17882
rect 1032 17818 1084 17824
rect 1030 17776 1086 17785
rect 1030 17711 1086 17720
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 940 5840 992 5846
rect 938 5808 940 5817
rect 992 5808 994 5817
rect 938 5743 994 5752
rect 952 5302 980 5743
rect 940 5296 992 5302
rect 940 5238 992 5244
rect 848 5092 900 5098
rect 848 5034 900 5040
rect 940 5024 992 5030
rect 938 4992 940 5001
rect 992 4992 994 5001
rect 938 4927 994 4936
rect 1044 2774 1072 17711
rect 1122 17096 1178 17105
rect 1122 17031 1178 17040
rect 1136 7546 1164 17031
rect 1124 7540 1176 7546
rect 1124 7482 1176 7488
rect 1124 7404 1176 7410
rect 1124 7346 1176 7352
rect 1136 2854 1164 7346
rect 1228 3126 1256 19479
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 18873 1532 19110
rect 1688 18902 1716 19790
rect 2688 19440 2740 19446
rect 2688 19382 2740 19388
rect 3148 19440 3200 19446
rect 3148 19382 3200 19388
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 2504 19372 2556 19378
rect 2504 19314 2556 19320
rect 2042 19272 2098 19281
rect 2042 19207 2044 19216
rect 2096 19207 2098 19216
rect 2044 19178 2096 19184
rect 2240 18970 2268 19314
rect 2516 18970 2544 19314
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 1676 18896 1728 18902
rect 1490 18864 1546 18873
rect 1676 18838 1728 18844
rect 1490 18799 1546 18808
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1504 18465 1532 18566
rect 1490 18456 1546 18465
rect 1490 18391 1546 18400
rect 1306 18184 1362 18193
rect 1306 18119 1362 18128
rect 1216 3120 1268 3126
rect 1216 3062 1268 3068
rect 1124 2848 1176 2854
rect 1124 2790 1176 2796
rect 1320 2774 1348 18119
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1544 18048 1546 18057
rect 1490 17983 1546 17992
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17241 1532 17478
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 16833 1532 16934
rect 1490 16824 1546 16833
rect 1490 16759 1546 16768
rect 1584 16720 1636 16726
rect 1584 16662 1636 16668
rect 1398 16552 1454 16561
rect 1398 16487 1400 16496
rect 1452 16487 1454 16496
rect 1400 16458 1452 16464
rect 1492 16448 1544 16454
rect 1490 16416 1492 16425
rect 1544 16416 1546 16425
rect 1490 16351 1546 16360
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1400 15632 1452 15638
rect 1504 15609 1532 15846
rect 1400 15574 1452 15580
rect 1490 15600 1546 15609
rect 1412 13002 1440 15574
rect 1490 15535 1546 15544
rect 1492 15496 1544 15502
rect 1490 15464 1492 15473
rect 1544 15464 1546 15473
rect 1490 15399 1546 15408
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15201 1532 15302
rect 1490 15192 1546 15201
rect 1490 15127 1546 15136
rect 1492 14816 1544 14822
rect 1490 14784 1492 14793
rect 1544 14784 1546 14793
rect 1490 14719 1546 14728
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 13977 1532 14214
rect 1490 13968 1546 13977
rect 1490 13903 1546 13912
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1504 13569 1532 13670
rect 1490 13560 1546 13569
rect 1490 13495 1546 13504
rect 1492 13184 1544 13190
rect 1490 13152 1492 13161
rect 1544 13152 1546 13161
rect 1490 13087 1546 13096
rect 1412 12974 1532 13002
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1412 4690 1440 10746
rect 1504 8498 1532 12974
rect 1596 10674 1624 16662
rect 1688 16590 1716 18566
rect 2148 18426 2176 18702
rect 2136 18420 2188 18426
rect 2136 18362 2188 18368
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 1676 16584 1728 16590
rect 1872 16574 1900 17750
rect 1964 17338 1992 18226
rect 2700 18034 2728 19382
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3068 18766 3096 19110
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 2780 18692 2832 18698
rect 2780 18634 2832 18640
rect 2792 18426 2820 18634
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 3068 18290 3096 18566
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2700 18006 2820 18034
rect 2792 17882 2820 18006
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2228 17672 2280 17678
rect 2042 17640 2098 17649
rect 2228 17614 2280 17620
rect 2042 17575 2098 17584
rect 2056 17542 2084 17575
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 1676 16526 1728 16532
rect 1780 16546 1900 16574
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 12442 1716 15438
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1584 10192 1636 10198
rect 1584 10134 1636 10140
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1596 7342 1624 10134
rect 1688 7954 1716 11086
rect 1780 9042 1808 16546
rect 2136 16448 2188 16454
rect 2136 16390 2188 16396
rect 2042 16008 2098 16017
rect 2042 15943 2044 15952
rect 2096 15943 2098 15952
rect 2044 15914 2096 15920
rect 2148 15026 2176 16390
rect 2240 15706 2268 17614
rect 2318 17232 2374 17241
rect 2318 17167 2374 17176
rect 2504 17196 2556 17202
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2226 15600 2282 15609
rect 2226 15535 2282 15544
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2240 14906 2268 15535
rect 2148 14878 2268 14906
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 2042 14376 2098 14385
rect 1964 14074 1992 14350
rect 2042 14311 2098 14320
rect 2056 14278 2084 14311
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1872 11898 1900 12718
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 1964 11354 1992 12786
rect 1952 11348 2004 11354
rect 1952 11290 2004 11296
rect 2056 11200 2084 12786
rect 2148 12306 2176 14878
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2332 11830 2360 17167
rect 2504 17138 2556 17144
rect 2688 17196 2740 17202
rect 2688 17138 2740 17144
rect 2516 16250 2544 17138
rect 2700 16969 2728 17138
rect 2686 16960 2742 16969
rect 2686 16895 2742 16904
rect 2976 16454 3004 18226
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2608 16114 2636 16390
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2516 15706 2544 15982
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2792 15502 2820 15914
rect 2872 15904 2924 15910
rect 2872 15846 2924 15852
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2424 13462 2452 15030
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2412 13456 2464 13462
rect 2412 13398 2464 13404
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2240 11529 2268 11630
rect 2424 11626 2452 12242
rect 2412 11620 2464 11626
rect 2412 11562 2464 11568
rect 2226 11520 2282 11529
rect 2226 11455 2282 11464
rect 1872 11172 2084 11200
rect 1872 10146 1900 11172
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1964 10266 1992 10950
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1872 10118 1992 10146
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1490 6624 1546 6633
rect 1490 6559 1546 6568
rect 1504 6390 1532 6559
rect 1688 6390 1716 7890
rect 1872 7834 1900 9386
rect 1964 8265 1992 10118
rect 1950 8256 2006 8265
rect 1950 8191 2006 8200
rect 1780 7806 1900 7834
rect 1492 6384 1544 6390
rect 1676 6384 1728 6390
rect 1492 6326 1544 6332
rect 1582 6352 1638 6361
rect 1676 6326 1728 6332
rect 1582 6287 1638 6296
rect 1596 6118 1624 6287
rect 1780 6186 1808 7806
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 7546 1900 7686
rect 2056 7546 2084 11018
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2148 10130 2176 10406
rect 2424 10130 2452 11562
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2148 8634 2176 9522
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2240 8673 2268 8910
rect 2226 8664 2282 8673
rect 2136 8628 2188 8634
rect 2226 8599 2282 8608
rect 2136 8570 2188 8576
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2240 8265 2268 8366
rect 2226 8256 2282 8265
rect 2226 8191 2282 8200
rect 2332 8090 2360 9454
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2318 7984 2374 7993
rect 2424 7954 2452 8842
rect 2318 7919 2374 7928
rect 2412 7948 2464 7954
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1964 7002 1992 7346
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 2148 6882 2176 7686
rect 2332 7426 2360 7919
rect 2412 7890 2464 7896
rect 2332 7398 2452 7426
rect 2318 7304 2374 7313
rect 2318 7239 2374 7248
rect 1964 6854 2176 6882
rect 2332 6866 2360 7239
rect 2320 6860 2372 6866
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1596 3641 1624 6054
rect 1858 5808 1914 5817
rect 1858 5743 1860 5752
rect 1912 5743 1914 5752
rect 1860 5714 1912 5720
rect 1674 5672 1730 5681
rect 1674 5607 1730 5616
rect 1688 5302 1716 5607
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 1688 4282 1716 5238
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1582 3632 1638 3641
rect 1582 3567 1638 3576
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 768 2746 1072 2774
rect 1228 2746 1348 2774
rect 664 2372 716 2378
rect 664 2314 716 2320
rect 768 2106 796 2746
rect 1228 2446 1256 2746
rect 1872 2650 1900 3130
rect 1964 3058 1992 6854
rect 2320 6802 2372 6808
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2148 6458 2176 6598
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2148 6322 2176 6394
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2056 3466 2084 3878
rect 2148 3602 2176 4966
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 2228 4616 2280 4622
rect 2226 4584 2228 4593
rect 2280 4584 2282 4593
rect 2226 4519 2282 4528
rect 2332 4146 2360 4626
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2136 3596 2188 3602
rect 2136 3538 2188 3544
rect 2044 3460 2096 3466
rect 2044 3402 2096 3408
rect 2424 3058 2452 7398
rect 2516 5914 2544 13466
rect 2608 12986 2636 13874
rect 2700 13462 2728 14214
rect 2780 14000 2832 14006
rect 2780 13942 2832 13948
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2792 13274 2820 13942
rect 2700 13246 2820 13274
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2700 12186 2728 13246
rect 2780 13184 2832 13190
rect 2884 13172 2912 15846
rect 3160 14906 3188 19382
rect 3436 19378 3464 20198
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3792 19848 3844 19854
rect 3896 19836 3924 20198
rect 4172 19961 4200 20198
rect 4158 19952 4214 19961
rect 4158 19887 4214 19896
rect 4344 19916 4396 19922
rect 4344 19858 4396 19864
rect 3844 19825 3924 19836
rect 3844 19816 3938 19825
rect 3844 19808 3882 19816
rect 3792 19790 3844 19796
rect 3882 19751 3938 19760
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3252 17678 3280 18022
rect 3240 17672 3292 17678
rect 3238 17640 3240 17649
rect 3292 17640 3294 17649
rect 3238 17575 3294 17584
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3252 16590 3280 16934
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3252 16153 3280 16526
rect 3344 16250 3372 16526
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3238 16144 3294 16153
rect 3436 16130 3464 19314
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 4264 18630 4292 19314
rect 4356 19242 4384 19858
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4344 19236 4396 19242
rect 4344 19178 4396 19184
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 3976 18080 4028 18086
rect 3974 18048 3976 18057
rect 4028 18048 4030 18057
rect 3549 17980 3857 17989
rect 3974 17983 4030 17992
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3988 17746 4016 17983
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3896 16266 3924 17138
rect 3238 16079 3294 16088
rect 3344 16102 3464 16130
rect 3528 16238 3924 16266
rect 3344 15434 3372 16102
rect 3528 15994 3556 16238
rect 3884 16176 3936 16182
rect 3884 16118 3936 16124
rect 3700 16040 3752 16046
rect 3436 15966 3556 15994
rect 3698 16008 3700 16017
rect 3752 16008 3754 16017
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 3240 15360 3292 15366
rect 3238 15328 3240 15337
rect 3292 15328 3294 15337
rect 3238 15263 3294 15272
rect 3344 15162 3372 15370
rect 3436 15162 3464 15966
rect 3698 15943 3754 15952
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3332 15156 3384 15162
rect 3332 15098 3384 15104
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 2964 14884 3016 14890
rect 3160 14878 3280 14906
rect 2964 14826 3016 14832
rect 2832 13144 2912 13172
rect 2780 13126 2832 13132
rect 2792 12345 2820 13126
rect 2870 12880 2926 12889
rect 2870 12815 2926 12824
rect 2884 12782 2912 12815
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2872 12368 2924 12374
rect 2778 12336 2834 12345
rect 2872 12310 2924 12316
rect 2778 12271 2834 12280
rect 2700 12158 2820 12186
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 9466 2636 12038
rect 2792 10690 2820 12158
rect 2884 11937 2912 12310
rect 2976 12238 3004 14826
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 3068 13530 3096 13874
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 3068 12617 3096 12786
rect 3054 12608 3110 12617
rect 3054 12543 3110 12552
rect 3160 12306 3188 14758
rect 3252 12434 3280 14878
rect 3332 13728 3384 13734
rect 3332 13670 3384 13676
rect 3344 12889 3372 13670
rect 3436 13410 3464 15098
rect 3514 14920 3570 14929
rect 3514 14855 3516 14864
rect 3568 14855 3570 14864
rect 3516 14826 3568 14832
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3804 13954 3832 14350
rect 3896 14074 3924 16118
rect 3988 15502 4016 17478
rect 4080 17270 4108 17750
rect 4448 17542 4476 19790
rect 4528 19712 4580 19718
rect 4528 19654 4580 19660
rect 4540 18426 4568 19654
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4632 18358 4660 19450
rect 4724 18902 4752 20266
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 4712 18896 4764 18902
rect 4712 18838 4764 18844
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4068 17264 4120 17270
rect 4068 17206 4120 17212
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 4172 16658 4200 17070
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4080 14890 4108 16050
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 4080 14006 4108 14486
rect 4068 14000 4120 14006
rect 3804 13926 3924 13954
rect 4068 13942 4120 13948
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3436 13382 3556 13410
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3436 12986 3464 13262
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3330 12880 3386 12889
rect 3528 12850 3556 13382
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 3620 12986 3648 13194
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3804 12850 3832 13126
rect 3330 12815 3386 12824
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 3344 12646 3372 12718
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3252 12406 3372 12434
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 2964 12232 3016 12238
rect 3016 12192 3096 12220
rect 2964 12174 3016 12180
rect 2870 11928 2926 11937
rect 2870 11863 2926 11872
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2884 11218 2912 11630
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2700 10662 2820 10690
rect 2700 9738 2728 10662
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2792 10305 2820 10474
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2792 9897 2820 9930
rect 2884 9926 2912 11154
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2976 10606 3004 10950
rect 3068 10606 3096 12192
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3252 11830 3280 12038
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 3344 11354 3372 12406
rect 3896 11626 3924 13926
rect 4066 13696 4122 13705
rect 4066 13631 4122 13640
rect 4080 13274 4108 13631
rect 3988 13246 4108 13274
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3988 11354 4016 13246
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 4080 12850 4108 13126
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4080 12753 4108 12786
rect 4066 12744 4122 12753
rect 4066 12679 4122 12688
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11898 4108 12038
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4172 11354 4200 15302
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4264 14482 4292 14758
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4356 13530 4384 13874
rect 4344 13524 4396 13530
rect 4344 13466 4396 13472
rect 4344 12776 4396 12782
rect 4342 12744 4344 12753
rect 4396 12744 4398 12753
rect 4342 12679 4398 12688
rect 4448 12434 4476 17478
rect 4528 16992 4580 16998
rect 4526 16960 4528 16969
rect 4580 16960 4582 16969
rect 4526 16895 4582 16904
rect 4528 15360 4580 15366
rect 4724 15337 4752 18838
rect 5000 18766 5028 19110
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15570 4844 15846
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4528 15302 4580 15308
rect 4710 15328 4766 15337
rect 4540 14414 4568 15302
rect 4710 15263 4766 15272
rect 4816 14958 4844 15506
rect 4908 15042 4936 18566
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 5000 16590 5028 17070
rect 5092 16794 5120 18906
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5092 16454 5120 16730
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 5184 15910 5212 20334
rect 7012 20324 7064 20330
rect 7012 20266 7064 20272
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 19553 5304 20198
rect 6920 19848 6972 19854
rect 6826 19816 6882 19825
rect 6920 19790 6972 19796
rect 6826 19751 6882 19760
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 5262 19544 5318 19553
rect 5368 19514 5396 19654
rect 5262 19479 5318 19488
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5644 18766 5672 19246
rect 5632 18760 5684 18766
rect 5632 18702 5684 18708
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5368 17746 5396 18022
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16522 5304 16934
rect 5264 16516 5316 16522
rect 5264 16458 5316 16464
rect 5368 16250 5396 17682
rect 5460 17338 5488 17682
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5368 15570 5396 16186
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 5000 15162 5028 15302
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 4908 15014 5028 15042
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4526 13016 4582 13025
rect 4526 12951 4528 12960
rect 4580 12951 4582 12960
rect 4528 12922 4580 12928
rect 4540 12617 4568 12922
rect 4526 12608 4582 12617
rect 4526 12543 4582 12552
rect 4264 12406 4476 12434
rect 4528 12436 4580 12442
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 3332 11144 3384 11150
rect 3238 11112 3294 11121
rect 4264 11098 4292 12406
rect 4528 12378 4580 12384
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11665 4384 12038
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4342 11656 4398 11665
rect 4342 11591 4398 11600
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 3332 11086 3384 11092
rect 3238 11047 3294 11056
rect 3148 10736 3200 10742
rect 3148 10678 3200 10684
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 2872 9920 2924 9926
rect 2778 9888 2834 9897
rect 2872 9862 2924 9868
rect 2778 9823 2834 9832
rect 2700 9710 2912 9738
rect 2608 9438 2728 9466
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 7546 2636 9318
rect 2700 8362 2728 9438
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2504 5636 2556 5642
rect 2504 5578 2556 5584
rect 2516 4185 2544 5578
rect 2502 4176 2558 4185
rect 2502 4111 2558 4120
rect 2608 3058 2636 7210
rect 2700 7041 2728 7346
rect 2686 7032 2742 7041
rect 2686 6967 2688 6976
rect 2740 6967 2742 6976
rect 2688 6938 2740 6944
rect 2700 6907 2728 6938
rect 2792 6798 2820 9318
rect 2884 7886 2912 9710
rect 2976 9654 3004 10542
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 8022 3004 9318
rect 3068 9110 3096 10542
rect 3160 10062 3188 10678
rect 3252 10062 3280 11047
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 3160 9042 3188 9522
rect 3238 9480 3294 9489
rect 3238 9415 3294 9424
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3160 8430 3188 8842
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2884 7449 2912 7822
rect 2870 7440 2926 7449
rect 2870 7375 2926 7384
rect 2872 7336 2924 7342
rect 3160 7313 3188 8366
rect 3252 7886 3280 9415
rect 3344 8022 3372 11086
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 4080 11070 4292 11098
rect 3896 10742 3924 11018
rect 4080 10810 4108 11070
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3884 10736 3936 10742
rect 3882 10704 3884 10713
rect 3936 10704 3938 10713
rect 3882 10639 3938 10648
rect 3422 10568 3478 10577
rect 3422 10503 3478 10512
rect 3436 10266 3464 10503
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3514 10160 3570 10169
rect 3424 10124 3476 10130
rect 4172 10130 4200 10950
rect 4356 10130 4384 11154
rect 4448 11014 4476 11834
rect 4436 11008 4488 11014
rect 4436 10950 4488 10956
rect 3514 10095 3570 10104
rect 4160 10124 4212 10130
rect 3424 10066 3476 10072
rect 3332 8016 3384 8022
rect 3332 7958 3384 7964
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3330 7440 3386 7449
rect 3330 7375 3332 7384
rect 3384 7375 3386 7384
rect 3332 7346 3384 7352
rect 2872 7278 2924 7284
rect 3146 7304 3202 7313
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 5710 2728 6598
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2700 4690 2728 5102
rect 2792 4826 2820 5714
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2778 4584 2834 4593
rect 2778 4519 2780 4528
rect 2832 4519 2834 4528
rect 2780 4490 2832 4496
rect 2884 4298 2912 7278
rect 3146 7239 3202 7248
rect 3436 7206 3464 10066
rect 3528 9382 3556 10095
rect 4160 10066 4212 10072
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3700 9512 3752 9518
rect 3698 9480 3700 9489
rect 3752 9480 3754 9489
rect 3698 9415 3754 9424
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3896 9081 3924 9522
rect 3882 9072 3938 9081
rect 3882 9007 3938 9016
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3804 8362 3832 8842
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3896 8090 3924 9007
rect 3988 8634 4016 9998
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 4172 9722 4200 9862
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3988 7970 4016 8298
rect 3896 7942 4016 7970
rect 3896 7426 3924 7942
rect 3976 7880 4028 7886
rect 3974 7848 3976 7857
rect 4028 7848 4030 7857
rect 3974 7783 4030 7792
rect 3896 7398 4016 7426
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3436 6730 3464 7142
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3790 6760 3846 6769
rect 3424 6724 3476 6730
rect 3790 6695 3846 6704
rect 3424 6666 3476 6672
rect 3804 6662 3832 6695
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3160 6458 3188 6598
rect 3896 6458 3924 7278
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2976 5778 3004 6258
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3422 6216 3478 6225
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 3068 5710 3096 6190
rect 3422 6151 3478 6160
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3160 4842 3188 6054
rect 3436 5710 3464 6151
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3988 5794 4016 7398
rect 3804 5766 4016 5794
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3330 5264 3386 5273
rect 3330 5199 3332 5208
rect 3384 5199 3386 5208
rect 3424 5228 3476 5234
rect 3332 5170 3384 5176
rect 3424 5170 3476 5176
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 2792 4270 2912 4298
rect 2976 4814 3188 4842
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2700 3738 2728 4014
rect 2792 3777 2820 4270
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2778 3768 2834 3777
rect 2688 3732 2740 3738
rect 2778 3703 2834 3712
rect 2688 3674 2740 3680
rect 2884 3670 2912 4082
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2976 3482 3004 4814
rect 3054 4720 3110 4729
rect 3054 4655 3110 4664
rect 3068 4010 3096 4655
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 2884 3454 3004 3482
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2424 2961 2452 2994
rect 2410 2952 2466 2961
rect 2410 2887 2466 2896
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 2792 2446 2820 2790
rect 1216 2440 1268 2446
rect 2780 2440 2832 2446
rect 1216 2382 1268 2388
rect 2226 2408 2282 2417
rect 2226 2343 2228 2352
rect 2280 2343 2282 2352
rect 2608 2400 2780 2428
rect 2228 2314 2280 2320
rect 756 2100 808 2106
rect 756 2042 808 2048
rect 2240 800 2268 2314
rect 2608 800 2636 2400
rect 2780 2382 2832 2388
rect 2884 1737 2912 3454
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2976 2582 3004 3334
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 2870 1728 2926 1737
rect 2870 1663 2926 1672
rect 3068 1170 3096 3674
rect 3160 3602 3188 4422
rect 3252 4282 3280 5102
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3252 2038 3280 2382
rect 3240 2032 3292 2038
rect 3240 1974 3292 1980
rect 2976 1142 3096 1170
rect 2976 800 3004 1142
rect 3344 800 3372 5034
rect 3436 5001 3464 5170
rect 3804 5030 3832 5766
rect 3974 5672 4030 5681
rect 3974 5607 4030 5616
rect 3988 5386 4016 5607
rect 4080 5574 4108 9590
rect 4264 8922 4292 9862
rect 4448 9738 4476 10950
rect 4172 8894 4292 8922
rect 4356 9710 4476 9738
rect 4172 8537 4200 8894
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4158 8528 4214 8537
rect 4158 8463 4214 8472
rect 4172 8430 4200 8463
rect 4264 8430 4292 8774
rect 4160 8424 4212 8430
rect 4252 8424 4304 8430
rect 4160 8366 4212 8372
rect 4250 8392 4252 8401
rect 4304 8392 4306 8401
rect 4250 8327 4306 8336
rect 4356 7750 4384 9710
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4448 9217 4476 9522
rect 4540 9450 4568 12378
rect 4632 11914 4660 13874
rect 4724 12986 4752 14894
rect 4896 14408 4948 14414
rect 4894 14376 4896 14385
rect 4948 14376 4950 14385
rect 4804 14340 4856 14346
rect 4894 14311 4950 14320
rect 4804 14282 4856 14288
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4816 12866 4844 14282
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4724 12838 4844 12866
rect 4724 12050 4752 12838
rect 4802 12472 4858 12481
rect 4802 12407 4858 12416
rect 4816 12238 4844 12407
rect 4804 12232 4856 12238
rect 4802 12200 4804 12209
rect 4856 12200 4858 12209
rect 4802 12135 4858 12144
rect 4816 12109 4844 12135
rect 4724 12022 4844 12050
rect 4632 11886 4752 11914
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4632 11694 4660 11766
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4618 11520 4674 11529
rect 4618 11455 4674 11464
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4434 9208 4490 9217
rect 4434 9143 4490 9152
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4448 7410 4476 8978
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4172 5914 4200 6598
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4158 5536 4214 5545
rect 4158 5471 4214 5480
rect 3988 5358 4108 5386
rect 3884 5092 3936 5098
rect 3884 5034 3936 5040
rect 3792 5024 3844 5030
rect 3422 4992 3478 5001
rect 3792 4966 3844 4972
rect 3422 4927 3478 4936
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3424 4548 3476 4554
rect 3424 4490 3476 4496
rect 3436 3398 3464 4490
rect 3804 4321 3832 4694
rect 3790 4312 3846 4321
rect 3790 4247 3846 4256
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3896 3058 3924 5034
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3988 4486 4016 4966
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 4080 4026 4108 5358
rect 3988 3998 4108 4026
rect 3988 3369 4016 3998
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3974 3360 4030 3369
rect 3974 3295 4030 3304
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3436 2530 3464 2790
rect 3988 2774 4016 3062
rect 4080 3058 4108 3878
rect 4172 3738 4200 5471
rect 4264 3738 4292 6598
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4342 5944 4398 5953
rect 4342 5879 4398 5888
rect 4356 5710 4384 5879
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4356 4622 4384 5238
rect 4448 5234 4476 6258
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4356 3602 4384 4558
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4172 3505 4200 3538
rect 4158 3496 4214 3505
rect 4158 3431 4214 3440
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 3194 4200 3334
rect 4448 3210 4476 5170
rect 4540 3398 4568 9046
rect 4632 7886 4660 11455
rect 4724 8498 4752 11886
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4620 6724 4672 6730
rect 4620 6666 4672 6672
rect 4632 6254 4660 6666
rect 4816 6322 4844 12022
rect 4908 11082 4936 13126
rect 5000 12730 5028 15014
rect 5092 12850 5120 15506
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5000 12702 5120 12730
rect 4986 12472 5042 12481
rect 4986 12407 5042 12416
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4908 10266 4936 10542
rect 4896 10260 4948 10266
rect 4896 10202 4948 10208
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4908 9625 4936 9862
rect 4894 9616 4950 9625
rect 4894 9551 4950 9560
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 4908 8974 4936 9454
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4908 6730 4936 8910
rect 5000 7410 5028 12407
rect 5092 11898 5120 12702
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5092 11121 5120 11698
rect 5078 11112 5134 11121
rect 5078 11047 5134 11056
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5092 10713 5120 10950
rect 5078 10704 5134 10713
rect 5078 10639 5134 10648
rect 5184 10554 5212 14350
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5276 13326 5304 14214
rect 5368 13938 5396 15302
rect 5460 15094 5488 16934
rect 5552 16538 5580 18634
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5828 18170 5856 18566
rect 5632 18148 5684 18154
rect 5828 18142 5948 18170
rect 5632 18090 5684 18096
rect 5644 17338 5672 18090
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5816 18080 5868 18086
rect 5816 18022 5868 18028
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5552 16510 5672 16538
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5460 14278 5488 14894
rect 5552 14346 5580 16390
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5460 13841 5488 14010
rect 5446 13832 5502 13841
rect 5446 13767 5502 13776
rect 5644 13546 5672 16510
rect 5736 15314 5764 18022
rect 5828 17338 5856 18022
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 5920 15706 5948 18142
rect 6012 17785 6040 19654
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6748 19174 6776 19314
rect 6736 19168 6788 19174
rect 6736 19110 6788 19116
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 5998 17776 6054 17785
rect 5998 17711 6054 17720
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 6012 17134 6040 17614
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6000 17128 6052 17134
rect 6000 17070 6052 17076
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 5736 15286 5856 15314
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5552 13518 5672 13546
rect 5552 13433 5580 13518
rect 5632 13456 5684 13462
rect 5538 13424 5594 13433
rect 5632 13398 5684 13404
rect 5538 13359 5594 13368
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5460 12434 5488 12718
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5276 12406 5488 12434
rect 5276 11218 5304 12406
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11830 5396 12038
rect 5552 11830 5580 12650
rect 5356 11824 5408 11830
rect 5354 11792 5356 11801
rect 5540 11824 5592 11830
rect 5408 11792 5410 11801
rect 5540 11766 5592 11772
rect 5354 11727 5410 11736
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5276 10606 5304 11154
rect 5092 10526 5212 10554
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5092 9654 5120 10526
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5092 7546 5120 8774
rect 5184 7954 5212 10406
rect 5368 10198 5396 11727
rect 5448 11688 5500 11694
rect 5446 11656 5448 11665
rect 5500 11656 5502 11665
rect 5446 11591 5502 11600
rect 5644 11506 5672 13398
rect 5736 13394 5764 13874
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5736 12986 5764 13126
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5460 11478 5672 11506
rect 5460 10810 5488 11478
rect 5736 11370 5764 12786
rect 5828 11529 5856 15286
rect 6012 15094 6040 17070
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6564 16232 6592 18702
rect 6644 18624 6696 18630
rect 6644 18566 6696 18572
rect 6656 16697 6684 18566
rect 6642 16688 6698 16697
rect 6642 16623 6698 16632
rect 6748 16538 6776 19110
rect 6840 17882 6868 19751
rect 6932 19417 6960 19790
rect 7024 19718 7052 20266
rect 7378 19952 7434 19961
rect 7378 19887 7434 19896
rect 7012 19712 7064 19718
rect 7012 19654 7064 19660
rect 6918 19408 6974 19417
rect 6918 19343 6974 19352
rect 7024 18630 7052 19654
rect 7392 19417 7420 19887
rect 7484 19786 7512 20402
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 7472 19780 7524 19786
rect 7472 19722 7524 19728
rect 7378 19408 7434 19417
rect 7378 19343 7434 19352
rect 7288 18692 7340 18698
rect 7288 18634 7340 18640
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7024 18358 7052 18566
rect 7012 18352 7064 18358
rect 7010 18320 7012 18329
rect 7064 18320 7066 18329
rect 7010 18255 7066 18264
rect 7024 18229 7052 18255
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6840 17338 6868 17818
rect 7102 17640 7158 17649
rect 7102 17575 7158 17584
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 7024 17202 7052 17478
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 6918 16960 6974 16969
rect 6918 16895 6974 16904
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6380 16204 6592 16232
rect 6656 16510 6776 16538
rect 6380 15570 6408 16204
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 6000 14952 6052 14958
rect 6000 14894 6052 14900
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5920 14006 5948 14214
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 5814 11520 5870 11529
rect 5814 11455 5870 11464
rect 5736 11342 5856 11370
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5446 10296 5502 10305
rect 5446 10231 5502 10240
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 5460 10062 5488 10231
rect 5552 10198 5580 10610
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5644 10062 5672 10950
rect 5736 10130 5764 11222
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5276 7886 5304 9862
rect 5460 9586 5488 9998
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5368 9110 5396 9522
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5552 8974 5580 9318
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5262 7712 5318 7721
rect 5262 7647 5318 7656
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 5000 6458 5028 7346
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 4620 6248 4672 6254
rect 4620 6190 4672 6196
rect 4618 5944 4674 5953
rect 4618 5879 4674 5888
rect 4632 4622 4660 5879
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4622 4752 4966
rect 4816 4690 4844 5714
rect 5000 5370 5028 6258
rect 5092 5846 5120 6598
rect 5170 6216 5226 6225
rect 5170 6151 5172 6160
rect 5224 6151 5226 6160
rect 5172 6122 5224 6128
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4896 5092 4948 5098
rect 4896 5034 4948 5040
rect 4908 4826 4936 5034
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4988 4752 5040 4758
rect 4988 4694 5040 4700
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4620 4480 4672 4486
rect 4618 4448 4620 4457
rect 4672 4448 4674 4457
rect 4674 4406 4752 4434
rect 4618 4383 4674 4392
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4632 3913 4660 4082
rect 4618 3904 4674 3913
rect 4618 3839 4674 3848
rect 4618 3632 4674 3641
rect 4618 3567 4674 3576
rect 4632 3466 4660 3567
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4160 3188 4212 3194
rect 4448 3182 4568 3210
rect 4160 3130 4212 3136
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3988 2746 4108 2774
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3976 2576 4028 2582
rect 3974 2544 3976 2553
rect 4028 2544 4030 2553
rect 3436 2502 3556 2530
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3436 1970 3464 2246
rect 3424 1964 3476 1970
rect 3424 1906 3476 1912
rect 3528 1834 3556 2502
rect 3700 2508 3752 2514
rect 3974 2479 4030 2488
rect 4080 2496 4108 2746
rect 4160 2508 4212 2514
rect 3700 2450 3752 2456
rect 4080 2468 4160 2496
rect 3516 1828 3568 1834
rect 3516 1770 3568 1776
rect 3712 800 3740 2450
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3988 2145 4016 2246
rect 3974 2136 4030 2145
rect 3974 2071 4030 2080
rect 4080 800 4108 2468
rect 4160 2450 4212 2456
rect 4356 1766 4384 2790
rect 4448 2009 4476 2994
rect 4540 2990 4568 3182
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4724 2774 4752 4406
rect 4816 3670 4844 4626
rect 4894 3904 4950 3913
rect 4894 3839 4950 3848
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 4540 2746 4752 2774
rect 4540 2650 4568 2746
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4804 2372 4856 2378
rect 4804 2314 4856 2320
rect 4816 2106 4844 2314
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 4434 2000 4490 2009
rect 4434 1935 4490 1944
rect 4344 1760 4396 1766
rect 4344 1702 4396 1708
rect 4448 800 4476 1935
rect 4816 800 4844 2042
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 4908 762 4936 3839
rect 5000 3602 5028 4694
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5000 2961 5028 3538
rect 5092 3126 5120 3878
rect 5184 3534 5212 5782
rect 5276 5574 5304 7647
rect 5368 7546 5396 8502
rect 5644 8498 5672 9454
rect 5736 9178 5764 9590
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5722 9072 5778 9081
rect 5722 9007 5778 9016
rect 5736 8838 5764 9007
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5354 7032 5410 7041
rect 5354 6967 5410 6976
rect 5368 6934 5396 6967
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5368 6118 5396 6394
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5460 5710 5488 8434
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5552 5914 5580 8366
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5644 5846 5672 8434
rect 5736 7954 5764 8774
rect 5828 8401 5856 11342
rect 5920 10146 5948 13806
rect 6012 13734 6040 14894
rect 6090 14648 6146 14657
rect 6090 14583 6146 14592
rect 6104 14482 6132 14583
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 6012 13530 6040 13670
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 6000 13252 6052 13258
rect 6000 13194 6052 13200
rect 6012 12968 6040 13194
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6012 12940 6132 12968
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6012 12306 6040 12650
rect 6000 12300 6052 12306
rect 6000 12242 6052 12248
rect 6104 12084 6132 12940
rect 6012 12056 6132 12084
rect 6012 10810 6040 12056
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 5998 10704 6054 10713
rect 5998 10639 6000 10648
rect 6052 10639 6054 10648
rect 6000 10610 6052 10616
rect 5920 10118 6040 10146
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5814 8392 5870 8401
rect 5814 8327 5870 8336
rect 5920 8090 5948 9930
rect 6012 9704 6040 10118
rect 6288 9994 6316 10746
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6472 10146 6500 10678
rect 6564 10266 6592 15438
rect 6656 13569 6684 16510
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6748 15881 6776 15982
rect 6734 15872 6790 15881
rect 6734 15807 6790 15816
rect 6840 15201 6868 16662
rect 6932 16425 6960 16895
rect 6918 16416 6974 16425
rect 6918 16351 6974 16360
rect 7024 16182 7052 17138
rect 7116 16726 7144 17575
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7208 16794 7236 17070
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 7104 16720 7156 16726
rect 7104 16662 7156 16668
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7012 16176 7064 16182
rect 7012 16118 7064 16124
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 6826 15192 6882 15201
rect 6826 15127 6882 15136
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6826 14784 6882 14793
rect 6826 14719 6882 14728
rect 6642 13560 6698 13569
rect 6642 13495 6698 13504
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6656 12646 6684 13330
rect 6644 12640 6696 12646
rect 6642 12608 6644 12617
rect 6840 12617 6868 14719
rect 6696 12608 6698 12617
rect 6642 12543 6698 12552
rect 6826 12608 6882 12617
rect 6826 12543 6882 12552
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6736 11688 6788 11694
rect 6840 11665 6868 12378
rect 6932 11898 6960 14962
rect 7024 14958 7052 15506
rect 7116 15094 7144 15982
rect 7104 15088 7156 15094
rect 7104 15030 7156 15036
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7116 14521 7144 14554
rect 7102 14512 7158 14521
rect 7208 14482 7236 16390
rect 7102 14447 7158 14456
rect 7196 14476 7248 14482
rect 7116 14074 7144 14447
rect 7196 14418 7248 14424
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6736 11630 6788 11636
rect 6826 11656 6882 11665
rect 6644 10736 6696 10742
rect 6748 10724 6776 11630
rect 6826 11591 6882 11600
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6840 11354 6868 11494
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6696 10696 6776 10724
rect 6644 10678 6696 10684
rect 6642 10568 6698 10577
rect 6642 10503 6698 10512
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6472 10118 6592 10146
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6012 9676 6132 9704
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6012 9382 6040 9522
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6012 9081 6040 9318
rect 5998 9072 6054 9081
rect 5998 9007 6054 9016
rect 6104 8888 6132 9676
rect 6012 8860 6132 8888
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 6012 7970 6040 8860
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6564 8294 6592 10118
rect 6656 8634 6684 10503
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6656 8362 6684 8570
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5920 7942 6040 7970
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5722 6896 5778 6905
rect 5722 6831 5778 6840
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 4986 2952 5042 2961
rect 4986 2887 5042 2896
rect 5276 2774 5304 5510
rect 5460 4690 5488 5510
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5552 4758 5580 4966
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5552 3738 5580 4422
rect 5736 4298 5764 6831
rect 5828 6322 5856 7686
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5920 5710 5948 7942
rect 6000 7880 6052 7886
rect 6748 7857 6776 10202
rect 6840 10130 6868 11290
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6840 9586 6868 10066
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8537 6868 8978
rect 6826 8528 6882 8537
rect 6826 8463 6882 8472
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6000 7822 6052 7828
rect 6734 7848 6790 7857
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5816 5636 5868 5642
rect 5816 5578 5868 5584
rect 5828 5166 5856 5578
rect 5920 5545 5948 5646
rect 5906 5536 5962 5545
rect 5906 5471 5962 5480
rect 5908 5228 5960 5234
rect 5908 5170 5960 5176
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5920 4826 5948 5170
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5736 4270 5856 4298
rect 6012 4282 6040 7822
rect 6734 7783 6790 7792
rect 6840 7750 6868 8026
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6380 6798 6408 7142
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6564 6458 6592 7482
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6656 6798 6684 7278
rect 6748 6866 6776 7686
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6644 6792 6696 6798
rect 6696 6740 6776 6746
rect 6644 6734 6776 6740
rect 6656 6718 6776 6734
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 6366 6352 6422 6361
rect 6288 5574 6316 6326
rect 6366 6287 6422 6296
rect 6380 5710 6408 6287
rect 6368 5704 6420 5710
rect 6366 5672 6368 5681
rect 6420 5672 6422 5681
rect 6366 5607 6422 5616
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6458 4720 6514 4729
rect 6458 4655 6460 4664
rect 6512 4655 6514 4664
rect 6460 4626 6512 4632
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 5722 4176 5778 4185
rect 5632 4140 5684 4146
rect 5722 4111 5778 4120
rect 5632 4082 5684 4088
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5356 3528 5408 3534
rect 5552 3482 5580 3538
rect 5408 3476 5580 3482
rect 5356 3470 5580 3476
rect 5368 3454 5580 3470
rect 5644 3398 5672 4082
rect 5736 4078 5764 4111
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5184 2746 5304 2774
rect 5184 2514 5212 2746
rect 5368 2650 5396 3334
rect 5736 2774 5764 4014
rect 5828 3194 5856 4270
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6564 4162 6592 6394
rect 6748 6118 6776 6718
rect 6828 6180 6880 6186
rect 6828 6122 6880 6128
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6734 5672 6790 5681
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6288 4134 6592 4162
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5920 2922 5948 4082
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 6090 4040 6146 4049
rect 6012 3641 6040 4014
rect 6090 3975 6092 3984
rect 6144 3975 6146 3984
rect 6092 3946 6144 3952
rect 5998 3632 6054 3641
rect 6288 3602 6316 4134
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6458 3632 6514 3641
rect 5998 3567 6054 3576
rect 6276 3596 6328 3602
rect 6458 3567 6514 3576
rect 6276 3538 6328 3544
rect 6000 3392 6052 3398
rect 6472 3380 6500 3567
rect 6564 3534 6592 4014
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6656 3482 6684 5646
rect 6734 5607 6790 5616
rect 6748 3738 6776 5607
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6656 3454 6776 3482
rect 6472 3352 6592 3380
rect 6000 3334 6052 3340
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 6012 2774 6040 3334
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6090 3088 6146 3097
rect 6090 3023 6092 3032
rect 6144 3023 6146 3032
rect 6368 3052 6420 3058
rect 6092 2994 6144 3000
rect 6368 2994 6420 3000
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 5552 2746 5764 2774
rect 5920 2746 6040 2774
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5092 870 5212 898
rect 5092 762 5120 870
rect 5184 800 5212 870
rect 5552 800 5580 2746
rect 5920 800 5948 2746
rect 6380 2553 6408 2994
rect 6472 2582 6500 2994
rect 6564 2632 6592 3352
rect 6644 3052 6696 3058
rect 6748 3040 6776 3454
rect 6840 3058 6868 6122
rect 6932 5710 6960 11018
rect 7024 9178 7052 13330
rect 7116 13326 7144 14010
rect 7196 13932 7248 13938
rect 7196 13874 7248 13880
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7116 12306 7144 12582
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7208 12170 7236 13874
rect 7300 12782 7328 18634
rect 7392 17882 7420 19343
rect 7484 18630 7512 19722
rect 7576 19718 7604 20334
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 10324 20256 10376 20262
rect 10324 20198 10376 20204
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7576 19242 7604 19654
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7472 18624 7524 18630
rect 7472 18566 7524 18572
rect 7564 18284 7616 18290
rect 7564 18226 7616 18232
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7392 17678 7420 17818
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 16153 7420 17478
rect 7576 17338 7604 18226
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7378 16144 7434 16153
rect 7378 16079 7434 16088
rect 7484 15609 7512 17138
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7470 15600 7526 15609
rect 7576 15570 7604 15914
rect 7470 15535 7526 15544
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7576 15434 7604 15506
rect 7564 15428 7616 15434
rect 7564 15370 7616 15376
rect 7576 15042 7604 15370
rect 7392 15014 7604 15042
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7392 11914 7420 15014
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7484 14822 7512 14894
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7470 14648 7526 14657
rect 7470 14583 7472 14592
rect 7524 14583 7526 14592
rect 7472 14554 7524 14560
rect 7576 14362 7604 14894
rect 7484 14334 7604 14362
rect 7484 13870 7512 14334
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7472 13864 7524 13870
rect 7576 13841 7604 14214
rect 7472 13806 7524 13812
rect 7562 13832 7618 13841
rect 7208 11886 7420 11914
rect 7104 11008 7156 11014
rect 7102 10976 7104 10985
rect 7156 10976 7158 10985
rect 7102 10911 7158 10920
rect 7116 10470 7144 10911
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7116 10169 7144 10406
rect 7102 10160 7158 10169
rect 7102 10095 7158 10104
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 7208 8566 7236 11886
rect 7484 11694 7512 13806
rect 7562 13767 7618 13776
rect 7668 13326 7696 20198
rect 8312 19961 8340 20198
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8298 19952 8354 19961
rect 8298 19887 8354 19896
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8484 19848 8536 19854
rect 8484 19790 8536 19796
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 7944 19174 7972 19246
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7760 18290 7788 19110
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7760 13938 7788 16458
rect 7852 14006 7880 18770
rect 7944 17610 7972 19110
rect 8312 18816 8340 19790
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8220 18788 8340 18816
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 8220 18578 8248 18788
rect 8404 18766 8432 19246
rect 8392 18760 8444 18766
rect 8298 18728 8354 18737
rect 8392 18702 8444 18708
rect 8298 18663 8300 18672
rect 8352 18663 8354 18672
rect 8300 18634 8352 18640
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 7944 17338 7972 17546
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8036 17134 8064 18566
rect 8220 18550 8340 18578
rect 8208 18352 8260 18358
rect 8208 18294 8260 18300
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8128 17882 8156 18158
rect 8116 17876 8168 17882
rect 8116 17818 8168 17824
rect 8220 17542 8248 18294
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 7944 16726 7972 16757
rect 7932 16720 7984 16726
rect 7930 16688 7932 16697
rect 7984 16688 7986 16697
rect 7930 16623 7986 16632
rect 7944 16590 7972 16623
rect 7932 16584 7984 16590
rect 7932 16526 7984 16532
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7944 15366 7972 15846
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7944 15026 7972 15302
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7852 13258 7880 13942
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7668 12918 7696 13126
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7300 10266 7328 10678
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 8974 7328 9318
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7102 8392 7158 8401
rect 7300 8362 7328 8774
rect 7102 8327 7158 8336
rect 7288 8356 7340 8362
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 7024 7206 7052 7890
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7024 5953 7052 7142
rect 7116 6458 7144 8327
rect 7288 8298 7340 8304
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7010 5944 7066 5953
rect 7010 5879 7066 5888
rect 7208 5710 7236 7210
rect 7300 6866 7328 7890
rect 7392 7886 7420 11630
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7484 10742 7512 11086
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7470 10296 7526 10305
rect 7470 10231 7526 10240
rect 7484 10198 7512 10231
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7470 10024 7526 10033
rect 7470 9959 7472 9968
rect 7524 9959 7526 9968
rect 7472 9930 7524 9936
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7392 6730 7420 6938
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6696 3012 6776 3040
rect 6828 3052 6880 3058
rect 6644 2994 6696 3000
rect 6828 2994 6880 3000
rect 6932 2774 6960 4966
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6748 2746 6960 2774
rect 6564 2604 6684 2632
rect 6460 2576 6512 2582
rect 6366 2544 6422 2553
rect 6460 2518 6512 2524
rect 6366 2479 6422 2488
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6276 2032 6328 2038
rect 6276 1974 6328 1980
rect 6288 800 6316 1974
rect 6656 800 6684 2604
rect 6748 2514 6776 2746
rect 7024 2582 7052 3130
rect 7208 2774 7236 5646
rect 7116 2746 7236 2774
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 6840 2106 6868 2382
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 7024 800 7052 2382
rect 7116 2310 7144 2746
rect 7300 2650 7328 6258
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 4690 7420 6190
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7484 4622 7512 9318
rect 7576 9110 7604 12106
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7576 7002 7604 7754
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7562 6488 7618 6497
rect 7562 6423 7618 6432
rect 7576 6390 7604 6423
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7472 4616 7524 4622
rect 7392 4564 7472 4570
rect 7392 4558 7524 4564
rect 7392 4542 7512 4558
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7392 800 7420 4542
rect 7576 4486 7604 6190
rect 7668 5166 7696 12854
rect 7852 12850 7880 13194
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 8036 12730 8064 17070
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8116 16176 8168 16182
rect 8220 16153 8248 16390
rect 8206 16144 8262 16153
rect 8168 16124 8206 16130
rect 8116 16118 8206 16124
rect 8128 16102 8206 16118
rect 8206 16079 8262 16088
rect 8208 16040 8260 16046
rect 8312 16028 8340 18550
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8404 17746 8432 17818
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8260 16000 8340 16028
rect 8208 15982 8260 15988
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8220 15638 8248 15846
rect 8312 15638 8340 16000
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8128 14890 8156 15506
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8206 15056 8262 15065
rect 8206 14991 8262 15000
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 7760 12702 8064 12730
rect 7760 6905 7788 12702
rect 8128 12442 8156 14826
rect 8220 14822 8248 14991
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14113 8248 14758
rect 8206 14104 8262 14113
rect 8206 14039 8262 14048
rect 8206 13288 8262 13297
rect 8206 13223 8208 13232
rect 8260 13223 8262 13232
rect 8208 13194 8260 13200
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 7886 7880 11698
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7746 6896 7802 6905
rect 7746 6831 7802 6840
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7668 4826 7696 5102
rect 7760 4826 7788 6598
rect 7852 5710 7880 7414
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7564 4480 7616 4486
rect 7470 4448 7526 4457
rect 7564 4422 7616 4428
rect 7470 4383 7526 4392
rect 7484 4282 7512 4383
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7576 4214 7604 4422
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7484 4049 7512 4082
rect 7470 4040 7526 4049
rect 7470 3975 7526 3984
rect 7564 4004 7616 4010
rect 7564 3946 7616 3952
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7484 3126 7512 3538
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 7576 2038 7604 3946
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7668 3738 7696 3878
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7668 3194 7696 3402
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7654 2680 7710 2689
rect 7654 2615 7710 2624
rect 7668 2514 7696 2615
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7564 2032 7616 2038
rect 7564 1974 7616 1980
rect 7760 800 7788 4558
rect 7944 4146 7972 12038
rect 8128 11558 8156 12378
rect 8312 12374 8340 15438
rect 8300 12368 8352 12374
rect 8220 12328 8300 12356
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8220 11150 8248 12328
rect 8300 12310 8352 12316
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8312 10826 8340 11494
rect 8128 10798 8340 10826
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8036 10130 8064 10610
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8036 5370 8064 9114
rect 8128 6497 8156 10798
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8206 10568 8262 10577
rect 8206 10503 8262 10512
rect 8220 9994 8248 10503
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8312 9926 8340 10678
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8208 8560 8260 8566
rect 8206 8528 8208 8537
rect 8260 8528 8262 8537
rect 8206 8463 8262 8472
rect 8312 8430 8340 9454
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7313 8248 7686
rect 8206 7304 8262 7313
rect 8206 7239 8262 7248
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8114 6488 8170 6497
rect 8114 6423 8170 6432
rect 8116 6384 8168 6390
rect 8114 6352 8116 6361
rect 8168 6352 8170 6361
rect 8114 6287 8170 6296
rect 8220 5778 8248 6598
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8036 5030 8064 5306
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 8128 4826 8156 5102
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 8036 3584 8064 4626
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8128 4282 8156 4490
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8036 3556 8156 3584
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8036 2514 8064 2790
rect 8024 2508 8076 2514
rect 8024 2450 8076 2456
rect 8128 800 8156 3556
rect 8220 3534 8248 4422
rect 8312 4010 8340 7822
rect 8404 7410 8432 16390
rect 8496 15502 8524 19790
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8588 18426 8616 18566
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8588 18086 8616 18158
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8588 17134 8616 18022
rect 8680 17134 8708 18770
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8956 18222 8984 18566
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8484 14816 8536 14822
rect 8482 14784 8484 14793
rect 8536 14784 8538 14793
rect 8482 14719 8538 14728
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8588 14362 8616 17070
rect 8680 15706 8708 17070
rect 8772 16998 8800 17750
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8680 14498 8708 15642
rect 8758 15600 8814 15609
rect 8758 15535 8760 15544
rect 8812 15535 8814 15544
rect 8760 15506 8812 15512
rect 9034 15056 9090 15065
rect 9034 14991 9090 15000
rect 9048 14822 9076 14991
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 8680 14470 8892 14498
rect 8496 13734 8524 14350
rect 8588 14334 8708 14362
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 13394 8524 13670
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8496 11354 8524 13194
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10538 8524 10950
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8496 9500 8524 9998
rect 8588 9654 8616 14214
rect 8680 12646 8708 14334
rect 8864 14006 8892 14470
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 9140 13802 9168 18226
rect 9232 18193 9260 19110
rect 9218 18184 9274 18193
rect 9218 18119 9274 18128
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 9036 13320 9088 13326
rect 9088 13280 9168 13308
rect 9036 13262 9088 13268
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8666 12336 8722 12345
rect 8666 12271 8722 12280
rect 8680 10169 8708 12271
rect 9140 12238 9168 13280
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9048 11694 9076 12106
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 9140 11218 9168 12174
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9232 11150 9260 16594
rect 9324 16590 9352 19654
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9968 18970 9996 19382
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 9680 18896 9732 18902
rect 9678 18864 9680 18873
rect 9732 18864 9734 18873
rect 9678 18799 9734 18808
rect 9496 18760 9548 18766
rect 9496 18702 9548 18708
rect 9508 17202 9536 18702
rect 10060 18358 10088 19450
rect 10140 18420 10192 18426
rect 10140 18362 10192 18368
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 17338 9720 17478
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9496 17196 9548 17202
rect 9496 17138 9548 17144
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9416 16250 9444 16390
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9416 15337 9444 15846
rect 9402 15328 9458 15337
rect 9402 15263 9458 15272
rect 9508 14906 9536 16594
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9692 15178 9720 15438
rect 9600 15150 9720 15178
rect 9600 15026 9628 15150
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9324 14878 9536 14906
rect 9680 14884 9732 14890
rect 9324 14346 9352 14878
rect 9680 14826 9732 14832
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9324 13938 9352 14282
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9416 14074 9444 14214
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9312 13796 9364 13802
rect 9312 13738 9364 13744
rect 9324 13682 9352 13738
rect 9496 13728 9548 13734
rect 9324 13654 9444 13682
rect 9496 13670 9548 13676
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8666 10160 8722 10169
rect 8666 10095 8722 10104
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8496 9472 8616 9500
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8404 3534 8432 7210
rect 8496 5234 8524 9046
rect 8588 7970 8616 9472
rect 8680 8090 8708 10095
rect 9140 9654 9168 10406
rect 9232 10266 9260 11086
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9220 9648 9272 9654
rect 9220 9590 9272 9596
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9036 9104 9088 9110
rect 9036 9046 9088 9052
rect 8758 8664 8814 8673
rect 8758 8599 8760 8608
rect 8812 8599 8814 8608
rect 8760 8570 8812 8576
rect 9048 8514 9076 9046
rect 9140 8634 9168 9454
rect 9232 9178 9260 9590
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9048 8486 9168 8514
rect 9140 8294 9168 8486
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8588 7942 8708 7970
rect 8574 7576 8630 7585
rect 8574 7511 8630 7520
rect 8588 7342 8616 7511
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8680 6866 8708 7942
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8588 6322 8616 6802
rect 9140 6390 9168 8230
rect 9128 6384 9180 6390
rect 9128 6326 9180 6332
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 5914 8616 6054
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8496 3670 8524 4762
rect 8588 4457 8616 5714
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9048 5370 9076 5646
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8574 4448 8630 4457
rect 8574 4383 8630 4392
rect 8680 4146 8708 4966
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 9140 4690 9168 5850
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9128 4480 9180 4486
rect 9126 4448 9128 4457
rect 9180 4448 9182 4457
rect 9126 4383 9182 4392
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8576 3392 8628 3398
rect 8206 3360 8262 3369
rect 8576 3334 8628 3340
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 8206 3295 8262 3304
rect 8220 2446 8248 3295
rect 8588 3126 8616 3334
rect 8576 3120 8628 3126
rect 8482 3088 8538 3097
rect 8576 3062 8628 3068
rect 8482 3023 8538 3032
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8404 1902 8432 2246
rect 8392 1896 8444 1902
rect 8392 1838 8444 1844
rect 8496 800 8524 3023
rect 9048 2990 9076 3334
rect 9036 2984 9088 2990
rect 9034 2952 9036 2961
rect 9088 2952 9090 2961
rect 9034 2887 9090 2896
rect 8576 2848 8628 2854
rect 8574 2816 8576 2825
rect 8628 2816 8630 2825
rect 8574 2751 8630 2760
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 8850 2544 8906 2553
rect 8850 2479 8906 2488
rect 8864 800 8892 2479
rect 9140 1170 9168 4014
rect 9232 2774 9260 8774
rect 9324 8566 9352 12718
rect 9416 9382 9444 13654
rect 9508 12646 9536 13670
rect 9586 13424 9642 13433
rect 9586 13359 9642 13368
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9508 11121 9536 11494
rect 9494 11112 9550 11121
rect 9600 11082 9628 13359
rect 9494 11047 9550 11056
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9508 8838 9536 9658
rect 9600 9178 9628 11018
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9692 8906 9720 14826
rect 9784 14074 9812 18090
rect 9876 17066 9904 18158
rect 10152 17542 10180 18362
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10140 17536 10192 17542
rect 10138 17504 10140 17513
rect 10192 17504 10194 17513
rect 10138 17439 10194 17448
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9956 16720 10008 16726
rect 9954 16688 9956 16697
rect 10008 16688 10010 16697
rect 9954 16623 10010 16632
rect 10060 16114 10088 16730
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10060 15473 10088 15846
rect 10046 15464 10102 15473
rect 10046 15399 10102 15408
rect 10046 15192 10102 15201
rect 10046 15127 10102 15136
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 13190 9996 13330
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9784 11898 9812 12854
rect 10060 12434 10088 15127
rect 10152 14006 10180 17070
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10152 13530 10180 13942
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10244 12918 10272 17682
rect 10336 17338 10364 20198
rect 10796 19922 10824 20198
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 10796 19825 10824 19858
rect 10782 19816 10838 19825
rect 10782 19751 10838 19760
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10428 18970 10456 19246
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10428 17921 10456 18906
rect 10612 18834 10640 19450
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10414 17912 10470 17921
rect 10414 17847 10470 17856
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10322 16688 10378 16697
rect 10322 16623 10324 16632
rect 10376 16623 10378 16632
rect 10324 16594 10376 16600
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 9876 12406 10088 12434
rect 9876 12170 9904 12406
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9876 11626 9904 12106
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9876 11506 9904 11562
rect 9876 11478 9996 11506
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9494 8664 9550 8673
rect 9692 8622 9812 8650
rect 9692 8616 9720 8622
rect 9494 8599 9496 8608
rect 9548 8599 9550 8608
rect 9496 8570 9548 8576
rect 9646 8588 9720 8616
rect 9312 8560 9364 8566
rect 9646 8514 9674 8588
rect 9784 8566 9812 8622
rect 9312 8502 9364 8508
rect 9324 7546 9352 8502
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9508 8486 9674 8514
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9416 8362 9444 8434
rect 9508 8412 9536 8486
rect 9508 8401 9628 8412
rect 9494 8392 9628 8401
rect 9404 8356 9456 8362
rect 9550 8384 9628 8392
rect 9494 8327 9550 8336
rect 9404 8298 9456 8304
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9324 7177 9352 7278
rect 9310 7168 9366 7177
rect 9310 7103 9366 7112
rect 9416 6934 9444 7482
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9404 6928 9456 6934
rect 9508 6905 9536 7210
rect 9404 6870 9456 6876
rect 9494 6896 9550 6905
rect 9494 6831 9550 6840
rect 9600 6780 9628 8384
rect 9678 8256 9734 8265
rect 9678 8191 9734 8200
rect 9692 8090 9720 8191
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9772 8016 9824 8022
rect 9876 8004 9904 10610
rect 9824 7976 9904 8004
rect 9772 7958 9824 7964
rect 9968 7857 9996 11478
rect 10060 9994 10088 12038
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10140 10736 10192 10742
rect 10244 10690 10272 10950
rect 10192 10684 10272 10690
rect 10140 10678 10272 10684
rect 10152 10662 10272 10678
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 10060 8634 10088 9930
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10152 8265 10180 8842
rect 10138 8256 10194 8265
rect 10138 8191 10194 8200
rect 10048 7880 10100 7886
rect 9954 7848 10010 7857
rect 10048 7822 10100 7828
rect 9954 7783 10010 7792
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9508 6752 9628 6780
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9310 5944 9366 5953
rect 9310 5879 9366 5888
rect 9324 5098 9352 5879
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 9416 4978 9444 6326
rect 9508 5234 9536 6752
rect 9692 5914 9720 7686
rect 9968 7041 9996 7783
rect 9954 7032 10010 7041
rect 9954 6967 10010 6976
rect 10060 6848 10088 7822
rect 9968 6820 10088 6848
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9784 6458 9812 6734
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9876 5642 9904 6666
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9496 5092 9548 5098
rect 9496 5034 9548 5040
rect 9324 4950 9444 4978
rect 9324 4264 9352 4950
rect 9324 4236 9444 4264
rect 9310 4176 9366 4185
rect 9310 4111 9366 4120
rect 9324 3058 9352 4111
rect 9416 3670 9444 4236
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9508 3398 9536 5034
rect 9600 4146 9628 5306
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9692 3058 9720 3334
rect 9312 3052 9364 3058
rect 9680 3052 9732 3058
rect 9364 3012 9536 3040
rect 9312 2994 9364 3000
rect 9232 2746 9352 2774
rect 9324 2446 9352 2746
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9140 1142 9260 1170
rect 9232 800 9260 1142
rect 4908 734 5120 762
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9324 762 9352 2382
rect 9508 1970 9536 3012
rect 9680 2994 9732 3000
rect 9784 2990 9812 4218
rect 9876 4146 9904 4762
rect 9968 4321 9996 6820
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 9954 4312 10010 4321
rect 9954 4247 10010 4256
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9772 2984 9824 2990
rect 9772 2926 9824 2932
rect 9876 2650 9904 2994
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 10060 2446 10088 5578
rect 10152 3534 10180 6598
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10244 2774 10272 10662
rect 10336 10577 10364 15914
rect 10428 15434 10456 17682
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10428 14618 10456 15370
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10416 11348 10468 11354
rect 10416 11290 10468 11296
rect 10322 10568 10378 10577
rect 10322 10503 10378 10512
rect 10428 4690 10456 11290
rect 10520 6474 10548 17546
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10796 16833 10824 16934
rect 10782 16824 10838 16833
rect 10782 16759 10838 16768
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10612 14550 10640 16594
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10612 10742 10640 14010
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10612 8974 10640 9318
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10612 7410 10640 8910
rect 10704 7886 10732 16662
rect 10888 16250 10916 19994
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11256 19514 11284 19654
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10980 18057 11008 19110
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 10966 18048 11022 18057
rect 10966 17983 11022 17992
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11072 17746 11100 17818
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11164 16794 11192 18566
rect 11256 18426 11284 19246
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11244 18420 11296 18426
rect 11244 18362 11296 18368
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11520 17128 11572 17134
rect 11518 17096 11520 17105
rect 11716 17105 11744 19858
rect 11794 19408 11850 19417
rect 11794 19343 11796 19352
rect 11848 19343 11850 19352
rect 11796 19314 11848 19320
rect 11808 18737 11836 19314
rect 11900 19242 11928 19858
rect 12084 19854 12112 20470
rect 16132 20466 16160 20742
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 17236 20602 17264 22200
rect 17958 21312 18014 21321
rect 17958 21247 18014 21256
rect 17972 20806 18000 21247
rect 20626 20904 20682 20913
rect 20626 20839 20682 20848
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 19892 20528 19944 20534
rect 19892 20470 19944 20476
rect 20166 20496 20222 20505
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 11980 19712 12032 19718
rect 11980 19654 12032 19660
rect 11992 19417 12020 19654
rect 11978 19408 12034 19417
rect 11978 19343 12034 19352
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 12254 19272 12310 19281
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11794 18728 11850 18737
rect 11794 18663 11850 18672
rect 11796 18148 11848 18154
rect 11796 18090 11848 18096
rect 11572 17096 11574 17105
rect 11518 17031 11574 17040
rect 11702 17096 11758 17105
rect 11702 17031 11758 17040
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10888 15910 10916 16050
rect 10968 15972 11020 15978
rect 10968 15914 11020 15920
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10796 14618 10824 15030
rect 10888 14793 10916 15846
rect 10874 14784 10930 14793
rect 10874 14719 10930 14728
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10796 12986 10824 13262
rect 10784 12980 10836 12986
rect 10836 12940 10916 12968
rect 10784 12922 10836 12928
rect 10888 12442 10916 12940
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10888 11830 10916 12378
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10888 11694 10916 11766
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 11354 10916 11630
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10888 11218 10916 11290
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10782 10976 10838 10985
rect 10782 10911 10838 10920
rect 10796 10606 10824 10911
rect 10888 10810 10916 11154
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10888 10674 10916 10746
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10888 10266 10916 10610
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10888 9722 10916 10202
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10796 8294 10824 9590
rect 10888 9178 10916 9658
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10888 9042 10916 9114
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10980 8378 11008 15914
rect 11072 14521 11100 16594
rect 11702 16552 11758 16561
rect 11702 16487 11758 16496
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11164 15162 11192 15642
rect 11348 15609 11376 15642
rect 11334 15600 11390 15609
rect 11440 15570 11468 16118
rect 11716 15706 11744 16487
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11334 15535 11390 15544
rect 11428 15564 11480 15570
rect 11428 15506 11480 15512
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11256 15162 11284 15438
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11164 14890 11192 15098
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11058 14512 11114 14521
rect 11058 14447 11114 14456
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 11072 13870 11100 14282
rect 11164 14074 11192 14554
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12434 11100 13126
rect 11164 12782 11192 13194
rect 11256 12782 11284 14350
rect 11348 14346 11376 14758
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11716 13705 11744 15438
rect 11702 13696 11758 13705
rect 11702 13631 11758 13640
rect 11704 13456 11756 13462
rect 11704 13398 11756 13404
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11072 12406 11192 12434
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11072 10849 11100 12038
rect 11164 11257 11192 12406
rect 11150 11248 11206 11257
rect 11150 11183 11206 11192
rect 11256 11150 11284 12718
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11624 12170 11652 12378
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11058 10840 11114 10849
rect 11346 10843 11654 10852
rect 11058 10775 11114 10784
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11150 10704 11206 10713
rect 11072 9722 11100 10678
rect 11150 10639 11206 10648
rect 11060 9716 11112 9722
rect 11060 9658 11112 9664
rect 11164 9110 11192 10639
rect 11242 10296 11298 10305
rect 11242 10231 11298 10240
rect 11256 10062 11284 10231
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11716 9926 11744 13398
rect 11808 10062 11836 18090
rect 11900 14618 11928 19178
rect 11992 18630 12020 19246
rect 12254 19207 12256 19216
rect 12308 19207 12310 19216
rect 12256 19178 12308 19184
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11992 18193 12020 18362
rect 11978 18184 12034 18193
rect 11978 18119 12034 18128
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11992 15366 12020 17546
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 13462 11928 13670
rect 11888 13456 11940 13462
rect 11888 13398 11940 13404
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12442 11928 13126
rect 11992 12481 12020 15302
rect 12084 14346 12112 18022
rect 12452 17678 12480 19110
rect 12544 18970 12572 19314
rect 12636 18970 12664 19790
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12176 17338 12204 17478
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12176 15502 12204 16730
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12164 14816 12216 14822
rect 12162 14784 12164 14793
rect 12216 14784 12218 14793
rect 12162 14719 12218 14728
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 12084 14074 12112 14282
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12268 13818 12296 17614
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12360 16794 12388 17546
rect 12544 17066 12572 17750
rect 12728 17746 12756 20198
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 12900 19304 12952 19310
rect 12898 19272 12900 19281
rect 12952 19272 12954 19281
rect 12898 19207 12954 19216
rect 13372 19224 13400 19926
rect 13464 19514 13492 20334
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 14648 20324 14700 20330
rect 14648 20266 14700 20272
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 19854 13584 20198
rect 13832 19922 13860 20266
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 14660 19922 14688 20266
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13556 19310 13584 19790
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13452 19236 13504 19242
rect 13372 19196 13452 19224
rect 13452 19178 13504 19184
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12820 18698 12848 18770
rect 12898 18728 12954 18737
rect 12808 18692 12860 18698
rect 12898 18663 12954 18672
rect 12808 18634 12860 18640
rect 12820 18426 12848 18634
rect 12912 18630 12940 18663
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 18465 12940 18566
rect 12898 18456 12954 18465
rect 12808 18420 12860 18426
rect 12898 18391 12954 18400
rect 12808 18362 12860 18368
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12636 16250 12664 16458
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12360 15609 12388 15846
rect 12346 15600 12402 15609
rect 12346 15535 12402 15544
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12360 15162 12388 15370
rect 12440 15360 12492 15366
rect 12624 15360 12676 15366
rect 12440 15302 12492 15308
rect 12544 15320 12624 15348
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12360 14482 12388 15098
rect 12452 14521 12480 15302
rect 12438 14512 12494 14521
rect 12348 14476 12400 14482
rect 12438 14447 12494 14456
rect 12348 14418 12400 14424
rect 12360 14006 12388 14418
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12176 13790 12296 13818
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 11978 12472 12034 12481
rect 11888 12436 11940 12442
rect 11978 12407 12034 12416
rect 11888 12378 11940 12384
rect 12176 12374 12204 13790
rect 12360 12850 12388 13806
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12254 12336 12310 12345
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11152 9104 11204 9110
rect 11152 9046 11204 9052
rect 10888 8350 11008 8378
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10704 6866 10732 7278
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10520 6446 10640 6474
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10520 5234 10548 5714
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10520 4826 10548 5170
rect 10612 4826 10640 6446
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10520 4214 10548 4762
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10612 4282 10640 4626
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10428 3738 10456 3946
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10520 3602 10548 4150
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3738 10640 3878
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10704 3466 10732 6054
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10322 3088 10378 3097
rect 10796 3058 10824 7142
rect 10322 3023 10378 3032
rect 10784 3052 10836 3058
rect 10336 2854 10364 3023
rect 10784 2994 10836 3000
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10796 2774 10824 2994
rect 10152 2746 10272 2774
rect 10704 2746 10824 2774
rect 10888 2774 10916 8350
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 7886 11192 8230
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11164 7750 11192 7822
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11164 7342 11192 7686
rect 11152 7336 11204 7342
rect 11058 7304 11114 7313
rect 11152 7278 11204 7284
rect 11058 7239 11114 7248
rect 11072 6798 11100 7239
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10980 6644 11008 6734
rect 10980 6616 11100 6644
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 5778 11008 6258
rect 11072 6118 11100 6616
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10980 4758 11008 5306
rect 11072 5030 11100 5578
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 11072 4282 11100 4966
rect 11164 4622 11192 7142
rect 11256 6254 11284 9114
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11532 8974 11560 9046
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11716 6390 11744 9386
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11256 4826 11284 6054
rect 11716 5953 11744 6326
rect 11702 5944 11758 5953
rect 11702 5879 11758 5888
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 11072 3058 11100 3975
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11164 2774 11192 4558
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11624 3466 11652 3878
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 11716 3398 11744 5578
rect 11808 5302 11836 9658
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11796 5160 11848 5166
rect 11796 5102 11848 5108
rect 11808 4622 11836 5102
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11796 3460 11848 3466
rect 11796 3402 11848 3408
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11716 2854 11744 3130
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 10888 2746 11008 2774
rect 10152 2514 10180 2746
rect 10598 2680 10654 2689
rect 10598 2615 10654 2624
rect 10612 2514 10640 2615
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 9496 1964 9548 1970
rect 9496 1906 9548 1912
rect 9508 870 9628 898
rect 9508 762 9536 870
rect 9600 800 9628 870
rect 9968 800 9996 2042
rect 9324 734 9536 762
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10060 762 10088 2382
rect 10244 870 10364 898
rect 10244 762 10272 870
rect 10336 800 10364 870
rect 10704 800 10732 2746
rect 10980 2106 11008 2746
rect 11072 2746 11192 2774
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 11072 800 11100 2746
rect 11624 2446 11652 2790
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11256 1748 11284 2246
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11256 1720 11468 1748
rect 11440 800 11468 1720
rect 11808 800 11836 3402
rect 11900 2774 11928 11290
rect 11992 11121 12020 12038
rect 12084 11506 12112 12106
rect 12176 11830 12204 12310
rect 12254 12271 12310 12280
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 12084 11478 12204 11506
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11978 11112 12034 11121
rect 11978 11047 12034 11056
rect 12084 11014 12112 11290
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12070 10432 12126 10441
rect 12070 10367 12126 10376
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11992 8906 12020 9862
rect 12084 9450 12112 10367
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 12176 7546 12204 11478
rect 12268 9625 12296 12271
rect 12254 9616 12310 9625
rect 12360 9586 12388 12786
rect 12452 10849 12480 13126
rect 12438 10840 12494 10849
rect 12438 10775 12494 10784
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 9722 12480 10406
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12254 9551 12310 9560
rect 12348 9580 12400 9586
rect 12268 8634 12296 9551
rect 12348 9522 12400 9528
rect 12360 8906 12388 9522
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12256 8628 12308 8634
rect 12256 8570 12308 8576
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11992 6662 12020 7346
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12084 7002 12112 7142
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12360 6730 12388 7414
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12164 6724 12216 6730
rect 12164 6666 12216 6672
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11992 3534 12020 5510
rect 12084 5234 12112 6394
rect 12176 5817 12204 6666
rect 12256 6112 12308 6118
rect 12256 6054 12308 6060
rect 12162 5808 12218 5817
rect 12162 5743 12218 5752
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12084 3670 12112 5170
rect 12176 5098 12204 5743
rect 12164 5092 12216 5098
rect 12164 5034 12216 5040
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 12268 3534 12296 6054
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11992 2961 12020 2994
rect 11978 2952 12034 2961
rect 11978 2887 12034 2896
rect 12268 2774 12296 3470
rect 12360 3398 12388 5238
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 11900 2746 12020 2774
rect 11992 2310 12020 2746
rect 12176 2746 12296 2774
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 12084 1902 12112 2246
rect 12072 1896 12124 1902
rect 12072 1838 12124 1844
rect 12176 800 12204 2746
rect 12254 2680 12310 2689
rect 12254 2615 12256 2624
rect 12308 2615 12310 2624
rect 12256 2586 12308 2592
rect 12452 2514 12480 7142
rect 12544 6769 12572 15320
rect 12624 15302 12676 15308
rect 12728 15042 12756 17682
rect 12820 15450 12848 18362
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13082 16688 13138 16697
rect 13082 16623 13084 16632
rect 13136 16623 13138 16632
rect 13084 16594 13136 16600
rect 13188 16590 13216 18158
rect 13372 18057 13400 18158
rect 13358 18048 13414 18057
rect 13358 17983 13414 17992
rect 13266 17776 13322 17785
rect 13266 17711 13322 17720
rect 13280 17338 13308 17711
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13176 16176 13228 16182
rect 13176 16118 13228 16124
rect 12820 15422 13032 15450
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12636 15014 12756 15042
rect 12636 13326 12664 15014
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12728 13938 12756 14826
rect 12912 14414 12940 15302
rect 12900 14408 12952 14414
rect 12820 14368 12900 14396
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12636 12986 12664 13262
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12728 12434 12756 13126
rect 12636 12406 12756 12434
rect 12636 7426 12664 12406
rect 12714 10296 12770 10305
rect 12714 10231 12770 10240
rect 12728 7954 12756 10231
rect 12820 8906 12848 14368
rect 12900 14350 12952 14356
rect 12898 10024 12954 10033
rect 12898 9959 12954 9968
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12806 7984 12862 7993
rect 12716 7948 12768 7954
rect 12806 7919 12862 7928
rect 12716 7890 12768 7896
rect 12820 7886 12848 7919
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12636 7398 12756 7426
rect 12622 7304 12678 7313
rect 12622 7239 12624 7248
rect 12676 7239 12678 7248
rect 12624 7210 12676 7216
rect 12530 6760 12586 6769
rect 12530 6695 12586 6704
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12544 5914 12572 6598
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12728 5574 12756 7398
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12820 6662 12848 6802
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12820 6458 12848 6598
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12820 6322 12848 6394
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12820 5778 12848 6258
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12820 4826 12848 5714
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12530 3632 12586 3641
rect 12530 3567 12586 3576
rect 12544 3058 12572 3567
rect 12728 3058 12756 3878
rect 12912 3738 12940 9959
rect 13004 9382 13032 15422
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 11626 13124 13126
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13188 10538 13216 16118
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 15337 13400 15846
rect 13464 15502 13492 19178
rect 13556 18766 13584 19246
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13556 16726 13584 17478
rect 13648 17270 13676 18566
rect 13832 17338 13860 19654
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14188 18896 14240 18902
rect 14188 18838 14240 18844
rect 14200 18222 14228 18838
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 14292 17270 14320 19314
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14384 18329 14412 18566
rect 14370 18320 14426 18329
rect 14370 18255 14426 18264
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 13636 17264 13688 17270
rect 13636 17206 13688 17212
rect 14280 17264 14332 17270
rect 14384 17241 14412 17478
rect 14476 17338 14504 18226
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14568 17270 14596 17614
rect 14660 17542 14688 19858
rect 14740 18964 14792 18970
rect 14740 18906 14792 18912
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14556 17264 14608 17270
rect 14280 17206 14332 17212
rect 14370 17232 14426 17241
rect 14556 17206 14608 17212
rect 14370 17167 14426 17176
rect 14464 17196 14516 17202
rect 14384 17134 14412 17167
rect 14464 17138 14516 17144
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13358 15328 13414 15337
rect 13358 15263 13414 15272
rect 13464 15162 13492 15438
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13280 11626 13308 12174
rect 13360 12096 13412 12102
rect 13360 12038 13412 12044
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12990 7848 13046 7857
rect 12990 7783 13046 7792
rect 13004 6458 13032 7783
rect 13096 6662 13124 9522
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13004 4146 13032 6054
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 13096 2990 13124 6598
rect 13188 4622 13216 10474
rect 13280 9994 13308 11562
rect 13372 11257 13400 12038
rect 13358 11248 13414 11257
rect 13358 11183 13414 11192
rect 13464 10033 13492 12242
rect 13556 11801 13584 16662
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13648 12238 13676 16594
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13740 14278 13768 16526
rect 13832 15042 13860 17002
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 14476 16561 14504 17138
rect 14462 16552 14518 16561
rect 14384 16510 14462 16538
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 13832 15026 14044 15042
rect 14292 15026 14320 15370
rect 13832 15020 14056 15026
rect 13832 15014 14004 15020
rect 13832 14600 13860 15014
rect 14004 14962 14056 14968
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13912 14612 13964 14618
rect 13832 14572 13912 14600
rect 13912 14554 13964 14560
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14016 14006 14044 14214
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13832 13530 13860 13874
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13740 12617 13768 12650
rect 13726 12608 13782 12617
rect 13726 12543 13782 12552
rect 13832 12434 13860 12854
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13740 12406 13860 12434
rect 13740 12306 13768 12406
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13542 11792 13598 11801
rect 13542 11727 13598 11736
rect 13648 11694 13676 12174
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13832 11286 13860 12310
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13832 10266 13860 10678
rect 14292 10554 14320 12650
rect 14384 10810 14412 16510
rect 14462 16487 14518 16496
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14476 12345 14504 12378
rect 14462 12336 14518 12345
rect 14462 12271 14518 12280
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14568 10742 14596 15982
rect 14660 15910 14688 16390
rect 14648 15904 14700 15910
rect 14646 15872 14648 15881
rect 14700 15872 14702 15881
rect 14646 15807 14702 15816
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14660 12374 14688 12718
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14292 10526 14596 10554
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 13820 10056 13872 10062
rect 13450 10024 13506 10033
rect 13268 9988 13320 9994
rect 13820 9998 13872 10004
rect 13450 9959 13506 9968
rect 13268 9930 13320 9936
rect 13832 9926 13860 9998
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 9518 13860 9862
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 8906 13492 9318
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13280 5914 13308 8434
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 3738 13216 4422
rect 13280 4146 13308 4626
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13372 2990 13400 8570
rect 13464 7206 13492 8842
rect 13556 8430 13584 9386
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 14292 9110 14320 10202
rect 14372 10124 14424 10130
rect 14372 10066 14424 10072
rect 14280 9104 14332 9110
rect 14280 9046 14332 9052
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13648 7449 13676 7686
rect 13634 7440 13690 7449
rect 13556 7384 13634 7392
rect 13556 7364 13636 7384
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13556 4214 13584 7364
rect 13688 7375 13690 7384
rect 13636 7346 13688 7352
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 14292 6866 14320 7754
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13648 5098 13676 6598
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 14292 5914 14320 6326
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13740 4622 13768 5510
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 12268 1834 12296 2314
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 12452 2106 12480 2246
rect 12440 2100 12492 2106
rect 12440 2042 12492 2048
rect 12256 1828 12308 1834
rect 12256 1770 12308 1776
rect 12544 800 12572 2246
rect 12636 1766 12664 2382
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12912 800 12940 2246
rect 13188 2038 13216 2382
rect 13464 2106 13492 3062
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13452 2100 13504 2106
rect 13452 2042 13504 2048
rect 13176 2032 13228 2038
rect 13176 1974 13228 1980
rect 13280 870 13400 898
rect 13280 800 13308 870
rect 10060 734 10272 762
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13372 762 13400 870
rect 13556 762 13584 2246
rect 13648 800 13676 2518
rect 13740 2106 13768 4558
rect 14384 4146 14412 10066
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14476 7177 14504 9930
rect 14568 8974 14596 10526
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14660 8498 14688 11494
rect 14648 8492 14700 8498
rect 14568 8452 14648 8480
rect 14462 7168 14518 7177
rect 14462 7103 14518 7112
rect 14464 6996 14516 7002
rect 14464 6938 14516 6944
rect 14476 6322 14504 6938
rect 14568 6458 14596 8452
rect 14648 8434 14700 8440
rect 14752 7834 14780 18906
rect 14936 18850 14964 20198
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15212 19378 15240 19858
rect 15396 19854 15424 20334
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 14844 18834 14964 18850
rect 15396 18850 15424 19314
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15488 18970 15516 19246
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 14832 18828 14964 18834
rect 14884 18822 14964 18828
rect 15108 18828 15160 18834
rect 14832 18770 14884 18776
rect 15396 18822 15516 18850
rect 15108 18770 15160 18776
rect 15120 18290 15148 18770
rect 15290 18728 15346 18737
rect 15290 18663 15346 18672
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15014 17912 15070 17921
rect 15014 17847 15070 17856
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14844 16658 14872 17138
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14936 16522 14964 17478
rect 14924 16516 14976 16522
rect 14924 16458 14976 16464
rect 14936 16114 14964 16458
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14830 12880 14886 12889
rect 14830 12815 14886 12824
rect 14844 11558 14872 12815
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14936 11014 14964 11630
rect 15028 11121 15056 17847
rect 15120 15366 15148 18226
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15212 17270 15240 17478
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 15304 16794 15332 18663
rect 15382 17096 15438 17105
rect 15382 17031 15438 17040
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15304 16182 15332 16730
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15396 15366 15424 17031
rect 15488 16658 15516 18822
rect 15580 18222 15608 18906
rect 15764 18426 15792 19654
rect 15856 19514 15884 19654
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 16132 18850 16160 20402
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 16316 19922 16344 20334
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16040 18822 16160 18850
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15580 17338 15608 17478
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15488 15570 15516 16186
rect 15580 16114 15608 17002
rect 15672 16454 15700 18294
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15752 16992 15804 16998
rect 15752 16934 15804 16940
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15120 12753 15148 15098
rect 15292 13932 15344 13938
rect 15292 13874 15344 13880
rect 15304 13462 15332 13874
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15106 12744 15162 12753
rect 15106 12679 15162 12688
rect 15396 12238 15424 15302
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 15580 14414 15608 15030
rect 15764 14550 15792 16934
rect 15752 14544 15804 14550
rect 15752 14486 15804 14492
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15580 13870 15608 14350
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15580 13530 15608 13806
rect 15856 13530 15884 17682
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 15948 16250 15976 17138
rect 16040 16794 16068 18822
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16132 18290 16160 18634
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 16132 16130 16160 17750
rect 16224 17134 16252 19790
rect 16316 19394 16344 19858
rect 17236 19786 17264 20198
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17224 19780 17276 19786
rect 17224 19722 17276 19728
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 16408 19514 16436 19654
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16948 19440 17000 19446
rect 16946 19408 16948 19417
rect 17000 19408 17002 19417
rect 16316 19366 16436 19394
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16040 16102 16160 16130
rect 16040 14906 16068 16102
rect 16118 16008 16174 16017
rect 16118 15943 16174 15952
rect 16132 15065 16160 15943
rect 16118 15056 16174 15065
rect 16118 14991 16174 15000
rect 16040 14878 16160 14906
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15476 13388 15528 13394
rect 15476 13330 15528 13336
rect 15488 12986 15516 13330
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15580 12753 15608 13126
rect 15566 12744 15622 12753
rect 15566 12679 15622 12688
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15856 11830 15884 13466
rect 16040 12434 16068 14758
rect 16132 13938 16160 14878
rect 16224 14618 16252 17070
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16224 13326 16252 14554
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 15948 12406 16068 12434
rect 15948 12170 15976 12406
rect 15936 12164 15988 12170
rect 15936 12106 15988 12112
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 15014 11112 15070 11121
rect 15014 11047 15070 11056
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14936 10470 14964 10950
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14844 9926 14872 10202
rect 14936 10062 14964 10406
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14660 7806 14780 7834
rect 14660 7546 14688 7806
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14660 7002 14688 7346
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14832 6792 14884 6798
rect 14830 6760 14832 6769
rect 14884 6760 14886 6769
rect 14830 6695 14886 6704
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14476 5778 14504 6258
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14476 5370 14504 5714
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 14462 5264 14518 5273
rect 14462 5199 14518 5208
rect 14476 5098 14504 5199
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14278 4040 14334 4049
rect 14278 3975 14334 3984
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 14292 3534 14320 3975
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14200 2854 14228 3334
rect 14384 3058 14412 3538
rect 14372 3052 14424 3058
rect 14372 2994 14424 3000
rect 14568 2961 14596 4966
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14648 3664 14700 3670
rect 14648 3606 14700 3612
rect 14660 3126 14688 3606
rect 14752 3602 14780 4558
rect 14844 4010 14872 6598
rect 14936 5234 14964 7686
rect 15028 7313 15056 10678
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15856 9994 15884 10542
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15304 8566 15332 8842
rect 15200 8560 15252 8566
rect 15200 8502 15252 8508
rect 15292 8560 15344 8566
rect 15292 8502 15344 8508
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15014 7304 15070 7313
rect 15014 7239 15070 7248
rect 15120 6798 15148 7958
rect 15212 7041 15240 8502
rect 15198 7032 15254 7041
rect 15198 6967 15254 6976
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15028 6390 15056 6598
rect 15016 6384 15068 6390
rect 15304 6361 15332 8502
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15396 6730 15424 8298
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15016 6326 15068 6332
rect 15290 6352 15346 6361
rect 15290 6287 15346 6296
rect 15290 5944 15346 5953
rect 15290 5879 15346 5888
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14936 5001 14964 5170
rect 15200 5024 15252 5030
rect 14922 4992 14978 5001
rect 15200 4966 15252 4972
rect 14922 4927 14978 4936
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14830 3496 14886 3505
rect 14830 3431 14832 3440
rect 14884 3431 14886 3440
rect 14832 3402 14884 3408
rect 14648 3120 14700 3126
rect 14648 3062 14700 3068
rect 14554 2952 14610 2961
rect 14554 2887 14610 2896
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 13728 2100 13780 2106
rect 13728 2042 13780 2048
rect 14016 870 14136 898
rect 14016 800 14044 870
rect 13372 734 13584 762
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14108 762 14136 870
rect 14292 762 14320 2790
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14384 800 14412 2314
rect 14752 800 14780 2790
rect 14936 2650 14964 4422
rect 15120 3466 15148 4422
rect 15212 4214 15240 4966
rect 15304 4593 15332 5879
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15290 4584 15346 4593
rect 15396 4554 15424 4966
rect 15290 4519 15346 4528
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15200 4208 15252 4214
rect 15200 4150 15252 4156
rect 15488 4146 15516 9386
rect 15568 9376 15620 9382
rect 15566 9344 15568 9353
rect 15620 9344 15622 9353
rect 15566 9279 15622 9288
rect 15580 9042 15608 9279
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15580 6089 15608 6802
rect 15566 6080 15622 6089
rect 15566 6015 15622 6024
rect 15672 5846 15700 8910
rect 15856 7750 15884 9930
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15108 3460 15160 3466
rect 15108 3402 15160 3408
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15120 800 15148 2518
rect 15212 2446 15240 3878
rect 15580 2990 15608 5510
rect 15764 5234 15792 7346
rect 15856 6866 15884 7686
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15856 4078 15884 6802
rect 15948 5574 15976 12106
rect 16028 12096 16080 12102
rect 16028 12038 16080 12044
rect 16040 7750 16068 12038
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 9382 16252 11494
rect 16316 10606 16344 19110
rect 16408 18766 16436 19366
rect 16946 19343 17002 19352
rect 16948 18896 17000 18902
rect 16948 18838 17000 18844
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16408 17814 16436 18702
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16960 17649 16988 18838
rect 16946 17640 17002 17649
rect 17052 17610 17080 19654
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 16946 17575 17002 17584
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8634 16160 8774
rect 16316 8634 16344 9114
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 7818 16160 8230
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16132 6866 16160 7210
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 16040 4706 16068 6258
rect 16120 5704 16172 5710
rect 16118 5672 16120 5681
rect 16172 5672 16174 5681
rect 16118 5607 16174 5616
rect 16224 5302 16252 6598
rect 16316 5370 16344 6802
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16118 4720 16174 4729
rect 16040 4678 16118 4706
rect 16118 4655 16174 4664
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15948 4282 15976 4558
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15844 4072 15896 4078
rect 15948 4049 15976 4082
rect 15844 4014 15896 4020
rect 15934 4040 15990 4049
rect 15934 3975 15990 3984
rect 16132 3738 16160 4655
rect 16316 4593 16344 5170
rect 16302 4584 16358 4593
rect 16302 4519 16358 4528
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15764 2446 15792 3674
rect 16408 3534 16436 17478
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16960 14249 16988 15914
rect 17040 15564 17092 15570
rect 17040 15506 17092 15512
rect 17052 14346 17080 15506
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 16946 14240 17002 14249
rect 16544 14172 16852 14181
rect 16946 14175 17002 14184
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 17052 14090 17080 14282
rect 16960 14062 17080 14090
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16488 12640 16540 12646
rect 16486 12608 16488 12617
rect 16580 12640 16632 12646
rect 16540 12608 16542 12617
rect 16580 12582 16632 12588
rect 16486 12543 16542 12552
rect 16592 12442 16620 12582
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16960 12374 16988 14062
rect 17040 12912 17092 12918
rect 17040 12854 17092 12860
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 17052 12186 17080 12854
rect 16960 12158 17080 12186
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16592 11558 16620 11698
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16960 10198 16988 12158
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 11354 17080 12038
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17040 11008 17092 11014
rect 17040 10950 17092 10956
rect 17052 10742 17080 10950
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16946 10024 17002 10033
rect 16946 9959 17002 9968
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16960 8480 16988 9959
rect 17052 8906 17080 10678
rect 17144 10266 17172 19246
rect 17236 18766 17264 19722
rect 17512 19514 17540 19790
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17604 18766 17632 19654
rect 18248 19514 18276 20334
rect 18892 19854 18920 20334
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18052 19236 18104 19242
rect 18052 19178 18104 19184
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17236 17882 17264 18702
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17420 18154 17448 18226
rect 17408 18148 17460 18154
rect 17408 18090 17460 18096
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17236 17626 17264 17818
rect 17880 17678 17908 19110
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 17814 18000 18566
rect 17960 17808 18012 17814
rect 17960 17750 18012 17756
rect 17868 17672 17920 17678
rect 17236 17598 17356 17626
rect 17868 17614 17920 17620
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17236 16658 17264 17478
rect 17328 16794 17356 17598
rect 17592 17604 17644 17610
rect 17592 17546 17644 17552
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17236 15162 17264 16594
rect 17420 15638 17448 17002
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17512 16182 17540 16662
rect 17500 16176 17552 16182
rect 17500 16118 17552 16124
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 17512 15502 17540 15642
rect 17500 15496 17552 15502
rect 17314 15464 17370 15473
rect 17500 15438 17552 15444
rect 17314 15399 17370 15408
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17236 14414 17264 14962
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17328 14278 17356 15399
rect 17408 15360 17460 15366
rect 17408 15302 17460 15308
rect 17420 15026 17448 15302
rect 17408 15020 17460 15026
rect 17408 14962 17460 14968
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17236 12918 17264 14214
rect 17420 14074 17448 14350
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17328 12730 17356 13942
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17236 12702 17356 12730
rect 17236 12170 17264 12702
rect 17420 12646 17448 13262
rect 17512 12850 17540 15438
rect 17604 14414 17632 17546
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17696 17338 17724 17478
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17776 17332 17828 17338
rect 17776 17274 17828 17280
rect 17684 17196 17736 17202
rect 17684 17138 17736 17144
rect 17696 15706 17724 17138
rect 17788 16794 17816 17274
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17774 16688 17830 16697
rect 17774 16623 17776 16632
rect 17828 16623 17830 16632
rect 17776 16594 17828 16600
rect 17776 16516 17828 16522
rect 17776 16458 17828 16464
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17788 14822 17816 16458
rect 17868 15632 17920 15638
rect 17868 15574 17920 15580
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17682 14376 17738 14385
rect 17682 14311 17738 14320
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17408 12640 17460 12646
rect 17314 12608 17370 12617
rect 17408 12582 17460 12588
rect 17314 12543 17370 12552
rect 17328 12186 17356 12543
rect 17420 12442 17448 12582
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17224 12164 17276 12170
rect 17328 12158 17540 12186
rect 17224 12106 17276 12112
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17040 8900 17092 8906
rect 17040 8842 17092 8848
rect 16960 8452 17080 8480
rect 17052 8294 17080 8452
rect 17040 8288 17092 8294
rect 17040 8230 17092 8236
rect 17144 7886 17172 10202
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17236 9178 17264 10066
rect 17328 10010 17356 11834
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17420 10810 17448 11494
rect 17408 10804 17460 10810
rect 17408 10746 17460 10752
rect 17328 9982 17448 10010
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 17236 8566 17264 8842
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17040 7812 17092 7818
rect 17040 7754 17092 7760
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 17052 7410 17080 7754
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17052 7002 17080 7346
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 16578 6760 16634 6769
rect 16578 6695 16634 6704
rect 16592 6662 16620 6695
rect 16580 6656 16632 6662
rect 16948 6656 17000 6662
rect 16580 6598 16632 6604
rect 16946 6624 16948 6633
rect 17000 6624 17002 6633
rect 16544 6556 16852 6565
rect 16946 6559 17002 6568
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 17052 6390 17080 6938
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 16854 5808 16910 5817
rect 17052 5778 17080 6326
rect 16854 5743 16856 5752
rect 16908 5743 16910 5752
rect 17040 5772 17092 5778
rect 16856 5714 16908 5720
rect 17040 5714 17092 5720
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16960 4729 16988 5646
rect 17144 5370 17172 7346
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17236 6458 17264 7278
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17236 5914 17264 6394
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17328 5794 17356 9862
rect 17420 9217 17448 9982
rect 17512 9654 17540 12158
rect 17604 11937 17632 14214
rect 17590 11928 17646 11937
rect 17590 11863 17646 11872
rect 17604 11354 17632 11863
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17500 9512 17552 9518
rect 17500 9454 17552 9460
rect 17592 9512 17644 9518
rect 17592 9454 17644 9460
rect 17406 9208 17462 9217
rect 17406 9143 17462 9152
rect 17512 8634 17540 9454
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 17420 6866 17448 8502
rect 17604 6934 17632 9454
rect 17696 9450 17724 14311
rect 17788 12617 17816 14758
rect 17880 13802 17908 15574
rect 17972 14278 18000 16934
rect 18064 16250 18092 19178
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18524 18970 18552 19110
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18248 18290 18368 18306
rect 18248 18284 18380 18290
rect 18248 18278 18328 18284
rect 18248 17882 18276 18278
rect 18328 18226 18380 18232
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18144 17740 18196 17746
rect 18144 17682 18196 17688
rect 18156 17202 18184 17682
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18064 15858 18092 16186
rect 18142 16008 18198 16017
rect 18142 15943 18144 15952
rect 18196 15943 18198 15952
rect 18144 15914 18196 15920
rect 18064 15830 18276 15858
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 18064 14006 18092 15302
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 18156 13852 18184 14350
rect 18064 13824 18184 13852
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17774 12608 17830 12617
rect 17774 12543 17830 12552
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17776 11824 17828 11830
rect 17880 11812 17908 12106
rect 18064 11898 18092 13824
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18156 12442 18184 13466
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18142 12336 18198 12345
rect 18142 12271 18198 12280
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17828 11784 17908 11812
rect 17776 11766 17828 11772
rect 17880 11558 17908 11784
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17972 11286 18000 11698
rect 17960 11280 18012 11286
rect 18156 11234 18184 12271
rect 18248 11830 18276 15830
rect 18340 15026 18368 18090
rect 18432 18086 18460 18702
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 18432 17785 18460 17818
rect 18418 17776 18474 17785
rect 18418 17711 18474 17720
rect 18524 17678 18552 18906
rect 18616 17921 18644 19654
rect 19064 19508 19116 19514
rect 19064 19450 19116 19456
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18892 18970 18920 19314
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18696 18760 18748 18766
rect 18694 18728 18696 18737
rect 18748 18728 18750 18737
rect 18694 18663 18750 18672
rect 19076 18290 19104 19450
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19352 18834 19380 18906
rect 19536 18850 19564 20198
rect 19720 20058 19748 20402
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 19812 19990 19840 20402
rect 19800 19984 19852 19990
rect 19706 19952 19762 19961
rect 19800 19926 19852 19932
rect 19706 19887 19762 19896
rect 19616 19304 19668 19310
rect 19616 19246 19668 19252
rect 19628 19174 19656 19246
rect 19616 19168 19668 19174
rect 19616 19110 19668 19116
rect 19340 18828 19392 18834
rect 19536 18822 19656 18850
rect 19340 18770 19392 18776
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19536 18426 19564 18702
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18602 17912 18658 17921
rect 18602 17847 18658 17856
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18432 13530 18460 17138
rect 18616 16998 18644 17546
rect 19076 17338 19104 18226
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19536 17882 19564 18158
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19628 17746 19656 18822
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19720 17610 19748 19887
rect 19800 19848 19852 19854
rect 19800 19790 19852 19796
rect 19812 19514 19840 19790
rect 19800 19508 19852 19514
rect 19800 19450 19852 19456
rect 19904 17785 19932 20470
rect 20166 20431 20222 20440
rect 20180 20262 20208 20431
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20640 20058 20668 20839
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 20732 20097 20760 20198
rect 20718 20088 20774 20097
rect 20628 20052 20680 20058
rect 20718 20023 20774 20032
rect 20628 19994 20680 20000
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19996 19514 20024 19654
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 19890 17776 19946 17785
rect 19800 17740 19852 17746
rect 19890 17711 19946 17720
rect 19800 17682 19852 17688
rect 19812 17649 19840 17682
rect 19798 17640 19854 17649
rect 19708 17604 19760 17610
rect 19798 17575 19854 17584
rect 19708 17546 19760 17552
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 18696 17128 18748 17134
rect 18696 17070 18748 17076
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18524 16590 18552 16934
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18524 15978 18552 16390
rect 18512 15972 18564 15978
rect 18512 15914 18564 15920
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18236 11824 18288 11830
rect 18236 11766 18288 11772
rect 18248 11286 18276 11766
rect 17960 11222 18012 11228
rect 17972 11121 18000 11222
rect 18064 11206 18184 11234
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 17958 11112 18014 11121
rect 17958 11047 18014 11056
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17880 9586 17908 10202
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17684 9444 17736 9450
rect 17684 9386 17736 9392
rect 17696 8566 17724 9386
rect 17958 9344 18014 9353
rect 17958 9279 18014 9288
rect 17866 9208 17922 9217
rect 17866 9143 17922 9152
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17420 5914 17448 6802
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17236 5766 17356 5794
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 17144 4826 17172 5170
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 16946 4720 17002 4729
rect 16946 4655 17002 4664
rect 17132 4684 17184 4690
rect 17132 4626 17184 4632
rect 16856 4616 16908 4622
rect 16908 4564 16988 4570
rect 16856 4558 16988 4564
rect 16868 4542 16988 4558
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16592 3534 16620 3878
rect 16960 3738 16988 4542
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17052 3738 17080 4082
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 15934 3088 15990 3097
rect 17144 3058 17172 4626
rect 17236 4622 17264 5766
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 15934 3023 15936 3032
rect 15988 3023 15990 3032
rect 17132 3052 17184 3058
rect 15936 2994 15988 3000
rect 17132 2994 17184 3000
rect 16580 2984 16632 2990
rect 16302 2952 16358 2961
rect 16580 2926 16632 2932
rect 16302 2887 16358 2896
rect 16316 2854 16344 2887
rect 15844 2848 15896 2854
rect 15844 2790 15896 2796
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15488 800 15516 2246
rect 15856 800 15884 2790
rect 16592 2446 16620 2926
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16580 2440 16632 2446
rect 16580 2382 16632 2388
rect 16212 2372 16264 2378
rect 16212 2314 16264 2320
rect 16224 800 16252 2314
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16960 1170 16988 2790
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 16868 1142 16988 1170
rect 16592 870 16712 898
rect 16592 800 16620 870
rect 14108 734 14320 762
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16684 762 16712 870
rect 16868 762 16896 1142
rect 17144 898 17172 2518
rect 17236 2446 17264 4422
rect 17328 3534 17356 5170
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17420 2774 17448 5306
rect 17512 5250 17540 6666
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17604 6322 17632 6598
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17682 6216 17738 6225
rect 17682 6151 17738 6160
rect 17590 5400 17646 5409
rect 17590 5335 17592 5344
rect 17644 5335 17646 5344
rect 17592 5306 17644 5312
rect 17512 5222 17632 5250
rect 17498 4720 17554 4729
rect 17498 4655 17554 4664
rect 17512 4486 17540 4655
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17512 4078 17540 4422
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17604 3126 17632 5222
rect 17696 4486 17724 6151
rect 17788 5234 17816 9046
rect 17880 7818 17908 9143
rect 17972 8974 18000 9279
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17868 7812 17920 7818
rect 17868 7754 17920 7760
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 7274 18000 7686
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17880 7002 17908 7142
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17880 6322 17908 6938
rect 18064 6497 18092 11206
rect 18248 11098 18276 11222
rect 18156 11070 18276 11098
rect 18156 9926 18184 11070
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18248 10266 18276 10610
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18248 8820 18276 9522
rect 18340 8922 18368 13126
rect 18432 9058 18460 13194
rect 18708 12986 18736 17070
rect 18892 16794 18920 17138
rect 19616 17128 19668 17134
rect 19616 17070 19668 17076
rect 19708 17128 19760 17134
rect 19708 17070 19760 17076
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19628 16794 19656 17070
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 18878 16688 18934 16697
rect 18788 16652 18840 16658
rect 18878 16623 18934 16632
rect 18788 16594 18840 16600
rect 18800 13530 18828 16594
rect 18892 16114 18920 16623
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18892 14618 18920 14962
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18524 10266 18552 12922
rect 18800 12918 18828 13466
rect 18788 12912 18840 12918
rect 18788 12854 18840 12860
rect 18788 12776 18840 12782
rect 18786 12744 18788 12753
rect 18840 12744 18842 12753
rect 18786 12679 18842 12688
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 18602 12200 18658 12209
rect 18602 12135 18658 12144
rect 18616 10810 18644 12135
rect 18800 11354 18828 12242
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 18696 11144 18748 11150
rect 18694 11112 18696 11121
rect 18748 11112 18750 11121
rect 18694 11047 18750 11056
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18432 9030 18828 9058
rect 18340 8894 18644 8922
rect 18248 8792 18368 8820
rect 18340 8566 18368 8792
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 18248 6866 18276 8502
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18050 6488 18106 6497
rect 18050 6423 18106 6432
rect 18234 6488 18290 6497
rect 18234 6423 18290 6432
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 17958 6080 18014 6089
rect 17958 6015 18014 6024
rect 17972 5574 18000 6015
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 17420 2746 17540 2774
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17512 2009 17540 2746
rect 17788 2446 17816 4694
rect 17880 3670 17908 5510
rect 17972 5370 18000 5510
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 18064 5114 18092 6258
rect 18248 5930 18276 6423
rect 18156 5902 18276 5930
rect 18156 5778 18184 5902
rect 18340 5817 18368 7686
rect 18418 7440 18474 7449
rect 18418 7375 18474 7384
rect 18432 7342 18460 7375
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18510 7032 18566 7041
rect 18510 6967 18566 6976
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18326 5808 18382 5817
rect 18144 5772 18196 5778
rect 18326 5743 18382 5752
rect 18144 5714 18196 5720
rect 18142 5400 18198 5409
rect 18142 5335 18198 5344
rect 18156 5234 18184 5335
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 17972 5086 18092 5114
rect 17972 5030 18000 5086
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 18050 4992 18106 5001
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17972 3534 18000 4966
rect 18050 4927 18106 4936
rect 17960 3528 18012 3534
rect 18064 3505 18092 4927
rect 18156 4729 18184 5170
rect 18142 4720 18198 4729
rect 18142 4655 18198 4664
rect 18144 4616 18196 4622
rect 18144 4558 18196 4564
rect 18156 3602 18184 4558
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3738 18276 3878
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18340 3618 18368 5743
rect 18432 3942 18460 6802
rect 18524 6322 18552 6967
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18524 6225 18552 6258
rect 18510 6216 18566 6225
rect 18616 6186 18644 8894
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8566 18736 8774
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18708 8430 18736 8502
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18708 7886 18736 8026
rect 18800 8022 18828 9030
rect 18788 8016 18840 8022
rect 18788 7958 18840 7964
rect 18696 7880 18748 7886
rect 18694 7848 18696 7857
rect 18748 7848 18750 7857
rect 18694 7783 18750 7792
rect 18892 7478 18920 14214
rect 18984 11898 19012 15438
rect 19076 15094 19104 16390
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19064 15088 19116 15094
rect 19064 15030 19116 15036
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19076 13530 19104 14010
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 19444 12986 19472 13466
rect 19536 13258 19564 15982
rect 19628 15570 19656 16390
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19628 15065 19656 15302
rect 19614 15056 19670 15065
rect 19614 14991 19670 15000
rect 19616 13796 19668 13802
rect 19616 13738 19668 13744
rect 19628 13394 19656 13738
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19524 13252 19576 13258
rect 19524 13194 19576 13200
rect 19628 13002 19656 13330
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19536 12974 19656 13002
rect 19536 12714 19564 12974
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 18972 11892 19024 11898
rect 18972 11834 19024 11840
rect 19076 11642 19104 12378
rect 18984 11614 19104 11642
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 18984 7342 19012 11614
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11234 19104 11494
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19524 11280 19576 11286
rect 19076 11206 19196 11234
rect 19524 11222 19576 11228
rect 19168 11150 19196 11206
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 19156 11144 19208 11150
rect 19156 11086 19208 11092
rect 19168 10674 19196 11086
rect 19260 10674 19288 11154
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19168 10554 19196 10610
rect 19076 10526 19196 10554
rect 19076 10130 19104 10526
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 19062 9480 19118 9489
rect 19062 9415 19118 9424
rect 19076 8974 19104 9415
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 19076 8498 19104 8910
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19352 8566 19380 8842
rect 19536 8566 19564 11222
rect 19628 10742 19656 12854
rect 19616 10736 19668 10742
rect 19616 10678 19668 10684
rect 19720 10690 19748 17070
rect 19812 12442 19840 17138
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19904 15609 19932 15846
rect 19890 15600 19946 15609
rect 19890 15535 19946 15544
rect 19996 15502 20024 18566
rect 20088 18290 20116 18566
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20180 18193 20208 18226
rect 20166 18184 20222 18193
rect 20166 18119 20222 18128
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20166 16688 20222 16697
rect 20166 16623 20222 16632
rect 20180 16454 20208 16623
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19892 13864 19944 13870
rect 19944 13824 20024 13852
rect 19892 13806 19944 13812
rect 19890 13288 19946 13297
rect 19890 13223 19946 13232
rect 19904 13190 19932 13223
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19996 12850 20024 13824
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19798 11928 19854 11937
rect 19798 11863 19800 11872
rect 19852 11863 19854 11872
rect 19800 11834 19852 11840
rect 19720 10662 19840 10690
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19524 8560 19576 8566
rect 19524 8502 19576 8508
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 18788 7200 18840 7206
rect 18788 7142 18840 7148
rect 18970 7168 19026 7177
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18510 6151 18566 6160
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 18248 3590 18368 3618
rect 17960 3470 18012 3476
rect 18050 3496 18106 3505
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17880 3097 17908 3334
rect 17972 3194 18000 3470
rect 18050 3431 18106 3440
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 17866 3088 17922 3097
rect 17866 3023 17922 3032
rect 18156 2922 18184 3538
rect 18248 2990 18276 3590
rect 18328 3460 18380 3466
rect 18328 3402 18380 3408
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18236 2984 18288 2990
rect 18236 2926 18288 2932
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 18052 2576 18104 2582
rect 18052 2518 18104 2524
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17684 2372 17736 2378
rect 17684 2314 17736 2320
rect 17592 2304 17644 2310
rect 17592 2246 17644 2252
rect 17498 2000 17554 2009
rect 17498 1935 17554 1944
rect 16960 870 17172 898
rect 17328 870 17448 898
rect 16960 800 16988 870
rect 17328 800 17356 870
rect 16684 734 16896 762
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17420 762 17448 870
rect 17604 762 17632 2246
rect 17696 800 17724 2314
rect 18064 800 18092 2518
rect 18340 2446 18368 3402
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18432 800 18460 3402
rect 18524 2446 18552 4966
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 18616 2961 18644 4150
rect 18708 4146 18736 6598
rect 18800 4622 18828 7142
rect 18970 7103 19026 7112
rect 18984 6322 19012 7103
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18984 6202 19012 6258
rect 18892 6174 19012 6202
rect 18892 5817 18920 6174
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18878 5808 18934 5817
rect 18878 5743 18934 5752
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18892 5273 18920 5646
rect 18878 5264 18934 5273
rect 18878 5199 18934 5208
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18880 4548 18932 4554
rect 18880 4490 18932 4496
rect 18892 4282 18920 4490
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18984 4146 19012 6054
rect 19076 5234 19104 8230
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19536 7750 19564 7958
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19246 6760 19302 6769
rect 19302 6718 19380 6746
rect 19246 6695 19302 6704
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19260 6361 19288 6598
rect 19246 6352 19302 6361
rect 19246 6287 19302 6296
rect 19352 6202 19380 6718
rect 19260 6174 19380 6202
rect 19260 6118 19288 6174
rect 19248 6112 19300 6118
rect 19248 6054 19300 6060
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19536 5914 19564 7686
rect 19628 6730 19656 9522
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 19720 8294 19748 9454
rect 19812 9178 19840 10662
rect 19904 9450 19932 12174
rect 19996 11354 20024 12650
rect 20088 12442 20116 15506
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 20180 14793 20208 15302
rect 20166 14784 20222 14793
rect 20166 14719 20222 14728
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20076 12436 20128 12442
rect 20180 12434 20208 14350
rect 20272 13326 20300 18022
rect 20456 17898 20484 19858
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20812 19848 20864 19854
rect 21284 19825 21312 20198
rect 20812 19790 20864 19796
rect 21270 19816 21326 19825
rect 20548 18970 20576 19790
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20640 19281 20668 19450
rect 20824 19446 20852 19790
rect 21270 19751 21326 19760
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20626 19272 20682 19281
rect 20626 19207 20682 19216
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20456 17870 20576 17898
rect 20444 17740 20496 17746
rect 20444 17682 20496 17688
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20364 13462 20392 17478
rect 20456 14346 20484 17682
rect 20548 16561 20576 17870
rect 20640 17338 20668 18702
rect 20732 18222 20760 19314
rect 21284 18873 21312 19654
rect 21548 19236 21600 19242
rect 21548 19178 21600 19184
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21270 18864 21326 18873
rect 21270 18799 21326 18808
rect 21178 18728 21234 18737
rect 21178 18663 21234 18672
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20718 17640 20774 17649
rect 20718 17575 20774 17584
rect 20732 17542 20760 17575
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20732 16833 20760 16934
rect 20718 16824 20774 16833
rect 20718 16759 20774 16768
rect 20824 16590 20852 18226
rect 20902 16960 20958 16969
rect 20902 16895 20958 16904
rect 20916 16658 20944 16895
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20812 16584 20864 16590
rect 20534 16552 20590 16561
rect 20812 16526 20864 16532
rect 20534 16487 20590 16496
rect 20548 15586 20576 16487
rect 20628 16448 20680 16454
rect 20628 16390 20680 16396
rect 20640 16250 20668 16390
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20548 15558 20668 15586
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20456 14074 20484 14282
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20352 13456 20404 13462
rect 20352 13398 20404 13404
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20548 12986 20576 15438
rect 20640 15162 20668 15558
rect 21008 15502 21036 18362
rect 21088 18148 21140 18154
rect 21088 18090 21140 18096
rect 21100 17202 21128 18090
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21192 16776 21220 18663
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21284 18057 21312 18566
rect 21376 18329 21404 19110
rect 21362 18320 21418 18329
rect 21362 18255 21418 18264
rect 21364 18080 21416 18086
rect 21270 18048 21326 18057
rect 21364 18022 21416 18028
rect 21270 17983 21326 17992
rect 21376 17241 21404 18022
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21362 17232 21418 17241
rect 21362 17167 21418 17176
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21100 16748 21220 16776
rect 21100 16454 21128 16748
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20732 14385 20760 15302
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20812 14408 20864 14414
rect 20718 14376 20774 14385
rect 20916 14396 20944 14962
rect 20864 14368 20944 14396
rect 21088 14408 21140 14414
rect 20812 14350 20864 14356
rect 21088 14350 21140 14356
rect 20718 14311 20774 14320
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20824 13954 20852 14350
rect 20640 13394 20668 13942
rect 20824 13938 20944 13954
rect 20824 13932 20956 13938
rect 20824 13926 20904 13932
rect 20824 13530 20852 13926
rect 20904 13874 20956 13880
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20352 12436 20404 12442
rect 20180 12406 20300 12434
rect 20076 12378 20128 12384
rect 20272 12186 20300 12406
rect 20352 12378 20404 12384
rect 20088 12158 20300 12186
rect 19984 11348 20036 11354
rect 19984 11290 20036 11296
rect 19982 10160 20038 10169
rect 19982 10095 19984 10104
rect 20036 10095 20038 10104
rect 19984 10066 20036 10072
rect 20088 10062 20116 12158
rect 20168 12096 20220 12102
rect 20168 12038 20220 12044
rect 20180 11898 20208 12038
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 20166 10296 20222 10305
rect 20166 10231 20222 10240
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 20180 9994 20208 10231
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 19892 9444 19944 9450
rect 19892 9386 19944 9392
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19996 8650 20024 9318
rect 20180 9042 20208 9658
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 20272 8922 20300 11766
rect 19812 8622 20024 8650
rect 20088 8894 20300 8922
rect 19708 8288 19760 8294
rect 19708 8230 19760 8236
rect 19812 7154 19840 8622
rect 19892 8492 19944 8498
rect 19892 8434 19944 8440
rect 19720 7126 19840 7154
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19614 6352 19670 6361
rect 19614 6287 19670 6296
rect 19628 6254 19656 6287
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19156 5840 19208 5846
rect 19156 5782 19208 5788
rect 19168 5545 19196 5782
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19154 5536 19210 5545
rect 19154 5471 19210 5480
rect 19156 5364 19208 5370
rect 19260 5352 19288 5578
rect 19352 5370 19380 5850
rect 19720 5794 19748 7126
rect 19904 6984 19932 8434
rect 19812 6956 19932 6984
rect 19812 5846 19840 6956
rect 19982 6896 20038 6905
rect 19982 6831 20038 6840
rect 19996 6322 20024 6831
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 19892 6112 19944 6118
rect 19892 6054 19944 6060
rect 19444 5766 19748 5794
rect 19800 5840 19852 5846
rect 19800 5782 19852 5788
rect 19208 5324 19288 5352
rect 19340 5364 19392 5370
rect 19156 5306 19208 5312
rect 19340 5306 19392 5312
rect 19064 5228 19116 5234
rect 19064 5170 19116 5176
rect 19444 5114 19472 5766
rect 19904 5710 19932 6054
rect 19892 5704 19944 5710
rect 19614 5672 19670 5681
rect 19892 5646 19944 5652
rect 19614 5607 19670 5616
rect 19984 5636 20036 5642
rect 19444 5086 19564 5114
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19156 4616 19208 4622
rect 19536 4570 19564 5086
rect 19628 4758 19656 5607
rect 19984 5578 20036 5584
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19720 5166 19748 5306
rect 19708 5160 19760 5166
rect 19708 5102 19760 5108
rect 19616 4752 19668 4758
rect 19616 4694 19668 4700
rect 19156 4558 19208 4564
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 19076 4282 19104 4490
rect 19168 4486 19196 4558
rect 19444 4542 19564 4570
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 19444 4146 19472 4542
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 18708 3194 18736 3946
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18800 3534 18828 3878
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 19246 3632 19302 3641
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18602 2952 18658 2961
rect 18602 2887 18658 2896
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18800 800 18828 3334
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18892 2650 18920 2994
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 18892 2514 18920 2586
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 18984 1737 19012 3062
rect 18970 1728 19026 1737
rect 19076 1714 19104 3606
rect 19246 3567 19302 3576
rect 19156 3460 19208 3466
rect 19156 3402 19208 3408
rect 19168 3097 19196 3402
rect 19260 3194 19288 3567
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19154 3088 19210 3097
rect 19154 3023 19210 3032
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19246 2544 19302 2553
rect 19246 2479 19302 2488
rect 19260 2106 19288 2479
rect 19248 2100 19300 2106
rect 19248 2042 19300 2048
rect 19076 1686 19196 1714
rect 18970 1663 19026 1672
rect 19168 800 19196 1686
rect 19536 800 19564 4422
rect 19628 3777 19656 4694
rect 19708 4548 19760 4554
rect 19708 4490 19760 4496
rect 19614 3768 19670 3777
rect 19614 3703 19670 3712
rect 19720 3534 19748 4490
rect 19812 3738 19840 5510
rect 19996 5234 20024 5578
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19904 5001 19932 5170
rect 20088 5030 20116 8894
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20180 5914 20208 8774
rect 20272 7546 20300 8774
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20364 5846 20392 12378
rect 20548 12345 20576 12718
rect 20534 12336 20590 12345
rect 20444 12300 20496 12306
rect 20534 12271 20590 12280
rect 20444 12242 20496 12248
rect 20456 11694 20484 12242
rect 20640 11830 20668 13126
rect 20824 11898 20852 13126
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20916 11694 20944 13738
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21008 12442 21036 13466
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20456 9722 20484 11630
rect 20536 11620 20588 11626
rect 20536 11562 20588 11568
rect 20548 11082 20576 11562
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 20548 10810 20576 11018
rect 20536 10804 20588 10810
rect 20536 10746 20588 10752
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20548 10033 20576 10066
rect 20534 10024 20590 10033
rect 20534 9959 20590 9968
rect 20444 9716 20496 9722
rect 20444 9658 20496 9664
rect 20442 9616 20498 9625
rect 20442 9551 20498 9560
rect 20536 9580 20588 9586
rect 20456 8634 20484 9551
rect 20536 9522 20588 9528
rect 20548 9081 20576 9522
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20534 9072 20590 9081
rect 20534 9007 20590 9016
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20444 8628 20496 8634
rect 20444 8570 20496 8576
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20352 5840 20404 5846
rect 20352 5782 20404 5788
rect 20168 5296 20220 5302
rect 20168 5238 20220 5244
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20076 5024 20128 5030
rect 19890 4992 19946 5001
rect 20076 4966 20128 4972
rect 19890 4927 19946 4936
rect 19892 4752 19944 4758
rect 19892 4694 19944 4700
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19904 800 19932 4694
rect 20088 4622 20116 4966
rect 20180 4758 20208 5238
rect 20168 4752 20220 4758
rect 20168 4694 20220 4700
rect 20272 4690 20300 5238
rect 20260 4684 20312 4690
rect 20260 4626 20312 4632
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20272 4078 20300 4626
rect 20456 4146 20484 8230
rect 20548 7818 20576 8774
rect 20640 8430 20668 9318
rect 20732 8498 20760 11630
rect 21008 11218 21036 12378
rect 21100 12374 21128 14350
rect 21192 13410 21220 16594
rect 21284 16017 21312 16934
rect 21468 16561 21496 17478
rect 21454 16552 21510 16561
rect 21454 16487 21510 16496
rect 21454 16144 21510 16153
rect 21454 16079 21510 16088
rect 21270 16008 21326 16017
rect 21270 15943 21326 15952
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15026 21312 15846
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21284 13569 21312 14214
rect 21376 13977 21404 15302
rect 21362 13968 21418 13977
rect 21362 13903 21418 13912
rect 21270 13560 21326 13569
rect 21270 13495 21326 13504
rect 21192 13382 21312 13410
rect 21178 12880 21234 12889
rect 21178 12815 21234 12824
rect 21192 12442 21220 12815
rect 21180 12436 21232 12442
rect 21284 12434 21312 13382
rect 21284 12406 21404 12434
rect 21180 12378 21232 12384
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21284 11801 21312 12174
rect 21270 11792 21326 11801
rect 21270 11727 21326 11736
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 21270 11520 21326 11529
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 20824 8537 20852 9454
rect 20902 9208 20958 9217
rect 20902 9143 20958 9152
rect 20810 8528 20866 8537
rect 20720 8492 20772 8498
rect 20810 8463 20866 8472
rect 20720 8434 20772 8440
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 7886 20668 8230
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20534 7440 20590 7449
rect 20534 7375 20590 7384
rect 20548 7206 20576 7375
rect 20640 7342 20668 7822
rect 20732 7546 20760 8434
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 20628 7336 20680 7342
rect 20628 7278 20680 7284
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 20548 6730 20576 7142
rect 20640 6798 20668 7278
rect 20916 6866 20944 9143
rect 21086 8936 21142 8945
rect 21086 8871 21088 8880
rect 21140 8871 21142 8880
rect 21088 8842 21140 8848
rect 21088 8356 21140 8362
rect 21088 8298 21140 8304
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 20904 6860 20956 6866
rect 20904 6802 20956 6808
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20718 6760 20774 6769
rect 20536 6724 20588 6730
rect 20536 6666 20588 6672
rect 20640 6390 20668 6734
rect 20718 6695 20774 6704
rect 20628 6384 20680 6390
rect 20628 6326 20680 6332
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20548 5370 20576 5714
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20548 4078 20576 5306
rect 20640 5302 20668 6326
rect 20732 6254 20760 6695
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20810 6352 20866 6361
rect 20810 6287 20866 6296
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20628 5296 20680 5302
rect 20628 5238 20680 5244
rect 20824 4690 20852 6287
rect 20916 5642 20944 6394
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20812 4684 20864 4690
rect 20864 4644 20944 4672
rect 20812 4626 20864 4632
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 20640 4185 20668 4422
rect 20812 4208 20864 4214
rect 20626 4176 20682 4185
rect 20812 4150 20864 4156
rect 20626 4111 20682 4120
rect 20260 4072 20312 4078
rect 20536 4072 20588 4078
rect 20260 4014 20312 4020
rect 20442 4040 20498 4049
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 19982 3088 20038 3097
rect 19982 3023 19984 3032
rect 20036 3023 20038 3032
rect 19984 2994 20036 3000
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 20088 2446 20116 2790
rect 20076 2440 20128 2446
rect 20076 2382 20128 2388
rect 20180 1986 20208 3538
rect 20272 2990 20300 4014
rect 20536 4014 20588 4020
rect 20442 3975 20444 3984
rect 20496 3975 20498 3984
rect 20444 3946 20496 3952
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20180 1958 20300 1986
rect 20272 800 20300 1958
rect 20640 800 20668 2994
rect 20824 2650 20852 4150
rect 20916 3602 20944 4644
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 20916 2582 20944 3538
rect 21008 3058 21036 8026
rect 21100 6361 21128 8298
rect 21192 7698 21220 11494
rect 21270 11455 21326 11464
rect 21284 11082 21312 11455
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21270 10704 21326 10713
rect 21270 10639 21272 10648
rect 21324 10639 21326 10648
rect 21272 10610 21324 10616
rect 21272 8968 21324 8974
rect 21270 8936 21272 8945
rect 21324 8936 21326 8945
rect 21270 8871 21326 8880
rect 21376 8838 21404 12406
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 21376 8566 21404 8774
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21270 8256 21326 8265
rect 21270 8191 21326 8200
rect 21284 7818 21312 8191
rect 21468 8090 21496 16079
rect 21560 15094 21588 19178
rect 21548 15088 21600 15094
rect 21548 15030 21600 15036
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21560 12753 21588 13874
rect 21652 13802 21680 20538
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 22006 18184 22062 18193
rect 22062 18142 22140 18170
rect 22006 18119 22062 18128
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21640 13796 21692 13802
rect 21640 13738 21692 13744
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21546 12744 21602 12753
rect 21546 12679 21602 12688
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21456 8084 21508 8090
rect 21456 8026 21508 8032
rect 21272 7812 21324 7818
rect 21272 7754 21324 7760
rect 21192 7670 21312 7698
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21086 6352 21142 6361
rect 21086 6287 21142 6296
rect 21086 5128 21142 5137
rect 21086 5063 21088 5072
rect 21140 5063 21142 5072
rect 21088 5034 21140 5040
rect 20996 3052 21048 3058
rect 20996 2994 21048 3000
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 21192 2378 21220 7414
rect 21284 7342 21312 7670
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21284 7002 21312 7278
rect 21362 7032 21418 7041
rect 21272 6996 21324 7002
rect 21362 6967 21418 6976
rect 21272 6938 21324 6944
rect 21284 5778 21312 6938
rect 21272 5772 21324 5778
rect 21272 5714 21324 5720
rect 21376 5302 21404 6967
rect 21560 5710 21588 11698
rect 22112 11354 22140 18142
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21560 5409 21588 5646
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21546 5400 21602 5409
rect 21742 5403 22050 5412
rect 21546 5335 21602 5344
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 21560 3534 21588 5335
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 21548 3528 21600 3534
rect 21548 3470 21600 3476
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 21180 2372 21232 2378
rect 21180 2314 21232 2320
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 17420 734 17632 762
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
<< via2 >>
rect 2962 21256 3018 21312
rect 1950 20848 2006 20904
rect 1490 20032 1546 20088
rect 2042 20440 2098 20496
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 2686 19896 2742 19952
rect 1490 19660 1492 19680
rect 1492 19660 1544 19680
rect 1544 19660 1546 19680
rect 1490 19624 1546 19660
rect 1214 19488 1270 19544
rect 938 18672 994 18728
rect 1030 18536 1086 18592
rect 1030 17720 1086 17776
rect 938 5788 940 5808
rect 940 5788 992 5808
rect 992 5788 994 5808
rect 938 5752 994 5788
rect 938 4972 940 4992
rect 940 4972 992 4992
rect 992 4972 994 4992
rect 938 4936 994 4972
rect 1122 17040 1178 17096
rect 2042 19236 2098 19272
rect 2042 19216 2044 19236
rect 2044 19216 2096 19236
rect 2096 19216 2098 19236
rect 1490 18808 1546 18864
rect 1490 18400 1546 18456
rect 1306 18128 1362 18184
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 1490 17176 1546 17232
rect 1490 16768 1546 16824
rect 1398 16516 1454 16552
rect 1398 16496 1400 16516
rect 1400 16496 1452 16516
rect 1452 16496 1454 16516
rect 1490 16396 1492 16416
rect 1492 16396 1544 16416
rect 1544 16396 1546 16416
rect 1490 16360 1546 16396
rect 1490 15544 1546 15600
rect 1490 15444 1492 15464
rect 1492 15444 1544 15464
rect 1544 15444 1546 15464
rect 1490 15408 1546 15444
rect 1490 15136 1546 15192
rect 1490 14764 1492 14784
rect 1492 14764 1544 14784
rect 1544 14764 1546 14784
rect 1490 14728 1546 14764
rect 1490 13912 1546 13968
rect 1490 13504 1546 13560
rect 1490 13132 1492 13152
rect 1492 13132 1544 13152
rect 1544 13132 1546 13152
rect 1490 13096 1546 13132
rect 2042 17584 2098 17640
rect 2042 15972 2098 16008
rect 2042 15952 2044 15972
rect 2044 15952 2096 15972
rect 2096 15952 2098 15972
rect 2318 17176 2374 17232
rect 2226 15544 2282 15600
rect 2042 14320 2098 14376
rect 2686 16904 2742 16960
rect 2226 11464 2282 11520
rect 1490 6568 1546 6624
rect 1950 8200 2006 8256
rect 1582 6296 1638 6352
rect 2226 8608 2282 8664
rect 2226 8200 2282 8256
rect 2318 7928 2374 7984
rect 2318 7248 2374 7304
rect 1858 5772 1914 5808
rect 1858 5752 1860 5772
rect 1860 5752 1912 5772
rect 1912 5752 1914 5772
rect 1674 5616 1730 5672
rect 1582 3576 1638 3632
rect 2226 4564 2228 4584
rect 2228 4564 2280 4584
rect 2280 4564 2282 4584
rect 2226 4528 2282 4564
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 4158 19896 4214 19952
rect 3882 19760 3938 19816
rect 3238 17620 3240 17640
rect 3240 17620 3292 17640
rect 3292 17620 3294 17640
rect 3238 17584 3294 17620
rect 3238 16088 3294 16144
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3974 18028 3976 18048
rect 3976 18028 4028 18048
rect 4028 18028 4030 18048
rect 3974 17992 4030 18028
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3698 15988 3700 16008
rect 3700 15988 3752 16008
rect 3752 15988 3754 16008
rect 3238 15308 3240 15328
rect 3240 15308 3292 15328
rect 3292 15308 3294 15328
rect 3238 15272 3294 15308
rect 3698 15952 3754 15988
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 2870 12824 2926 12880
rect 2778 12280 2834 12336
rect 3054 12552 3110 12608
rect 3514 14884 3570 14920
rect 3514 14864 3516 14884
rect 3516 14864 3568 14884
rect 3568 14864 3570 14884
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3330 12824 3386 12880
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 2870 11872 2926 11928
rect 2778 10240 2834 10296
rect 4066 13640 4122 13696
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 4066 12688 4122 12744
rect 4342 12724 4344 12744
rect 4344 12724 4396 12744
rect 4396 12724 4398 12744
rect 4342 12688 4398 12724
rect 4526 16940 4528 16960
rect 4528 16940 4580 16960
rect 4580 16940 4582 16960
rect 4526 16904 4582 16940
rect 4710 15272 4766 15328
rect 6826 19760 6882 19816
rect 5262 19488 5318 19544
rect 4526 12980 4582 13016
rect 4526 12960 4528 12980
rect 4528 12960 4580 12980
rect 4580 12960 4582 12980
rect 4526 12552 4582 12608
rect 3238 11056 3294 11112
rect 4342 11600 4398 11656
rect 2778 9832 2834 9888
rect 2502 4120 2558 4176
rect 2686 6996 2742 7032
rect 2686 6976 2688 6996
rect 2688 6976 2740 6996
rect 2740 6976 2742 6996
rect 3238 9424 3294 9480
rect 2870 7384 2926 7440
rect 3882 10684 3884 10704
rect 3884 10684 3936 10704
rect 3936 10684 3938 10704
rect 3882 10648 3938 10684
rect 3422 10512 3478 10568
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3514 10104 3570 10160
rect 3330 7404 3386 7440
rect 3330 7384 3332 7404
rect 3332 7384 3384 7404
rect 3384 7384 3386 7404
rect 2778 4548 2834 4584
rect 2778 4528 2780 4548
rect 2780 4528 2832 4548
rect 2832 4528 2834 4548
rect 3146 7248 3202 7304
rect 3698 9460 3700 9480
rect 3700 9460 3752 9480
rect 3752 9460 3754 9480
rect 3698 9424 3754 9460
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3882 9016 3938 9072
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3974 7828 3976 7848
rect 3976 7828 4028 7848
rect 4028 7828 4030 7848
rect 3974 7792 4030 7828
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3790 6704 3846 6760
rect 3422 6160 3478 6216
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3330 5228 3386 5264
rect 3330 5208 3332 5228
rect 3332 5208 3384 5228
rect 3384 5208 3386 5228
rect 2778 3712 2834 3768
rect 3054 4664 3110 4720
rect 2410 2896 2466 2952
rect 2226 2372 2282 2408
rect 2226 2352 2228 2372
rect 2228 2352 2280 2372
rect 2280 2352 2282 2372
rect 2870 1672 2926 1728
rect 3974 5616 4030 5672
rect 4158 8472 4214 8528
rect 4250 8372 4252 8392
rect 4252 8372 4304 8392
rect 4304 8372 4306 8392
rect 4250 8336 4306 8372
rect 4894 14356 4896 14376
rect 4896 14356 4948 14376
rect 4948 14356 4950 14376
rect 4894 14320 4950 14356
rect 4802 12416 4858 12472
rect 4802 12180 4804 12200
rect 4804 12180 4856 12200
rect 4856 12180 4858 12200
rect 4802 12144 4858 12180
rect 4618 11464 4674 11520
rect 4434 9152 4490 9208
rect 4158 5480 4214 5536
rect 3422 4936 3478 4992
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3790 4256 3846 4312
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3974 3304 4030 3360
rect 4342 5888 4398 5944
rect 4158 3440 4214 3496
rect 4986 12416 5042 12472
rect 4894 9560 4950 9616
rect 5078 11056 5134 11112
rect 5078 10648 5134 10704
rect 5446 13776 5502 13832
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 5998 17720 6054 17776
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 5538 13368 5594 13424
rect 5354 11772 5356 11792
rect 5356 11772 5408 11792
rect 5408 11772 5410 11792
rect 5354 11736 5410 11772
rect 5446 11636 5448 11656
rect 5448 11636 5500 11656
rect 5500 11636 5502 11656
rect 5446 11600 5502 11636
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6642 16632 6698 16688
rect 7378 19896 7434 19952
rect 6918 19352 6974 19408
rect 7378 19352 7434 19408
rect 7010 18300 7012 18320
rect 7012 18300 7064 18320
rect 7064 18300 7066 18320
rect 7010 18264 7066 18300
rect 7102 17584 7158 17640
rect 6918 16904 6974 16960
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 5814 11464 5870 11520
rect 5446 10240 5502 10296
rect 5262 7656 5318 7712
rect 4618 5888 4674 5944
rect 5170 6180 5226 6216
rect 5170 6160 5172 6180
rect 5172 6160 5224 6180
rect 5224 6160 5226 6180
rect 4618 4428 4620 4448
rect 4620 4428 4672 4448
rect 4672 4428 4674 4448
rect 4618 4392 4674 4428
rect 4618 3848 4674 3904
rect 4618 3576 4674 3632
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3974 2524 3976 2544
rect 3976 2524 4028 2544
rect 4028 2524 4030 2544
rect 3974 2488 4030 2524
rect 3974 2080 4030 2136
rect 4894 3848 4950 3904
rect 4434 1944 4490 2000
rect 5722 9016 5778 9072
rect 5354 6976 5410 7032
rect 6090 14592 6146 14648
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 5998 10668 6054 10704
rect 5998 10648 6000 10668
rect 6000 10648 6052 10668
rect 6052 10648 6054 10668
rect 5814 8336 5870 8392
rect 6734 15816 6790 15872
rect 6918 16360 6974 16416
rect 6826 15136 6882 15192
rect 6826 14728 6882 14784
rect 6642 13504 6698 13560
rect 6642 12588 6644 12608
rect 6644 12588 6696 12608
rect 6696 12588 6698 12608
rect 6642 12552 6698 12588
rect 6826 12552 6882 12608
rect 7102 14456 7158 14512
rect 6826 11600 6882 11656
rect 6642 10512 6698 10568
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 5998 9016 6054 9072
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 5722 6840 5778 6896
rect 4986 2896 5042 2952
rect 6826 8472 6882 8528
rect 5906 5480 5962 5536
rect 6734 7792 6790 7848
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6366 6296 6422 6352
rect 6366 5652 6368 5672
rect 6368 5652 6420 5672
rect 6420 5652 6422 5672
rect 6366 5616 6422 5652
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6458 4684 6514 4720
rect 6458 4664 6460 4684
rect 6460 4664 6512 4684
rect 6512 4664 6514 4684
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 5722 4120 5778 4176
rect 6090 4004 6146 4040
rect 6090 3984 6092 4004
rect 6092 3984 6144 4004
rect 6144 3984 6146 4004
rect 5998 3576 6054 3632
rect 6458 3576 6514 3632
rect 6734 5616 6790 5672
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6090 3052 6146 3088
rect 6090 3032 6092 3052
rect 6092 3032 6144 3052
rect 6144 3032 6146 3052
rect 7378 16088 7434 16144
rect 7470 15544 7526 15600
rect 7470 14612 7526 14648
rect 7470 14592 7472 14612
rect 7472 14592 7524 14612
rect 7524 14592 7526 14612
rect 7102 10956 7104 10976
rect 7104 10956 7156 10976
rect 7156 10956 7158 10976
rect 7102 10920 7158 10956
rect 7102 10104 7158 10160
rect 7562 13776 7618 13832
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8298 19896 8354 19952
rect 8298 18692 8354 18728
rect 8298 18672 8300 18692
rect 8300 18672 8352 18692
rect 8352 18672 8354 18692
rect 7930 16668 7932 16688
rect 7932 16668 7984 16688
rect 7984 16668 7986 16688
rect 7930 16632 7986 16668
rect 7102 8336 7158 8392
rect 7010 5888 7066 5944
rect 7470 10240 7526 10296
rect 7470 9988 7526 10024
rect 7470 9968 7472 9988
rect 7472 9968 7524 9988
rect 7524 9968 7526 9988
rect 6366 2488 6422 2544
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 7562 6432 7618 6488
rect 8206 16088 8262 16144
rect 8206 15000 8262 15056
rect 8206 14048 8262 14104
rect 8206 13252 8262 13288
rect 8206 13232 8208 13252
rect 8208 13232 8260 13252
rect 8260 13232 8262 13252
rect 7746 6840 7802 6896
rect 7470 4392 7526 4448
rect 7470 3984 7526 4040
rect 7654 2624 7710 2680
rect 8206 10512 8262 10568
rect 8206 8508 8208 8528
rect 8208 8508 8260 8528
rect 8260 8508 8262 8528
rect 8206 8472 8262 8508
rect 8206 7248 8262 7304
rect 8114 6432 8170 6488
rect 8114 6332 8116 6352
rect 8116 6332 8168 6352
rect 8168 6332 8170 6352
rect 8114 6296 8170 6332
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8482 14764 8484 14784
rect 8484 14764 8536 14784
rect 8536 14764 8538 14784
rect 8482 14728 8538 14764
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8758 15564 8814 15600
rect 8758 15544 8760 15564
rect 8760 15544 8812 15564
rect 8812 15544 8814 15564
rect 9034 15000 9090 15056
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 9218 18128 9274 18184
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8666 12280 8722 12336
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 9678 18844 9680 18864
rect 9680 18844 9732 18864
rect 9732 18844 9734 18864
rect 9678 18808 9734 18844
rect 9402 15272 9458 15328
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8666 10104 8722 10160
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8758 8628 8814 8664
rect 8758 8608 8760 8628
rect 8760 8608 8812 8628
rect 8812 8608 8814 8628
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8574 7520 8630 7576
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8574 4392 8630 4448
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9126 4428 9128 4448
rect 9128 4428 9180 4448
rect 9180 4428 9182 4448
rect 9126 4392 9182 4428
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8206 3304 8262 3360
rect 8482 3032 8538 3088
rect 9034 2932 9036 2952
rect 9036 2932 9088 2952
rect 9088 2932 9090 2952
rect 9034 2896 9090 2932
rect 8574 2796 8576 2816
rect 8576 2796 8628 2816
rect 8628 2796 8630 2816
rect 8574 2760 8630 2796
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 8850 2488 8906 2544
rect 9586 13368 9642 13424
rect 9494 11056 9550 11112
rect 10138 17484 10140 17504
rect 10140 17484 10192 17504
rect 10192 17484 10194 17504
rect 10138 17448 10194 17484
rect 9954 16668 9956 16688
rect 9956 16668 10008 16688
rect 10008 16668 10010 16688
rect 9954 16632 10010 16668
rect 10046 15408 10102 15464
rect 10046 15136 10102 15192
rect 10782 19760 10838 19816
rect 10414 17856 10470 17912
rect 10322 16652 10378 16688
rect 10322 16632 10324 16652
rect 10324 16632 10376 16652
rect 10376 16632 10378 16652
rect 9494 8628 9550 8664
rect 9494 8608 9496 8628
rect 9496 8608 9548 8628
rect 9548 8608 9550 8628
rect 9494 8336 9550 8392
rect 9310 7112 9366 7168
rect 9494 6840 9550 6896
rect 9678 8200 9734 8256
rect 10138 8200 10194 8256
rect 9954 7792 10010 7848
rect 9310 5888 9366 5944
rect 9954 6976 10010 7032
rect 9310 4120 9366 4176
rect 9954 4256 10010 4312
rect 10322 10512 10378 10568
rect 10782 16768 10838 16824
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 10966 17992 11022 18048
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11794 19372 11850 19408
rect 11794 19352 11796 19372
rect 11796 19352 11848 19372
rect 11848 19352 11850 19372
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 17958 21256 18014 21312
rect 20626 20848 20682 20904
rect 11978 19352 12034 19408
rect 11794 18672 11850 18728
rect 11518 17076 11520 17096
rect 11520 17076 11572 17096
rect 11572 17076 11574 17096
rect 11518 17040 11574 17076
rect 11702 17040 11758 17096
rect 10874 14728 10930 14784
rect 10782 10920 10838 10976
rect 11702 16496 11758 16552
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11334 15544 11390 15600
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11058 14456 11114 14512
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11702 13640 11758 13696
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11150 11192 11206 11248
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11058 10784 11114 10840
rect 11150 10648 11206 10704
rect 11242 10240 11298 10296
rect 12254 19236 12310 19272
rect 12254 19216 12256 19236
rect 12256 19216 12308 19236
rect 12308 19216 12310 19236
rect 11978 18128 12034 18184
rect 12162 14764 12164 14784
rect 12164 14764 12216 14784
rect 12216 14764 12218 14784
rect 12162 14728 12218 14764
rect 12898 19252 12900 19272
rect 12900 19252 12952 19272
rect 12952 19252 12954 19272
rect 12898 19216 12954 19252
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 12898 18672 12954 18728
rect 12898 18400 12954 18456
rect 12346 15544 12402 15600
rect 12438 14456 12494 14512
rect 11978 12416 12034 12472
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 10322 3032 10378 3088
rect 11058 7248 11114 7304
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11702 5888 11758 5944
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11058 3984 11114 4040
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 10598 2624 10654 2680
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12254 12280 12310 12336
rect 11978 11056 12034 11112
rect 12070 10376 12126 10432
rect 12254 9560 12310 9616
rect 12438 10784 12494 10840
rect 12162 5752 12218 5808
rect 11978 2896 12034 2952
rect 12254 2644 12310 2680
rect 12254 2624 12256 2644
rect 12256 2624 12308 2644
rect 12308 2624 12310 2644
rect 13082 16652 13138 16688
rect 13082 16632 13084 16652
rect 13084 16632 13136 16652
rect 13136 16632 13138 16652
rect 13358 17992 13414 18048
rect 13266 17720 13322 17776
rect 12714 10240 12770 10296
rect 12898 9968 12954 10024
rect 12806 7928 12862 7984
rect 12622 7268 12678 7304
rect 12622 7248 12624 7268
rect 12624 7248 12676 7268
rect 12676 7248 12678 7268
rect 12530 6704 12586 6760
rect 12530 3576 12586 3632
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 14370 18264 14426 18320
rect 14370 17176 14426 17232
rect 13358 15272 13414 15328
rect 12990 7792 13046 7848
rect 13358 11192 13414 11248
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13726 12552 13782 12608
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13542 11736 13598 11792
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 14462 16496 14518 16552
rect 14462 12280 14518 12336
rect 14646 15852 14648 15872
rect 14648 15852 14700 15872
rect 14700 15852 14702 15872
rect 14646 15816 14702 15852
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13450 9968 13506 10024
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13634 7404 13690 7440
rect 13634 7384 13636 7404
rect 13636 7384 13688 7404
rect 13688 7384 13690 7404
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 14462 7112 14518 7168
rect 15290 18672 15346 18728
rect 15014 17856 15070 17912
rect 14830 12824 14886 12880
rect 15382 17040 15438 17096
rect 15106 12688 15162 12744
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16118 15952 16174 16008
rect 16118 15000 16174 15056
rect 15566 12688 15622 12744
rect 15014 11056 15070 11112
rect 14830 6740 14832 6760
rect 14832 6740 14884 6760
rect 14884 6740 14886 6760
rect 14830 6704 14886 6740
rect 14462 5208 14518 5264
rect 14278 3984 14334 4040
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 15014 7248 15070 7304
rect 15198 6976 15254 7032
rect 15290 6296 15346 6352
rect 15290 5888 15346 5944
rect 14922 4936 14978 4992
rect 14830 3460 14886 3496
rect 14830 3440 14832 3460
rect 14832 3440 14884 3460
rect 14884 3440 14886 3460
rect 14554 2896 14610 2952
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 15290 4528 15346 4584
rect 15566 9324 15568 9344
rect 15568 9324 15620 9344
rect 15620 9324 15622 9344
rect 15566 9288 15622 9324
rect 15566 6024 15622 6080
rect 16946 19388 16948 19408
rect 16948 19388 17000 19408
rect 17000 19388 17002 19408
rect 16946 19352 17002 19388
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16946 17584 17002 17640
rect 16118 5652 16120 5672
rect 16120 5652 16172 5672
rect 16172 5652 16174 5672
rect 16118 5616 16174 5652
rect 16118 4664 16174 4720
rect 15934 3984 15990 4040
rect 16302 4528 16358 4584
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16946 14184 17002 14240
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16486 12588 16488 12608
rect 16488 12588 16540 12608
rect 16540 12588 16542 12608
rect 16486 12552 16542 12588
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16946 9968 17002 10024
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 17314 15408 17370 15464
rect 17774 16652 17830 16688
rect 17774 16632 17776 16652
rect 17776 16632 17828 16652
rect 17828 16632 17830 16652
rect 17682 14320 17738 14376
rect 17314 12552 17370 12608
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16578 6704 16634 6760
rect 16946 6604 16948 6624
rect 16948 6604 17000 6624
rect 17000 6604 17002 6624
rect 16946 6568 17002 6604
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16854 5772 16910 5808
rect 16854 5752 16856 5772
rect 16856 5752 16908 5772
rect 16908 5752 16910 5772
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 17590 11872 17646 11928
rect 17406 9152 17462 9208
rect 18142 15972 18198 16008
rect 18142 15952 18144 15972
rect 18144 15952 18196 15972
rect 18196 15952 18198 15972
rect 17774 12552 17830 12608
rect 18142 12280 18198 12336
rect 18418 17720 18474 17776
rect 18694 18708 18696 18728
rect 18696 18708 18748 18728
rect 18748 18708 18750 18728
rect 18694 18672 18750 18708
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19706 19896 19762 19952
rect 18602 17856 18658 17912
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 20166 20440 20222 20496
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 20718 20032 20774 20088
rect 19890 17720 19946 17776
rect 19798 17584 19854 17640
rect 17958 11056 18014 11112
rect 17958 9288 18014 9344
rect 17866 9152 17922 9208
rect 16946 4664 17002 4720
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 15934 3052 15990 3088
rect 15934 3032 15936 3052
rect 15936 3032 15988 3052
rect 15988 3032 15990 3052
rect 16302 2896 16358 2952
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 17682 6160 17738 6216
rect 17590 5364 17646 5400
rect 17590 5344 17592 5364
rect 17592 5344 17644 5364
rect 17644 5344 17646 5364
rect 17498 4664 17554 4720
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 18878 16632 18934 16688
rect 18786 12724 18788 12744
rect 18788 12724 18840 12744
rect 18840 12724 18842 12744
rect 18786 12688 18842 12724
rect 18602 12144 18658 12200
rect 18694 11092 18696 11112
rect 18696 11092 18748 11112
rect 18748 11092 18750 11112
rect 18694 11056 18750 11092
rect 18050 6432 18106 6488
rect 18234 6432 18290 6488
rect 17958 6024 18014 6080
rect 18418 7384 18474 7440
rect 18510 6976 18566 7032
rect 18326 5752 18382 5808
rect 18142 5344 18198 5400
rect 18050 4936 18106 4992
rect 18142 4664 18198 4720
rect 18510 6160 18566 6216
rect 18694 7828 18696 7848
rect 18696 7828 18748 7848
rect 18748 7828 18750 7848
rect 18694 7792 18750 7828
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19614 15000 19670 15056
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19062 9424 19118 9480
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19890 15544 19946 15600
rect 20166 18128 20222 18184
rect 20166 16632 20222 16688
rect 19890 13232 19946 13288
rect 19798 11892 19854 11928
rect 19798 11872 19800 11892
rect 19800 11872 19852 11892
rect 19852 11872 19854 11892
rect 18050 3440 18106 3496
rect 17866 3032 17922 3088
rect 17498 1944 17554 2000
rect 18970 7112 19026 7168
rect 18878 5752 18934 5808
rect 18878 5208 18934 5264
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19246 6704 19302 6760
rect 19246 6296 19302 6352
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 20166 14728 20222 14784
rect 21270 19760 21326 19816
rect 20626 19216 20682 19272
rect 21270 18808 21326 18864
rect 21178 18672 21234 18728
rect 20718 17584 20774 17640
rect 20718 16768 20774 16824
rect 20902 16904 20958 16960
rect 20534 16496 20590 16552
rect 21362 18264 21418 18320
rect 21270 17992 21326 18048
rect 21362 17176 21418 17232
rect 20718 14320 20774 14376
rect 19982 10124 20038 10160
rect 19982 10104 19984 10124
rect 19984 10104 20036 10124
rect 20036 10104 20038 10124
rect 20166 10240 20222 10296
rect 19614 6296 19670 6352
rect 19154 5480 19210 5536
rect 19982 6840 20038 6896
rect 19614 5616 19670 5672
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 18602 2896 18658 2952
rect 18970 1672 19026 1728
rect 19246 3576 19302 3632
rect 19154 3032 19210 3088
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19246 2488 19302 2544
rect 19614 3712 19670 3768
rect 20534 12280 20590 12336
rect 20534 9968 20590 10024
rect 20442 9560 20498 9616
rect 20534 9016 20590 9072
rect 19890 4936 19946 4992
rect 21454 16496 21510 16552
rect 21454 16088 21510 16144
rect 21270 15952 21326 16008
rect 21362 13912 21418 13968
rect 21270 13504 21326 13560
rect 21178 12824 21234 12880
rect 21270 11736 21326 11792
rect 20902 9152 20958 9208
rect 20810 8472 20866 8528
rect 20534 7384 20590 7440
rect 21086 8900 21142 8936
rect 21086 8880 21088 8900
rect 21088 8880 21140 8900
rect 21140 8880 21142 8900
rect 20718 6704 20774 6760
rect 20810 6296 20866 6352
rect 20626 4120 20682 4176
rect 19982 3052 20038 3088
rect 19982 3032 19984 3052
rect 19984 3032 20036 3052
rect 20036 3032 20038 3052
rect 20442 4004 20498 4040
rect 20442 3984 20444 4004
rect 20444 3984 20496 4004
rect 20496 3984 20498 4004
rect 21270 11464 21326 11520
rect 21270 10668 21326 10704
rect 21270 10648 21272 10668
rect 21272 10648 21324 10668
rect 21324 10648 21326 10668
rect 21270 8916 21272 8936
rect 21272 8916 21324 8936
rect 21324 8916 21326 8936
rect 21270 8880 21326 8916
rect 21270 8200 21326 8256
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 22006 18128 22062 18184
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21546 12688 21602 12744
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21086 6296 21142 6352
rect 21086 5092 21142 5128
rect 21086 5072 21088 5092
rect 21088 5072 21140 5092
rect 21140 5072 21142 5092
rect 21362 6976 21418 7032
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21546 5344 21602 5400
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 0 21314 800 21344
rect 2957 21314 3023 21317
rect 0 21312 3023 21314
rect 0 21256 2962 21312
rect 3018 21256 3023 21312
rect 0 21254 3023 21256
rect 0 21224 800 21254
rect 2957 21251 3023 21254
rect 17953 21314 18019 21317
rect 22200 21314 23000 21344
rect 17953 21312 23000 21314
rect 17953 21256 17958 21312
rect 18014 21256 23000 21312
rect 17953 21254 23000 21256
rect 17953 21251 18019 21254
rect 22200 21224 23000 21254
rect 0 20906 800 20936
rect 1945 20906 2011 20909
rect 0 20904 2011 20906
rect 0 20848 1950 20904
rect 2006 20848 2011 20904
rect 0 20846 2011 20848
rect 0 20816 800 20846
rect 1945 20843 2011 20846
rect 20621 20906 20687 20909
rect 22200 20906 23000 20936
rect 20621 20904 23000 20906
rect 20621 20848 20626 20904
rect 20682 20848 23000 20904
rect 20621 20846 23000 20848
rect 20621 20843 20687 20846
rect 22200 20816 23000 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 0 20498 800 20528
rect 2037 20498 2103 20501
rect 0 20496 2103 20498
rect 0 20440 2042 20496
rect 2098 20440 2103 20496
rect 0 20438 2103 20440
rect 0 20408 800 20438
rect 2037 20435 2103 20438
rect 20161 20498 20227 20501
rect 22200 20498 23000 20528
rect 20161 20496 23000 20498
rect 20161 20440 20166 20496
rect 20222 20440 23000 20496
rect 20161 20438 23000 20440
rect 20161 20435 20227 20438
rect 22200 20408 23000 20438
rect 3545 20160 3861 20161
rect 0 20090 800 20120
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 1485 20090 1551 20093
rect 0 20088 1551 20090
rect 0 20032 1490 20088
rect 1546 20032 1551 20088
rect 0 20030 1551 20032
rect 0 20000 800 20030
rect 1485 20027 1551 20030
rect 20713 20090 20779 20093
rect 22200 20090 23000 20120
rect 20713 20088 23000 20090
rect 20713 20032 20718 20088
rect 20774 20032 23000 20088
rect 20713 20030 23000 20032
rect 20713 20027 20779 20030
rect 22200 20000 23000 20030
rect 2681 19954 2747 19957
rect 4153 19954 4219 19957
rect 7373 19954 7439 19957
rect 2681 19952 7439 19954
rect 2681 19896 2686 19952
rect 2742 19896 4158 19952
rect 4214 19896 7378 19952
rect 7434 19896 7439 19952
rect 2681 19894 7439 19896
rect 2681 19891 2747 19894
rect 4153 19891 4219 19894
rect 7373 19891 7439 19894
rect 8293 19954 8359 19957
rect 19701 19954 19767 19957
rect 8293 19952 19767 19954
rect 8293 19896 8298 19952
rect 8354 19896 19706 19952
rect 19762 19896 19767 19952
rect 8293 19894 19767 19896
rect 8293 19891 8359 19894
rect 19701 19891 19767 19894
rect 3877 19818 3943 19821
rect 6821 19818 6887 19821
rect 10777 19818 10843 19821
rect 16246 19818 16252 19820
rect 3877 19816 16252 19818
rect 3877 19760 3882 19816
rect 3938 19760 6826 19816
rect 6882 19760 10782 19816
rect 10838 19760 16252 19816
rect 3877 19758 16252 19760
rect 3877 19755 3943 19758
rect 6821 19755 6887 19758
rect 10777 19755 10843 19758
rect 16246 19756 16252 19758
rect 16316 19756 16322 19820
rect 21265 19818 21331 19821
rect 21265 19816 22202 19818
rect 21265 19760 21270 19816
rect 21326 19760 22202 19816
rect 21265 19758 22202 19760
rect 21265 19755 21331 19758
rect 22142 19712 22202 19758
rect 0 19682 800 19712
rect 1485 19682 1551 19685
rect 0 19680 1551 19682
rect 0 19624 1490 19680
rect 1546 19624 1551 19680
rect 0 19622 1551 19624
rect 22142 19622 23000 19712
rect 0 19592 800 19622
rect 1485 19619 1551 19622
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 22200 19592 23000 19622
rect 21738 19551 22054 19552
rect 1209 19546 1275 19549
rect 5257 19546 5323 19549
rect 1209 19544 5323 19546
rect 1209 19488 1214 19544
rect 1270 19488 5262 19544
rect 5318 19488 5323 19544
rect 1209 19486 5323 19488
rect 1209 19483 1275 19486
rect 5257 19483 5323 19486
rect 3918 19348 3924 19412
rect 3988 19410 3994 19412
rect 6913 19410 6979 19413
rect 3988 19408 6979 19410
rect 3988 19352 6918 19408
rect 6974 19352 6979 19408
rect 3988 19350 6979 19352
rect 3988 19348 3994 19350
rect 6913 19347 6979 19350
rect 7373 19410 7439 19413
rect 11789 19410 11855 19413
rect 7373 19408 11855 19410
rect 7373 19352 7378 19408
rect 7434 19352 11794 19408
rect 11850 19352 11855 19408
rect 7373 19350 11855 19352
rect 7373 19347 7439 19350
rect 11789 19347 11855 19350
rect 11973 19410 12039 19413
rect 16941 19412 17007 19413
rect 15142 19410 15148 19412
rect 11973 19408 15148 19410
rect 11973 19352 11978 19408
rect 12034 19352 15148 19408
rect 11973 19350 15148 19352
rect 11973 19347 12039 19350
rect 15142 19348 15148 19350
rect 15212 19348 15218 19412
rect 16941 19408 16988 19412
rect 17052 19410 17058 19412
rect 16941 19352 16946 19408
rect 16941 19348 16988 19352
rect 17052 19350 17098 19410
rect 17052 19348 17058 19350
rect 16941 19347 17007 19348
rect 0 19274 800 19304
rect 2037 19274 2103 19277
rect 0 19272 2103 19274
rect 0 19216 2042 19272
rect 2098 19216 2103 19272
rect 0 19214 2103 19216
rect 0 19184 800 19214
rect 2037 19211 2103 19214
rect 12249 19274 12315 19277
rect 12893 19274 12959 19277
rect 12249 19272 12959 19274
rect 12249 19216 12254 19272
rect 12310 19216 12898 19272
rect 12954 19216 12959 19272
rect 12249 19214 12959 19216
rect 12249 19211 12315 19214
rect 12893 19211 12959 19214
rect 20621 19274 20687 19277
rect 22200 19274 23000 19304
rect 20621 19272 23000 19274
rect 20621 19216 20626 19272
rect 20682 19216 23000 19272
rect 20621 19214 23000 19216
rect 20621 19211 20687 19214
rect 22200 19184 23000 19214
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 0 18866 800 18896
rect 1485 18866 1551 18869
rect 9673 18866 9739 18869
rect 0 18864 1551 18866
rect 0 18808 1490 18864
rect 1546 18808 1551 18864
rect 0 18806 1551 18808
rect 0 18776 800 18806
rect 1485 18803 1551 18806
rect 1718 18864 9739 18866
rect 1718 18808 9678 18864
rect 9734 18808 9739 18864
rect 1718 18806 9739 18808
rect 933 18730 999 18733
rect 1718 18730 1778 18806
rect 9673 18803 9739 18806
rect 21265 18866 21331 18869
rect 22200 18866 23000 18896
rect 21265 18864 23000 18866
rect 21265 18808 21270 18864
rect 21326 18808 23000 18864
rect 21265 18806 23000 18808
rect 21265 18803 21331 18806
rect 22200 18776 23000 18806
rect 8293 18730 8359 18733
rect 933 18728 1778 18730
rect 933 18672 938 18728
rect 994 18672 1778 18728
rect 933 18670 1778 18672
rect 1902 18728 8359 18730
rect 1902 18672 8298 18728
rect 8354 18672 8359 18728
rect 1902 18670 8359 18672
rect 933 18667 999 18670
rect 1025 18594 1091 18597
rect 1902 18594 1962 18670
rect 8293 18667 8359 18670
rect 11789 18730 11855 18733
rect 12893 18730 12959 18733
rect 11789 18728 12959 18730
rect 11789 18672 11794 18728
rect 11850 18672 12898 18728
rect 12954 18672 12959 18728
rect 11789 18670 12959 18672
rect 11789 18667 11855 18670
rect 12893 18667 12959 18670
rect 15285 18730 15351 18733
rect 18689 18730 18755 18733
rect 21173 18730 21239 18733
rect 15285 18728 21239 18730
rect 15285 18672 15290 18728
rect 15346 18672 18694 18728
rect 18750 18672 21178 18728
rect 21234 18672 21239 18728
rect 15285 18670 21239 18672
rect 15285 18667 15351 18670
rect 18689 18667 18755 18670
rect 21173 18667 21239 18670
rect 1025 18592 1962 18594
rect 1025 18536 1030 18592
rect 1086 18536 1962 18592
rect 1025 18534 1962 18536
rect 1025 18531 1091 18534
rect 6144 18528 6460 18529
rect 0 18458 800 18488
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 1485 18458 1551 18461
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 12893 18458 12959 18461
rect 22200 18458 23000 18488
rect 12893 18456 14658 18458
rect 12893 18400 12898 18456
rect 12954 18400 14658 18456
rect 12893 18398 14658 18400
rect 12893 18395 12959 18398
rect 5574 18260 5580 18324
rect 5644 18322 5650 18324
rect 7005 18322 7071 18325
rect 5644 18320 7071 18322
rect 5644 18264 7010 18320
rect 7066 18264 7071 18320
rect 5644 18262 7071 18264
rect 5644 18260 5650 18262
rect 7005 18259 7071 18262
rect 8334 18260 8340 18324
rect 8404 18322 8410 18324
rect 14365 18322 14431 18325
rect 8404 18320 14431 18322
rect 8404 18264 14370 18320
rect 14426 18264 14431 18320
rect 8404 18262 14431 18264
rect 14598 18322 14658 18398
rect 22142 18368 23000 18458
rect 21357 18322 21423 18325
rect 22142 18322 22202 18368
rect 14598 18262 20362 18322
rect 8404 18260 8410 18262
rect 14365 18259 14431 18262
rect 1301 18186 1367 18189
rect 9213 18186 9279 18189
rect 1301 18184 9279 18186
rect 1301 18128 1306 18184
rect 1362 18128 9218 18184
rect 9274 18128 9279 18184
rect 1301 18126 9279 18128
rect 1301 18123 1367 18126
rect 9213 18123 9279 18126
rect 11973 18186 12039 18189
rect 20161 18186 20227 18189
rect 11973 18184 20227 18186
rect 11973 18128 11978 18184
rect 12034 18128 20166 18184
rect 20222 18128 20227 18184
rect 11973 18126 20227 18128
rect 20302 18186 20362 18262
rect 21357 18320 22202 18322
rect 21357 18264 21362 18320
rect 21418 18264 22202 18320
rect 21357 18262 22202 18264
rect 21357 18259 21423 18262
rect 22001 18186 22067 18189
rect 20302 18184 22067 18186
rect 20302 18128 22006 18184
rect 22062 18128 22067 18184
rect 20302 18126 22067 18128
rect 11973 18123 12039 18126
rect 20161 18123 20227 18126
rect 22001 18123 22067 18126
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 3969 18050 4035 18053
rect 8150 18050 8156 18052
rect 3969 18048 8156 18050
rect 3969 17992 3974 18048
rect 4030 17992 8156 18048
rect 3969 17990 8156 17992
rect 3969 17987 4035 17990
rect 8150 17988 8156 17990
rect 8220 17988 8226 18052
rect 10961 18050 11027 18053
rect 12198 18050 12204 18052
rect 10961 18048 12204 18050
rect 10961 17992 10966 18048
rect 11022 17992 12204 18048
rect 10961 17990 12204 17992
rect 10961 17987 11027 17990
rect 12198 17988 12204 17990
rect 12268 17988 12274 18052
rect 13353 18050 13419 18053
rect 13486 18050 13492 18052
rect 13353 18048 13492 18050
rect 13353 17992 13358 18048
rect 13414 17992 13492 18048
rect 13353 17990 13492 17992
rect 13353 17987 13419 17990
rect 13486 17988 13492 17990
rect 13556 17988 13562 18052
rect 21265 18050 21331 18053
rect 22200 18050 23000 18080
rect 21265 18048 23000 18050
rect 21265 17992 21270 18048
rect 21326 17992 23000 18048
rect 21265 17990 23000 17992
rect 21265 17987 21331 17990
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 22200 17960 23000 17990
rect 19139 17919 19455 17920
rect 10409 17914 10475 17917
rect 10726 17914 10732 17916
rect 10409 17912 10732 17914
rect 10409 17856 10414 17912
rect 10470 17856 10732 17912
rect 10409 17854 10732 17856
rect 10409 17851 10475 17854
rect 10726 17852 10732 17854
rect 10796 17852 10802 17916
rect 15009 17914 15075 17917
rect 18597 17914 18663 17917
rect 14414 17912 18663 17914
rect 14414 17856 15014 17912
rect 15070 17856 18602 17912
rect 18658 17856 18663 17912
rect 14414 17854 18663 17856
rect 1025 17778 1091 17781
rect 5993 17778 6059 17781
rect 1025 17776 6059 17778
rect 1025 17720 1030 17776
rect 1086 17720 5998 17776
rect 6054 17720 6059 17776
rect 1025 17718 6059 17720
rect 1025 17715 1091 17718
rect 5993 17715 6059 17718
rect 13261 17778 13327 17781
rect 14414 17778 14474 17854
rect 15009 17851 15075 17854
rect 18597 17851 18663 17854
rect 13261 17776 14474 17778
rect 13261 17720 13266 17776
rect 13322 17720 14474 17776
rect 13261 17718 14474 17720
rect 18413 17778 18479 17781
rect 19885 17778 19951 17781
rect 18413 17776 19951 17778
rect 18413 17720 18418 17776
rect 18474 17720 19890 17776
rect 19946 17720 19951 17776
rect 18413 17718 19951 17720
rect 13261 17715 13327 17718
rect 18413 17715 18479 17718
rect 19885 17715 19951 17718
rect 0 17642 800 17672
rect 2037 17642 2103 17645
rect 0 17640 2103 17642
rect 0 17584 2042 17640
rect 2098 17584 2103 17640
rect 0 17582 2103 17584
rect 0 17552 800 17582
rect 2037 17579 2103 17582
rect 3233 17642 3299 17645
rect 7097 17642 7163 17645
rect 3233 17640 7163 17642
rect 3233 17584 3238 17640
rect 3294 17584 7102 17640
rect 7158 17584 7163 17640
rect 3233 17582 7163 17584
rect 3233 17579 3299 17582
rect 7097 17579 7163 17582
rect 16941 17642 17007 17645
rect 19793 17642 19859 17645
rect 16941 17640 19859 17642
rect 16941 17584 16946 17640
rect 17002 17584 19798 17640
rect 19854 17584 19859 17640
rect 16941 17582 19859 17584
rect 16941 17579 17007 17582
rect 19793 17579 19859 17582
rect 20713 17642 20779 17645
rect 22200 17642 23000 17672
rect 20713 17640 23000 17642
rect 20713 17584 20718 17640
rect 20774 17584 23000 17640
rect 20713 17582 23000 17584
rect 20713 17579 20779 17582
rect 22200 17552 23000 17582
rect 8150 17444 8156 17508
rect 8220 17506 8226 17508
rect 10133 17506 10199 17509
rect 8220 17504 10199 17506
rect 8220 17448 10138 17504
rect 10194 17448 10199 17504
rect 8220 17446 10199 17448
rect 8220 17444 8226 17446
rect 10133 17443 10199 17446
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 2313 17234 2379 17237
rect 14365 17234 14431 17237
rect 2313 17232 14431 17234
rect 2313 17176 2318 17232
rect 2374 17176 14370 17232
rect 14426 17176 14431 17232
rect 2313 17174 14431 17176
rect 2313 17171 2379 17174
rect 14365 17171 14431 17174
rect 21357 17234 21423 17237
rect 22200 17234 23000 17264
rect 21357 17232 23000 17234
rect 21357 17176 21362 17232
rect 21418 17176 23000 17232
rect 21357 17174 23000 17176
rect 21357 17171 21423 17174
rect 22200 17144 23000 17174
rect 1117 17098 1183 17101
rect 11513 17098 11579 17101
rect 1117 17096 11579 17098
rect 1117 17040 1122 17096
rect 1178 17040 11518 17096
rect 11574 17040 11579 17096
rect 1117 17038 11579 17040
rect 1117 17035 1183 17038
rect 11513 17035 11579 17038
rect 11697 17098 11763 17101
rect 15377 17098 15443 17101
rect 11697 17096 15443 17098
rect 11697 17040 11702 17096
rect 11758 17040 15382 17096
rect 15438 17040 15443 17096
rect 11697 17038 15443 17040
rect 11697 17035 11763 17038
rect 15377 17035 15443 17038
rect 2681 16964 2747 16965
rect 2630 16962 2636 16964
rect 2590 16902 2636 16962
rect 2700 16960 2747 16964
rect 2742 16904 2747 16960
rect 2630 16900 2636 16902
rect 2700 16900 2747 16904
rect 2681 16899 2747 16900
rect 4521 16962 4587 16965
rect 6913 16962 6979 16965
rect 20897 16962 20963 16965
rect 4521 16960 6979 16962
rect 4521 16904 4526 16960
rect 4582 16904 6918 16960
rect 6974 16904 6979 16960
rect 4521 16902 6979 16904
rect 4521 16899 4587 16902
rect 6913 16899 6979 16902
rect 19934 16960 20963 16962
rect 19934 16904 20902 16960
rect 20958 16904 20963 16960
rect 19934 16902 20963 16904
rect 3545 16896 3861 16897
rect 0 16826 800 16856
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 1485 16826 1551 16829
rect 0 16824 1551 16826
rect 0 16768 1490 16824
rect 1546 16768 1551 16824
rect 0 16766 1551 16768
rect 0 16736 800 16766
rect 1485 16763 1551 16766
rect 10777 16826 10843 16829
rect 10777 16824 13370 16826
rect 10777 16768 10782 16824
rect 10838 16768 13370 16824
rect 10777 16766 13370 16768
rect 10777 16763 10843 16766
rect 5758 16628 5764 16692
rect 5828 16690 5834 16692
rect 6637 16690 6703 16693
rect 7925 16692 7991 16693
rect 9949 16692 10015 16693
rect 10317 16692 10383 16693
rect 13077 16692 13143 16693
rect 7925 16690 7972 16692
rect 5828 16688 6703 16690
rect 5828 16632 6642 16688
rect 6698 16632 6703 16688
rect 5828 16630 6703 16632
rect 7880 16688 7972 16690
rect 7880 16632 7930 16688
rect 7880 16630 7972 16632
rect 5828 16628 5834 16630
rect 6637 16627 6703 16630
rect 7925 16628 7972 16630
rect 8036 16628 8042 16692
rect 9949 16688 9996 16692
rect 10060 16690 10066 16692
rect 9949 16632 9954 16688
rect 9949 16628 9996 16632
rect 10060 16630 10106 16690
rect 10317 16688 10364 16692
rect 10428 16690 10434 16692
rect 10317 16632 10322 16688
rect 10060 16628 10066 16630
rect 10317 16628 10364 16632
rect 10428 16630 10474 16690
rect 13077 16688 13124 16692
rect 13188 16690 13194 16692
rect 13310 16690 13370 16766
rect 17769 16692 17835 16693
rect 14406 16690 14412 16692
rect 13077 16632 13082 16688
rect 10428 16628 10434 16630
rect 13077 16628 13124 16632
rect 13188 16630 13234 16690
rect 13310 16630 14412 16690
rect 13188 16628 13194 16630
rect 14406 16628 14412 16630
rect 14476 16628 14482 16692
rect 17718 16690 17724 16692
rect 17678 16630 17724 16690
rect 17788 16688 17835 16692
rect 17830 16632 17835 16688
rect 17718 16628 17724 16630
rect 17788 16628 17835 16632
rect 7925 16627 7991 16628
rect 9949 16627 10015 16628
rect 10317 16627 10383 16628
rect 13077 16627 13143 16628
rect 17769 16627 17835 16628
rect 18873 16690 18939 16693
rect 19934 16690 19994 16902
rect 20897 16899 20963 16902
rect 20713 16826 20779 16829
rect 22200 16826 23000 16856
rect 20713 16824 23000 16826
rect 20713 16768 20718 16824
rect 20774 16768 23000 16824
rect 20713 16766 23000 16768
rect 20713 16763 20779 16766
rect 22200 16736 23000 16766
rect 18873 16688 19994 16690
rect 18873 16632 18878 16688
rect 18934 16632 19994 16688
rect 18873 16630 19994 16632
rect 20161 16690 20227 16693
rect 20478 16690 20484 16692
rect 20161 16688 20484 16690
rect 20161 16632 20166 16688
rect 20222 16632 20484 16688
rect 20161 16630 20484 16632
rect 18873 16627 18939 16630
rect 20161 16627 20227 16630
rect 20478 16628 20484 16630
rect 20548 16628 20554 16692
rect 1393 16554 1459 16557
rect 11697 16554 11763 16557
rect 1393 16552 11763 16554
rect 1393 16496 1398 16552
rect 1454 16496 11702 16552
rect 11758 16496 11763 16552
rect 1393 16494 11763 16496
rect 1393 16491 1459 16494
rect 11697 16491 11763 16494
rect 14457 16554 14523 16557
rect 20529 16554 20595 16557
rect 14457 16552 20595 16554
rect 14457 16496 14462 16552
rect 14518 16496 20534 16552
rect 20590 16496 20595 16552
rect 14457 16494 20595 16496
rect 14457 16491 14523 16494
rect 20529 16491 20595 16494
rect 21449 16554 21515 16557
rect 21449 16552 22202 16554
rect 21449 16496 21454 16552
rect 21510 16496 22202 16552
rect 21449 16494 22202 16496
rect 21449 16491 21515 16494
rect 22142 16448 22202 16494
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 6913 16418 6979 16421
rect 8518 16418 8524 16420
rect 6913 16416 8524 16418
rect 6913 16360 6918 16416
rect 6974 16360 8524 16416
rect 6913 16358 8524 16360
rect 6913 16355 6979 16358
rect 8518 16356 8524 16358
rect 8588 16356 8594 16420
rect 22142 16358 23000 16448
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 22200 16328 23000 16358
rect 21738 16287 22054 16288
rect 3233 16146 3299 16149
rect 5390 16146 5396 16148
rect 3233 16144 5396 16146
rect 3233 16088 3238 16144
rect 3294 16088 5396 16144
rect 3233 16086 5396 16088
rect 3233 16083 3299 16086
rect 5390 16084 5396 16086
rect 5460 16146 5466 16148
rect 7373 16146 7439 16149
rect 5460 16144 7439 16146
rect 5460 16088 7378 16144
rect 7434 16088 7439 16144
rect 5460 16086 7439 16088
rect 5460 16084 5466 16086
rect 7373 16083 7439 16086
rect 8201 16146 8267 16149
rect 21449 16146 21515 16149
rect 8201 16144 21515 16146
rect 8201 16088 8206 16144
rect 8262 16088 21454 16144
rect 21510 16088 21515 16144
rect 8201 16086 21515 16088
rect 8201 16083 8267 16086
rect 21449 16083 21515 16086
rect 0 16010 800 16040
rect 2037 16010 2103 16013
rect 0 16008 2103 16010
rect 0 15952 2042 16008
rect 2098 15952 2103 16008
rect 0 15950 2103 15952
rect 0 15920 800 15950
rect 2037 15947 2103 15950
rect 3693 16010 3759 16013
rect 6862 16010 6868 16012
rect 3693 16008 6868 16010
rect 3693 15952 3698 16008
rect 3754 15952 6868 16008
rect 3693 15950 6868 15952
rect 3693 15947 3759 15950
rect 6862 15948 6868 15950
rect 6932 15948 6938 16012
rect 16113 16010 16179 16013
rect 18137 16010 18203 16013
rect 16113 16008 18203 16010
rect 16113 15952 16118 16008
rect 16174 15952 18142 16008
rect 18198 15952 18203 16008
rect 16113 15950 18203 15952
rect 16113 15947 16179 15950
rect 18137 15947 18203 15950
rect 21265 16010 21331 16013
rect 22200 16010 23000 16040
rect 21265 16008 23000 16010
rect 21265 15952 21270 16008
rect 21326 15952 23000 16008
rect 21265 15950 23000 15952
rect 21265 15947 21331 15950
rect 22200 15920 23000 15950
rect 6729 15874 6795 15877
rect 7230 15874 7236 15876
rect 6729 15872 7236 15874
rect 6729 15816 6734 15872
rect 6790 15816 7236 15872
rect 6729 15814 7236 15816
rect 6729 15811 6795 15814
rect 7230 15812 7236 15814
rect 7300 15812 7306 15876
rect 14641 15874 14707 15877
rect 14774 15874 14780 15876
rect 14641 15872 14780 15874
rect 14641 15816 14646 15872
rect 14702 15816 14780 15872
rect 14641 15814 14780 15816
rect 14641 15811 14707 15814
rect 14774 15812 14780 15814
rect 14844 15812 14850 15876
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 0 15602 800 15632
rect 1485 15602 1551 15605
rect 0 15600 1551 15602
rect 0 15544 1490 15600
rect 1546 15544 1551 15600
rect 0 15542 1551 15544
rect 0 15512 800 15542
rect 1485 15539 1551 15542
rect 2221 15602 2287 15605
rect 7465 15602 7531 15605
rect 2221 15600 7531 15602
rect 2221 15544 2226 15600
rect 2282 15544 7470 15600
rect 7526 15544 7531 15600
rect 2221 15542 7531 15544
rect 2221 15539 2287 15542
rect 7465 15539 7531 15542
rect 7782 15540 7788 15604
rect 7852 15602 7858 15604
rect 8753 15602 8819 15605
rect 7852 15600 10242 15602
rect 7852 15544 8758 15600
rect 8814 15544 10242 15600
rect 7852 15542 10242 15544
rect 7852 15540 7858 15542
rect 8753 15539 8819 15542
rect 1485 15466 1551 15469
rect 10041 15466 10107 15469
rect 1485 15464 10107 15466
rect 1485 15408 1490 15464
rect 1546 15408 10046 15464
rect 10102 15408 10107 15464
rect 1485 15406 10107 15408
rect 10182 15466 10242 15542
rect 11094 15540 11100 15604
rect 11164 15602 11170 15604
rect 11329 15602 11395 15605
rect 11164 15600 11395 15602
rect 11164 15544 11334 15600
rect 11390 15544 11395 15600
rect 11164 15542 11395 15544
rect 11164 15540 11170 15542
rect 11329 15539 11395 15542
rect 12341 15602 12407 15605
rect 14590 15602 14596 15604
rect 12341 15600 14596 15602
rect 12341 15544 12346 15600
rect 12402 15544 14596 15600
rect 12341 15542 14596 15544
rect 12341 15539 12407 15542
rect 14590 15540 14596 15542
rect 14660 15540 14666 15604
rect 19885 15602 19951 15605
rect 22200 15602 23000 15632
rect 19885 15600 23000 15602
rect 19885 15544 19890 15600
rect 19946 15544 23000 15600
rect 19885 15542 23000 15544
rect 19885 15539 19951 15542
rect 22200 15512 23000 15542
rect 17309 15466 17375 15469
rect 10182 15464 17375 15466
rect 10182 15408 17314 15464
rect 17370 15408 17375 15464
rect 10182 15406 17375 15408
rect 1485 15403 1551 15406
rect 10041 15403 10107 15406
rect 17309 15403 17375 15406
rect 3233 15330 3299 15333
rect 4102 15330 4108 15332
rect 3233 15328 4108 15330
rect 3233 15272 3238 15328
rect 3294 15272 4108 15328
rect 3233 15270 4108 15272
rect 3233 15267 3299 15270
rect 4102 15268 4108 15270
rect 4172 15268 4178 15332
rect 4470 15268 4476 15332
rect 4540 15330 4546 15332
rect 4705 15330 4771 15333
rect 4540 15328 4771 15330
rect 4540 15272 4710 15328
rect 4766 15272 4771 15328
rect 4540 15270 4771 15272
rect 4540 15268 4546 15270
rect 4705 15267 4771 15270
rect 9397 15332 9463 15333
rect 13353 15332 13419 15333
rect 9397 15328 9444 15332
rect 9508 15330 9514 15332
rect 13302 15330 13308 15332
rect 9397 15272 9402 15328
rect 9397 15268 9444 15272
rect 9508 15270 9554 15330
rect 13262 15270 13308 15330
rect 13372 15328 13419 15332
rect 13414 15272 13419 15328
rect 9508 15268 9514 15270
rect 13302 15268 13308 15270
rect 13372 15268 13419 15272
rect 9397 15267 9463 15268
rect 13353 15267 13419 15268
rect 6144 15264 6460 15265
rect 0 15194 800 15224
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 6821 15194 6887 15197
rect 10041 15194 10107 15197
rect 22200 15194 23000 15224
rect 6821 15192 10107 15194
rect 6821 15136 6826 15192
rect 6882 15136 10046 15192
rect 10102 15136 10107 15192
rect 6821 15134 10107 15136
rect 6821 15131 6887 15134
rect 10041 15131 10107 15134
rect 22142 15104 23000 15194
rect 8201 15060 8267 15061
rect 8150 15058 8156 15060
rect 8110 14998 8156 15058
rect 8220 15056 8267 15060
rect 8262 15000 8267 15056
rect 8150 14996 8156 14998
rect 8220 14996 8267 15000
rect 8201 14995 8267 14996
rect 9029 15058 9095 15061
rect 16113 15058 16179 15061
rect 9029 15056 16179 15058
rect 9029 15000 9034 15056
rect 9090 15000 16118 15056
rect 16174 15000 16179 15056
rect 9029 14998 16179 15000
rect 9029 14995 9095 14998
rect 16113 14995 16179 14998
rect 19609 15058 19675 15061
rect 22142 15058 22202 15104
rect 19609 15056 22202 15058
rect 19609 15000 19614 15056
rect 19670 15000 22202 15056
rect 19609 14998 22202 15000
rect 19609 14995 19675 14998
rect 3509 14922 3575 14925
rect 14774 14922 14780 14924
rect 3509 14920 14780 14922
rect 3509 14864 3514 14920
rect 3570 14864 14780 14920
rect 3509 14862 14780 14864
rect 3509 14859 3575 14862
rect 14774 14860 14780 14862
rect 14844 14860 14850 14924
rect 0 14786 800 14816
rect 1485 14786 1551 14789
rect 0 14784 1551 14786
rect 0 14728 1490 14784
rect 1546 14728 1551 14784
rect 0 14726 1551 14728
rect 0 14696 800 14726
rect 1485 14723 1551 14726
rect 6821 14786 6887 14789
rect 8477 14786 8543 14789
rect 6821 14784 8543 14786
rect 6821 14728 6826 14784
rect 6882 14728 8482 14784
rect 8538 14728 8543 14784
rect 6821 14726 8543 14728
rect 6821 14723 6887 14726
rect 8477 14723 8543 14726
rect 10869 14786 10935 14789
rect 12157 14786 12223 14789
rect 12382 14786 12388 14788
rect 10869 14784 12388 14786
rect 10869 14728 10874 14784
rect 10930 14728 12162 14784
rect 12218 14728 12388 14784
rect 10869 14726 12388 14728
rect 10869 14723 10935 14726
rect 12157 14723 12223 14726
rect 12382 14724 12388 14726
rect 12452 14724 12458 14788
rect 20161 14786 20227 14789
rect 22200 14786 23000 14816
rect 20161 14784 23000 14786
rect 20161 14728 20166 14784
rect 20222 14728 23000 14784
rect 20161 14726 23000 14728
rect 20161 14723 20227 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 22200 14696 23000 14726
rect 19139 14655 19455 14656
rect 6085 14650 6151 14653
rect 7465 14650 7531 14653
rect 6085 14648 7531 14650
rect 6085 14592 6090 14648
rect 6146 14592 7470 14648
rect 7526 14592 7531 14648
rect 6085 14590 7531 14592
rect 6085 14587 6151 14590
rect 7465 14587 7531 14590
rect 9630 14590 12450 14650
rect 7097 14514 7163 14517
rect 9630 14514 9690 14590
rect 12390 14517 12450 14590
rect 7097 14512 9690 14514
rect 7097 14456 7102 14512
rect 7158 14456 9690 14512
rect 7097 14454 9690 14456
rect 7097 14451 7163 14454
rect 10174 14452 10180 14516
rect 10244 14514 10250 14516
rect 11053 14514 11119 14517
rect 10244 14512 11119 14514
rect 10244 14456 11058 14512
rect 11114 14456 11119 14512
rect 10244 14454 11119 14456
rect 12390 14514 12499 14517
rect 19006 14514 19012 14516
rect 12390 14512 19012 14514
rect 12390 14456 12438 14512
rect 12494 14456 19012 14512
rect 12390 14454 19012 14456
rect 10244 14452 10250 14454
rect 11053 14451 11119 14454
rect 12433 14451 12499 14454
rect 19006 14452 19012 14454
rect 19076 14452 19082 14516
rect 0 14378 800 14408
rect 2037 14378 2103 14381
rect 0 14376 2103 14378
rect 0 14320 2042 14376
rect 2098 14320 2103 14376
rect 0 14318 2103 14320
rect 0 14288 800 14318
rect 2037 14315 2103 14318
rect 4889 14378 4955 14381
rect 17677 14378 17743 14381
rect 4889 14376 17743 14378
rect 4889 14320 4894 14376
rect 4950 14320 17682 14376
rect 17738 14320 17743 14376
rect 4889 14318 17743 14320
rect 4889 14315 4955 14318
rect 17677 14315 17743 14318
rect 20713 14378 20779 14381
rect 22200 14378 23000 14408
rect 20713 14376 23000 14378
rect 20713 14320 20718 14376
rect 20774 14320 23000 14376
rect 20713 14318 23000 14320
rect 20713 14315 20779 14318
rect 22200 14288 23000 14318
rect 16941 14242 17007 14245
rect 19926 14242 19932 14244
rect 16941 14240 19932 14242
rect 16941 14184 16946 14240
rect 17002 14184 19932 14240
rect 16941 14182 19932 14184
rect 16941 14179 17007 14182
rect 19926 14180 19932 14182
rect 19996 14180 20002 14244
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 8201 14106 8267 14109
rect 8201 14104 9690 14106
rect 8201 14048 8206 14104
rect 8262 14048 9690 14104
rect 8201 14046 9690 14048
rect 8201 14043 8267 14046
rect 0 13970 800 14000
rect 1485 13970 1551 13973
rect 0 13968 1551 13970
rect 0 13912 1490 13968
rect 1546 13912 1551 13968
rect 0 13910 1551 13912
rect 9630 13970 9690 14046
rect 11830 13970 11836 13972
rect 9630 13910 11836 13970
rect 0 13880 800 13910
rect 1485 13907 1551 13910
rect 11830 13908 11836 13910
rect 11900 13908 11906 13972
rect 21357 13970 21423 13973
rect 22200 13970 23000 14000
rect 21357 13968 23000 13970
rect 21357 13912 21362 13968
rect 21418 13912 23000 13968
rect 21357 13910 23000 13912
rect 21357 13907 21423 13910
rect 22200 13880 23000 13910
rect 5441 13834 5507 13837
rect 7557 13836 7623 13837
rect 7414 13834 7420 13836
rect 5441 13832 7420 13834
rect 5441 13776 5446 13832
rect 5502 13776 7420 13832
rect 5441 13774 7420 13776
rect 5441 13771 5507 13774
rect 7414 13772 7420 13774
rect 7484 13772 7490 13836
rect 7557 13832 7604 13836
rect 7668 13834 7674 13836
rect 7557 13776 7562 13832
rect 7557 13772 7604 13776
rect 7668 13774 7714 13834
rect 7790 13774 9690 13834
rect 7668 13772 7674 13774
rect 7557 13771 7623 13772
rect 4061 13698 4127 13701
rect 7790 13698 7850 13774
rect 4061 13696 7850 13698
rect 4061 13640 4066 13696
rect 4122 13640 7850 13696
rect 4061 13638 7850 13640
rect 9630 13698 9690 13774
rect 11697 13698 11763 13701
rect 9630 13696 11763 13698
rect 9630 13640 11702 13696
rect 11758 13640 11763 13696
rect 9630 13638 11763 13640
rect 4061 13635 4127 13638
rect 11697 13635 11763 13638
rect 3545 13632 3861 13633
rect 0 13562 800 13592
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 1485 13562 1551 13565
rect 0 13560 1551 13562
rect 0 13504 1490 13560
rect 1546 13504 1551 13560
rect 0 13502 1551 13504
rect 0 13472 800 13502
rect 1485 13499 1551 13502
rect 6637 13562 6703 13565
rect 7046 13562 7052 13564
rect 6637 13560 7052 13562
rect 6637 13504 6642 13560
rect 6698 13504 7052 13560
rect 6637 13502 7052 13504
rect 6637 13499 6703 13502
rect 7046 13500 7052 13502
rect 7116 13500 7122 13564
rect 21265 13562 21331 13565
rect 22200 13562 23000 13592
rect 21265 13560 23000 13562
rect 21265 13504 21270 13560
rect 21326 13504 23000 13560
rect 21265 13502 23000 13504
rect 21265 13499 21331 13502
rect 22200 13472 23000 13502
rect 2814 13364 2820 13428
rect 2884 13426 2890 13428
rect 5533 13426 5599 13429
rect 2884 13424 5599 13426
rect 2884 13368 5538 13424
rect 5594 13368 5599 13424
rect 2884 13366 5599 13368
rect 2884 13364 2890 13366
rect 5533 13363 5599 13366
rect 6862 13364 6868 13428
rect 6932 13426 6938 13428
rect 9581 13426 9647 13429
rect 6932 13424 9647 13426
rect 6932 13368 9586 13424
rect 9642 13368 9647 13424
rect 6932 13366 9647 13368
rect 6932 13364 6938 13366
rect 9581 13363 9647 13366
rect 3366 13228 3372 13292
rect 3436 13290 3442 13292
rect 8201 13290 8267 13293
rect 3436 13288 8267 13290
rect 3436 13232 8206 13288
rect 8262 13232 8267 13288
rect 3436 13230 8267 13232
rect 3436 13228 3442 13230
rect 8201 13227 8267 13230
rect 19885 13290 19951 13293
rect 19885 13288 22202 13290
rect 19885 13232 19890 13288
rect 19946 13232 22202 13288
rect 19885 13230 22202 13232
rect 19885 13227 19951 13230
rect 22142 13184 22202 13230
rect 0 13154 800 13184
rect 1485 13154 1551 13157
rect 0 13152 1551 13154
rect 0 13096 1490 13152
rect 1546 13096 1551 13152
rect 0 13094 1551 13096
rect 22142 13094 23000 13184
rect 0 13064 800 13094
rect 1485 13091 1551 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 22200 13064 23000 13094
rect 21738 13023 22054 13024
rect 4521 13020 4587 13021
rect 4470 12956 4476 13020
rect 4540 13018 4587 13020
rect 4540 13016 4632 13018
rect 4582 12960 4632 13016
rect 4540 12958 4632 12960
rect 4540 12956 4587 12958
rect 4521 12955 4587 12956
rect 2865 12882 2931 12885
rect 3325 12882 3391 12885
rect 14825 12882 14891 12885
rect 2865 12880 14891 12882
rect 2865 12824 2870 12880
rect 2926 12824 3330 12880
rect 3386 12824 14830 12880
rect 14886 12824 14891 12880
rect 2865 12822 14891 12824
rect 2865 12819 2931 12822
rect 3325 12819 3391 12822
rect 14825 12819 14891 12822
rect 16246 12820 16252 12884
rect 16316 12882 16322 12884
rect 21173 12882 21239 12885
rect 16316 12880 21239 12882
rect 16316 12824 21178 12880
rect 21234 12824 21239 12880
rect 16316 12822 21239 12824
rect 16316 12820 16322 12822
rect 21173 12819 21239 12822
rect 0 12746 800 12776
rect 4061 12746 4127 12749
rect 0 12744 4127 12746
rect 0 12688 4066 12744
rect 4122 12688 4127 12744
rect 0 12686 4127 12688
rect 0 12656 800 12686
rect 4061 12683 4127 12686
rect 4337 12746 4403 12749
rect 15101 12746 15167 12749
rect 4337 12744 15167 12746
rect 4337 12688 4342 12744
rect 4398 12688 15106 12744
rect 15162 12688 15167 12744
rect 4337 12686 15167 12688
rect 4337 12683 4403 12686
rect 15101 12683 15167 12686
rect 15561 12746 15627 12749
rect 18781 12746 18847 12749
rect 15561 12744 18847 12746
rect 15561 12688 15566 12744
rect 15622 12688 18786 12744
rect 18842 12688 18847 12744
rect 15561 12686 18847 12688
rect 15561 12683 15627 12686
rect 18781 12683 18847 12686
rect 21541 12746 21607 12749
rect 22200 12746 23000 12776
rect 21541 12744 23000 12746
rect 21541 12688 21546 12744
rect 21602 12688 23000 12744
rect 21541 12686 23000 12688
rect 21541 12683 21607 12686
rect 22200 12656 23000 12686
rect 3049 12612 3115 12613
rect 2998 12610 3004 12612
rect 2958 12550 3004 12610
rect 3068 12608 3115 12612
rect 3110 12552 3115 12608
rect 2998 12548 3004 12550
rect 3068 12548 3115 12552
rect 3049 12547 3115 12548
rect 4521 12610 4587 12613
rect 6637 12612 6703 12613
rect 6637 12610 6684 12612
rect 4521 12608 4860 12610
rect 4521 12552 4526 12608
rect 4582 12552 4860 12608
rect 4521 12550 4860 12552
rect 6592 12608 6684 12610
rect 6592 12552 6642 12608
rect 6592 12550 6684 12552
rect 4521 12547 4587 12550
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 4800 12477 4860 12550
rect 6637 12548 6684 12550
rect 6748 12548 6754 12612
rect 6821 12608 6887 12613
rect 6821 12552 6826 12608
rect 6882 12552 6887 12608
rect 6637 12547 6703 12548
rect 6821 12547 6887 12552
rect 10726 12548 10732 12612
rect 10796 12610 10802 12612
rect 13721 12610 13787 12613
rect 10796 12608 13787 12610
rect 10796 12552 13726 12608
rect 13782 12552 13787 12608
rect 10796 12550 13787 12552
rect 10796 12548 10802 12550
rect 13721 12547 13787 12550
rect 16481 12610 16547 12613
rect 17309 12610 17375 12613
rect 17769 12610 17835 12613
rect 16481 12608 17835 12610
rect 16481 12552 16486 12608
rect 16542 12552 17314 12608
rect 17370 12552 17774 12608
rect 17830 12552 17835 12608
rect 16481 12550 17835 12552
rect 16481 12547 16547 12550
rect 17309 12547 17375 12550
rect 17769 12547 17835 12550
rect 4797 12472 4863 12477
rect 4797 12416 4802 12472
rect 4858 12416 4863 12472
rect 4797 12411 4863 12416
rect 4981 12474 5047 12477
rect 6824 12474 6884 12547
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 11973 12476 12039 12477
rect 11973 12474 12020 12476
rect 4981 12472 6884 12474
rect 4981 12416 4986 12472
rect 5042 12416 6884 12472
rect 4981 12414 6884 12416
rect 11928 12472 12020 12474
rect 11928 12416 11978 12472
rect 11928 12414 12020 12416
rect 4981 12411 5047 12414
rect 11973 12412 12020 12414
rect 12084 12412 12090 12476
rect 11973 12411 12039 12412
rect 0 12338 800 12368
rect 2773 12338 2839 12341
rect 0 12336 2839 12338
rect 0 12280 2778 12336
rect 2834 12280 2839 12336
rect 0 12278 2839 12280
rect 0 12248 800 12278
rect 2773 12275 2839 12278
rect 7966 12276 7972 12340
rect 8036 12338 8042 12340
rect 8661 12338 8727 12341
rect 8036 12336 8727 12338
rect 8036 12280 8666 12336
rect 8722 12280 8727 12336
rect 8036 12278 8727 12280
rect 8036 12276 8042 12278
rect 8661 12275 8727 12278
rect 12014 12276 12020 12340
rect 12084 12338 12090 12340
rect 12249 12338 12315 12341
rect 12084 12336 12315 12338
rect 12084 12280 12254 12336
rect 12310 12280 12315 12336
rect 12084 12278 12315 12280
rect 12084 12276 12090 12278
rect 12249 12275 12315 12278
rect 14457 12338 14523 12341
rect 18137 12338 18203 12341
rect 14457 12336 18203 12338
rect 14457 12280 14462 12336
rect 14518 12280 18142 12336
rect 18198 12280 18203 12336
rect 14457 12278 18203 12280
rect 14457 12275 14523 12278
rect 18137 12275 18203 12278
rect 20529 12338 20595 12341
rect 22200 12338 23000 12368
rect 20529 12336 23000 12338
rect 20529 12280 20534 12336
rect 20590 12280 23000 12336
rect 20529 12278 23000 12280
rect 20529 12275 20595 12278
rect 22200 12248 23000 12278
rect 4797 12202 4863 12205
rect 18597 12202 18663 12205
rect 4797 12200 18663 12202
rect 4797 12144 4802 12200
rect 4858 12144 18602 12200
rect 18658 12144 18663 12200
rect 4797 12142 18663 12144
rect 4797 12139 4863 12142
rect 18597 12139 18663 12142
rect 6144 12000 6460 12001
rect 0 11930 800 11960
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 2865 11930 2931 11933
rect 0 11928 2931 11930
rect 0 11872 2870 11928
rect 2926 11872 2931 11928
rect 0 11870 2931 11872
rect 0 11840 800 11870
rect 2865 11867 2931 11870
rect 17585 11930 17651 11933
rect 19793 11930 19859 11933
rect 22200 11930 23000 11960
rect 17585 11928 19859 11930
rect 17585 11872 17590 11928
rect 17646 11872 19798 11928
rect 19854 11872 19859 11928
rect 17585 11870 19859 11872
rect 17585 11867 17651 11870
rect 19793 11867 19859 11870
rect 22142 11840 23000 11930
rect 5349 11794 5415 11797
rect 13537 11794 13603 11797
rect 5349 11792 13603 11794
rect 5349 11736 5354 11792
rect 5410 11736 13542 11792
rect 13598 11736 13603 11792
rect 5349 11734 13603 11736
rect 5349 11731 5415 11734
rect 13537 11731 13603 11734
rect 21265 11794 21331 11797
rect 22142 11794 22202 11840
rect 21265 11792 22202 11794
rect 21265 11736 21270 11792
rect 21326 11736 22202 11792
rect 21265 11734 22202 11736
rect 21265 11731 21331 11734
rect 4102 11596 4108 11660
rect 4172 11658 4178 11660
rect 4337 11658 4403 11661
rect 5206 11658 5212 11660
rect 4172 11656 5212 11658
rect 4172 11600 4342 11656
rect 4398 11600 5212 11656
rect 4172 11598 5212 11600
rect 4172 11596 4178 11598
rect 4337 11595 4403 11598
rect 5206 11596 5212 11598
rect 5276 11658 5282 11660
rect 5441 11658 5507 11661
rect 6821 11658 6887 11661
rect 5276 11656 5507 11658
rect 5276 11600 5446 11656
rect 5502 11600 5507 11656
rect 5276 11598 5507 11600
rect 5276 11596 5282 11598
rect 5441 11595 5507 11598
rect 5582 11656 6887 11658
rect 5582 11600 6826 11656
rect 6882 11600 6887 11656
rect 5582 11598 6887 11600
rect 0 11522 800 11552
rect 2221 11522 2287 11525
rect 0 11520 2287 11522
rect 0 11464 2226 11520
rect 2282 11464 2287 11520
rect 0 11462 2287 11464
rect 0 11432 800 11462
rect 2221 11459 2287 11462
rect 4613 11522 4679 11525
rect 5582 11522 5642 11598
rect 6821 11595 6887 11598
rect 4613 11520 5642 11522
rect 4613 11464 4618 11520
rect 4674 11464 5642 11520
rect 4613 11462 5642 11464
rect 5809 11522 5875 11525
rect 5942 11522 5948 11524
rect 5809 11520 5948 11522
rect 5809 11464 5814 11520
rect 5870 11464 5948 11520
rect 5809 11462 5948 11464
rect 4613 11459 4679 11462
rect 5809 11459 5875 11462
rect 5942 11460 5948 11462
rect 6012 11460 6018 11524
rect 21265 11522 21331 11525
rect 22200 11522 23000 11552
rect 21265 11520 23000 11522
rect 21265 11464 21270 11520
rect 21326 11464 23000 11520
rect 21265 11462 23000 11464
rect 21265 11459 21331 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 22200 11432 23000 11462
rect 19139 11391 19455 11392
rect 4470 11188 4476 11252
rect 4540 11250 4546 11252
rect 11145 11250 11211 11253
rect 4540 11248 11211 11250
rect 4540 11192 11150 11248
rect 11206 11192 11211 11248
rect 4540 11190 11211 11192
rect 4540 11188 4546 11190
rect 11145 11187 11211 11190
rect 13353 11250 13419 11253
rect 18086 11250 18092 11252
rect 13353 11248 18092 11250
rect 13353 11192 13358 11248
rect 13414 11192 18092 11248
rect 13353 11190 18092 11192
rect 13353 11187 13419 11190
rect 18086 11188 18092 11190
rect 18156 11188 18162 11252
rect 0 11114 800 11144
rect 3233 11114 3299 11117
rect 0 11112 3299 11114
rect 0 11056 3238 11112
rect 3294 11056 3299 11112
rect 0 11054 3299 11056
rect 0 11024 800 11054
rect 3233 11051 3299 11054
rect 5073 11114 5139 11117
rect 6678 11114 6684 11116
rect 5073 11112 6684 11114
rect 5073 11056 5078 11112
rect 5134 11056 6684 11112
rect 5073 11054 6684 11056
rect 5073 11051 5139 11054
rect 6678 11052 6684 11054
rect 6748 11052 6754 11116
rect 9489 11114 9555 11117
rect 11973 11116 12039 11117
rect 9622 11114 9628 11116
rect 9489 11112 9628 11114
rect 9489 11056 9494 11112
rect 9550 11056 9628 11112
rect 9489 11054 9628 11056
rect 9489 11051 9555 11054
rect 9622 11052 9628 11054
rect 9692 11052 9698 11116
rect 11973 11112 12020 11116
rect 12084 11114 12090 11116
rect 15009 11114 15075 11117
rect 16246 11114 16252 11116
rect 11973 11056 11978 11112
rect 11973 11052 12020 11056
rect 12084 11054 12130 11114
rect 15009 11112 16252 11114
rect 15009 11056 15014 11112
rect 15070 11056 16252 11112
rect 15009 11054 16252 11056
rect 12084 11052 12090 11054
rect 11973 11051 12039 11052
rect 15009 11051 15075 11054
rect 16246 11052 16252 11054
rect 16316 11052 16322 11116
rect 17953 11114 18019 11117
rect 17910 11112 18019 11114
rect 17910 11056 17958 11112
rect 18014 11056 18019 11112
rect 17910 11051 18019 11056
rect 18689 11114 18755 11117
rect 22200 11114 23000 11144
rect 18689 11112 23000 11114
rect 18689 11056 18694 11112
rect 18750 11056 23000 11112
rect 18689 11054 23000 11056
rect 18689 11051 18755 11054
rect 7097 10980 7163 10981
rect 10777 10980 10843 10981
rect 7046 10978 7052 10980
rect 7006 10918 7052 10978
rect 7116 10976 7163 10980
rect 7158 10920 7163 10976
rect 7046 10916 7052 10918
rect 7116 10916 7163 10920
rect 10726 10916 10732 10980
rect 10796 10978 10843 10980
rect 10796 10976 10888 10978
rect 10838 10920 10888 10976
rect 10796 10918 10888 10920
rect 10796 10916 10843 10918
rect 7097 10915 7163 10916
rect 10777 10915 10843 10916
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 11053 10842 11119 10845
rect 12433 10842 12499 10845
rect 6640 10840 11119 10842
rect 6640 10784 11058 10840
rect 11114 10784 11119 10840
rect 6640 10782 11119 10784
rect 0 10706 800 10736
rect 3877 10706 3943 10709
rect 0 10704 3943 10706
rect 0 10648 3882 10704
rect 3938 10648 3943 10704
rect 0 10646 3943 10648
rect 0 10616 800 10646
rect 3877 10643 3943 10646
rect 5073 10706 5139 10709
rect 5993 10706 6059 10709
rect 6640 10706 6700 10782
rect 11053 10779 11119 10782
rect 11792 10840 12499 10842
rect 11792 10784 12438 10840
rect 12494 10784 12499 10840
rect 11792 10782 12499 10784
rect 5073 10704 6700 10706
rect 5073 10648 5078 10704
rect 5134 10648 5998 10704
rect 6054 10648 6700 10704
rect 5073 10646 6700 10648
rect 11145 10706 11211 10709
rect 11792 10706 11852 10782
rect 12433 10779 12499 10782
rect 17910 10706 17970 11051
rect 22200 11024 23000 11054
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 11145 10704 11852 10706
rect 11145 10648 11150 10704
rect 11206 10648 11852 10704
rect 11145 10646 11852 10648
rect 12390 10646 17970 10706
rect 21265 10706 21331 10709
rect 22200 10706 23000 10736
rect 21265 10704 23000 10706
rect 21265 10648 21270 10704
rect 21326 10648 23000 10704
rect 21265 10646 23000 10648
rect 5073 10643 5139 10646
rect 5993 10643 6059 10646
rect 11145 10643 11211 10646
rect 3417 10570 3483 10573
rect 3918 10570 3924 10572
rect 3417 10568 3924 10570
rect 3417 10512 3422 10568
rect 3478 10512 3924 10568
rect 3417 10510 3924 10512
rect 3417 10507 3483 10510
rect 3918 10508 3924 10510
rect 3988 10508 3994 10572
rect 6637 10570 6703 10573
rect 7230 10570 7236 10572
rect 6637 10568 7236 10570
rect 6637 10512 6642 10568
rect 6698 10512 7236 10568
rect 6637 10510 7236 10512
rect 6637 10507 6703 10510
rect 7230 10508 7236 10510
rect 7300 10508 7306 10572
rect 8201 10570 8267 10573
rect 10317 10570 10383 10573
rect 12390 10570 12450 10646
rect 21265 10643 21331 10646
rect 22200 10616 23000 10646
rect 8201 10568 12450 10570
rect 8201 10512 8206 10568
rect 8262 10512 10322 10568
rect 10378 10512 12450 10568
rect 8201 10510 12450 10512
rect 8201 10507 8267 10510
rect 10317 10507 10383 10510
rect 12065 10434 12131 10437
rect 12382 10434 12388 10436
rect 12065 10432 12388 10434
rect 12065 10376 12070 10432
rect 12126 10376 12388 10432
rect 12065 10374 12388 10376
rect 12065 10371 12131 10374
rect 12382 10372 12388 10374
rect 12452 10372 12458 10436
rect 3545 10368 3861 10369
rect 0 10298 800 10328
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 2773 10298 2839 10301
rect 5441 10300 5507 10301
rect 7465 10300 7531 10301
rect 5390 10298 5396 10300
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 5350 10238 5396 10298
rect 5460 10296 5507 10300
rect 5502 10240 5507 10296
rect 0 10208 800 10238
rect 2773 10235 2839 10238
rect 5390 10236 5396 10238
rect 5460 10236 5507 10240
rect 7414 10236 7420 10300
rect 7484 10298 7531 10300
rect 11237 10298 11303 10301
rect 12709 10298 12775 10301
rect 7484 10296 8586 10298
rect 7526 10240 8586 10296
rect 7484 10238 8586 10240
rect 7484 10236 7531 10238
rect 5441 10235 5507 10236
rect 7465 10235 7531 10236
rect 3509 10162 3575 10165
rect 7097 10162 7163 10165
rect 3509 10160 7163 10162
rect 3509 10104 3514 10160
rect 3570 10104 7102 10160
rect 7158 10104 7163 10160
rect 3509 10102 7163 10104
rect 3509 10099 3575 10102
rect 7097 10099 7163 10102
rect 2078 9964 2084 10028
rect 2148 10026 2154 10028
rect 7465 10026 7531 10029
rect 2148 10024 7531 10026
rect 2148 9968 7470 10024
rect 7526 9968 7531 10024
rect 2148 9966 7531 9968
rect 8526 10026 8586 10238
rect 11237 10296 12775 10298
rect 11237 10240 11242 10296
rect 11298 10240 12714 10296
rect 12770 10240 12775 10296
rect 11237 10238 12775 10240
rect 11237 10235 11303 10238
rect 12709 10235 12775 10238
rect 20161 10298 20227 10301
rect 22200 10298 23000 10328
rect 20161 10296 23000 10298
rect 20161 10240 20166 10296
rect 20222 10240 23000 10296
rect 20161 10238 23000 10240
rect 20161 10235 20227 10238
rect 22200 10208 23000 10238
rect 8661 10162 8727 10165
rect 19977 10162 20043 10165
rect 8661 10160 20043 10162
rect 8661 10104 8666 10160
rect 8722 10104 19982 10160
rect 20038 10104 20043 10160
rect 8661 10102 20043 10104
rect 8661 10099 8727 10102
rect 19977 10099 20043 10102
rect 12893 10026 12959 10029
rect 8526 10024 12959 10026
rect 8526 9968 12898 10024
rect 12954 9968 12959 10024
rect 8526 9966 12959 9968
rect 2148 9964 2154 9966
rect 7465 9963 7531 9966
rect 12893 9963 12959 9966
rect 13445 10026 13511 10029
rect 16941 10026 17007 10029
rect 13445 10024 17007 10026
rect 13445 9968 13450 10024
rect 13506 9968 16946 10024
rect 17002 9968 17007 10024
rect 13445 9966 17007 9968
rect 13445 9963 13511 9966
rect 16941 9963 17007 9966
rect 20529 10026 20595 10029
rect 20529 10024 22202 10026
rect 20529 9968 20534 10024
rect 20590 9968 22202 10024
rect 20529 9966 22202 9968
rect 20529 9963 20595 9966
rect 22142 9920 22202 9966
rect 0 9890 800 9920
rect 2773 9890 2839 9893
rect 0 9888 2839 9890
rect 0 9832 2778 9888
rect 2834 9832 2839 9888
rect 0 9830 2839 9832
rect 22142 9830 23000 9920
rect 0 9800 800 9830
rect 2773 9827 2839 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 22200 9800 23000 9830
rect 21738 9759 22054 9760
rect 4889 9618 4955 9621
rect 12249 9618 12315 9621
rect 20437 9618 20503 9621
rect 4889 9616 20503 9618
rect 4889 9560 4894 9616
rect 4950 9560 12254 9616
rect 12310 9560 20442 9616
rect 20498 9560 20503 9616
rect 4889 9558 20503 9560
rect 4889 9555 4955 9558
rect 12249 9555 12315 9558
rect 20437 9555 20503 9558
rect 0 9482 800 9512
rect 3233 9482 3299 9485
rect 3693 9482 3759 9485
rect 0 9480 3759 9482
rect 0 9424 3238 9480
rect 3294 9424 3698 9480
rect 3754 9424 3759 9480
rect 0 9422 3759 9424
rect 0 9392 800 9422
rect 3233 9419 3299 9422
rect 3693 9419 3759 9422
rect 19057 9482 19123 9485
rect 22200 9482 23000 9512
rect 19057 9480 23000 9482
rect 19057 9424 19062 9480
rect 19118 9424 23000 9480
rect 19057 9422 23000 9424
rect 19057 9419 19123 9422
rect 22200 9392 23000 9422
rect 15561 9346 15627 9349
rect 17953 9346 18019 9349
rect 15561 9344 18019 9346
rect 15561 9288 15566 9344
rect 15622 9288 17958 9344
rect 18014 9288 18019 9344
rect 15561 9286 18019 9288
rect 15561 9283 15627 9286
rect 17953 9283 18019 9286
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 4429 9210 4495 9213
rect 5942 9210 5948 9212
rect 4429 9208 4538 9210
rect 4429 9152 4434 9208
rect 4490 9152 4538 9208
rect 4429 9147 4538 9152
rect 0 9074 800 9104
rect 3877 9074 3943 9077
rect 0 9072 3943 9074
rect 0 9016 3882 9072
rect 3938 9016 3943 9072
rect 0 9014 3943 9016
rect 4478 9074 4538 9147
rect 5766 9150 5948 9210
rect 5766 9077 5826 9150
rect 5942 9148 5948 9150
rect 6012 9148 6018 9212
rect 17401 9210 17467 9213
rect 17861 9210 17927 9213
rect 20897 9210 20963 9213
rect 17401 9208 17927 9210
rect 17401 9152 17406 9208
rect 17462 9152 17866 9208
rect 17922 9152 17927 9208
rect 17401 9150 17927 9152
rect 17401 9147 17467 9150
rect 17861 9147 17927 9150
rect 20302 9208 20963 9210
rect 20302 9152 20902 9208
rect 20958 9152 20963 9208
rect 20302 9150 20963 9152
rect 5717 9074 5826 9077
rect 4478 9072 5826 9074
rect 4478 9016 5722 9072
rect 5778 9016 5826 9072
rect 4478 9014 5826 9016
rect 5993 9074 6059 9077
rect 20302 9074 20362 9150
rect 20897 9147 20963 9150
rect 5993 9072 20362 9074
rect 5993 9016 5998 9072
rect 6054 9016 20362 9072
rect 5993 9014 20362 9016
rect 20529 9074 20595 9077
rect 22200 9074 23000 9104
rect 20529 9072 23000 9074
rect 20529 9016 20534 9072
rect 20590 9016 23000 9072
rect 20529 9014 23000 9016
rect 0 8984 800 9014
rect 3877 9011 3943 9014
rect 5717 9011 5783 9014
rect 5993 9011 6059 9014
rect 20529 9011 20595 9014
rect 22200 8984 23000 9014
rect 11830 8876 11836 8940
rect 11900 8938 11906 8940
rect 21081 8938 21147 8941
rect 11900 8936 21147 8938
rect 11900 8880 21086 8936
rect 21142 8880 21147 8936
rect 11900 8878 21147 8880
rect 11900 8876 11906 8878
rect 21081 8875 21147 8878
rect 21265 8938 21331 8941
rect 21265 8936 22018 8938
rect 21265 8880 21270 8936
rect 21326 8904 22018 8936
rect 21326 8880 22202 8904
rect 21265 8878 22202 8880
rect 21265 8875 21331 8878
rect 21958 8844 22202 8878
rect 6144 8736 6460 8737
rect 0 8666 800 8696
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 22142 8696 22202 8844
rect 2221 8666 2287 8669
rect 0 8664 2287 8666
rect 0 8608 2226 8664
rect 2282 8608 2287 8664
rect 0 8606 2287 8608
rect 0 8576 800 8606
rect 2221 8603 2287 8606
rect 8753 8666 8819 8669
rect 9489 8666 9555 8669
rect 8753 8664 9555 8666
rect 8753 8608 8758 8664
rect 8814 8608 9494 8664
rect 9550 8608 9555 8664
rect 8753 8606 9555 8608
rect 22142 8606 23000 8696
rect 8753 8603 8819 8606
rect 9489 8603 9555 8606
rect 22200 8576 23000 8606
rect 4153 8530 4219 8533
rect 4286 8530 4292 8532
rect 4153 8528 4292 8530
rect 4153 8472 4158 8528
rect 4214 8472 4292 8528
rect 4153 8470 4292 8472
rect 4153 8467 4219 8470
rect 4286 8468 4292 8470
rect 4356 8468 4362 8532
rect 6821 8530 6887 8533
rect 8201 8530 8267 8533
rect 20805 8530 20871 8533
rect 6821 8528 7298 8530
rect 6821 8472 6826 8528
rect 6882 8472 7298 8528
rect 6821 8470 7298 8472
rect 6821 8467 6887 8470
rect 4245 8394 4311 8397
rect 5390 8394 5396 8396
rect 4245 8392 5396 8394
rect 4245 8336 4250 8392
rect 4306 8336 5396 8392
rect 4245 8334 5396 8336
rect 4245 8331 4311 8334
rect 5390 8332 5396 8334
rect 5460 8332 5466 8396
rect 5809 8394 5875 8397
rect 7097 8394 7163 8397
rect 5809 8392 7163 8394
rect 5809 8336 5814 8392
rect 5870 8336 7102 8392
rect 7158 8336 7163 8392
rect 5809 8334 7163 8336
rect 7238 8394 7298 8470
rect 8201 8528 20871 8530
rect 8201 8472 8206 8528
rect 8262 8472 20810 8528
rect 20866 8472 20871 8528
rect 8201 8470 20871 8472
rect 8201 8467 8267 8470
rect 20805 8467 20871 8470
rect 9489 8394 9555 8397
rect 7238 8392 9555 8394
rect 7238 8336 9494 8392
rect 9550 8336 9555 8392
rect 7238 8334 9555 8336
rect 5809 8331 5875 8334
rect 7097 8331 7163 8334
rect 9489 8331 9555 8334
rect 0 8258 800 8288
rect 1945 8258 2011 8261
rect 2221 8258 2287 8261
rect 0 8256 2287 8258
rect 0 8200 1950 8256
rect 2006 8200 2226 8256
rect 2282 8200 2287 8256
rect 0 8198 2287 8200
rect 0 8168 800 8198
rect 1945 8195 2011 8198
rect 2221 8195 2287 8198
rect 9673 8258 9739 8261
rect 10133 8258 10199 8261
rect 9673 8256 10199 8258
rect 9673 8200 9678 8256
rect 9734 8200 10138 8256
rect 10194 8200 10199 8256
rect 9673 8198 10199 8200
rect 9673 8195 9739 8198
rect 10133 8195 10199 8198
rect 21265 8258 21331 8261
rect 22200 8258 23000 8288
rect 21265 8256 23000 8258
rect 21265 8200 21270 8256
rect 21326 8200 23000 8256
rect 21265 8198 23000 8200
rect 21265 8195 21331 8198
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 22200 8168 23000 8198
rect 19139 8127 19455 8128
rect 13118 8122 13124 8124
rect 9262 8062 13124 8122
rect 2313 7986 2379 7989
rect 9262 7986 9322 8062
rect 13118 8060 13124 8062
rect 13188 8060 13194 8124
rect 2313 7984 9322 7986
rect 2313 7928 2318 7984
rect 2374 7928 9322 7984
rect 2313 7926 9322 7928
rect 2313 7923 2379 7926
rect 12198 7924 12204 7988
rect 12268 7986 12274 7988
rect 12801 7986 12867 7989
rect 12268 7984 12867 7986
rect 12268 7928 12806 7984
rect 12862 7928 12867 7984
rect 12268 7926 12867 7928
rect 12268 7924 12274 7926
rect 12801 7923 12867 7926
rect 0 7850 800 7880
rect 3969 7850 4035 7853
rect 6729 7850 6795 7853
rect 0 7848 4035 7850
rect 0 7792 3974 7848
rect 4030 7792 4035 7848
rect 0 7790 4035 7792
rect 0 7760 800 7790
rect 3969 7787 4035 7790
rect 5950 7848 6795 7850
rect 5950 7792 6734 7848
rect 6790 7792 6795 7848
rect 5950 7790 6795 7792
rect 5257 7714 5323 7717
rect 5950 7714 6010 7790
rect 6729 7787 6795 7790
rect 9949 7850 10015 7853
rect 12985 7850 13051 7853
rect 9949 7848 13051 7850
rect 9949 7792 9954 7848
rect 10010 7792 12990 7848
rect 13046 7792 13051 7848
rect 9949 7790 13051 7792
rect 9949 7787 10015 7790
rect 12985 7787 13051 7790
rect 18689 7850 18755 7853
rect 22200 7850 23000 7880
rect 18689 7848 23000 7850
rect 18689 7792 18694 7848
rect 18750 7792 23000 7848
rect 18689 7790 23000 7792
rect 18689 7787 18755 7790
rect 22200 7760 23000 7790
rect 5257 7712 6010 7714
rect 5257 7656 5262 7712
rect 5318 7656 6010 7712
rect 5257 7654 6010 7656
rect 5257 7651 5323 7654
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 8334 7516 8340 7580
rect 8404 7578 8410 7580
rect 8569 7578 8635 7581
rect 8404 7576 8635 7578
rect 8404 7520 8574 7576
rect 8630 7520 8635 7576
rect 8404 7518 8635 7520
rect 8404 7516 8410 7518
rect 8569 7515 8635 7518
rect 0 7442 800 7472
rect 2865 7442 2931 7445
rect 3325 7444 3391 7445
rect 3325 7442 3372 7444
rect 0 7440 2931 7442
rect 0 7384 2870 7440
rect 2926 7384 2931 7440
rect 0 7382 2931 7384
rect 3280 7440 3372 7442
rect 3280 7384 3330 7440
rect 3280 7382 3372 7384
rect 0 7352 800 7382
rect 2865 7379 2931 7382
rect 3325 7380 3372 7382
rect 3436 7380 3442 7444
rect 13629 7442 13695 7445
rect 18413 7442 18479 7445
rect 5214 7382 12450 7442
rect 3325 7379 3391 7380
rect 2313 7306 2379 7309
rect 3141 7306 3207 7309
rect 5214 7306 5274 7382
rect 2313 7304 5274 7306
rect 2313 7248 2318 7304
rect 2374 7248 3146 7304
rect 3202 7248 5274 7304
rect 2313 7246 5274 7248
rect 8201 7306 8267 7309
rect 11053 7306 11119 7309
rect 8201 7304 11119 7306
rect 8201 7248 8206 7304
rect 8262 7248 11058 7304
rect 11114 7248 11119 7304
rect 8201 7246 11119 7248
rect 12390 7306 12450 7382
rect 13629 7440 18479 7442
rect 13629 7384 13634 7440
rect 13690 7384 18418 7440
rect 18474 7384 18479 7440
rect 13629 7382 18479 7384
rect 13629 7379 13695 7382
rect 18413 7379 18479 7382
rect 20529 7442 20595 7445
rect 22200 7442 23000 7472
rect 20529 7440 23000 7442
rect 20529 7384 20534 7440
rect 20590 7384 23000 7440
rect 20529 7382 23000 7384
rect 20529 7379 20595 7382
rect 22200 7352 23000 7382
rect 12617 7306 12683 7309
rect 12390 7304 12683 7306
rect 12390 7248 12622 7304
rect 12678 7248 12683 7304
rect 12390 7246 12683 7248
rect 2313 7243 2379 7246
rect 3141 7243 3207 7246
rect 8201 7243 8267 7246
rect 11053 7243 11119 7246
rect 12617 7243 12683 7246
rect 15009 7306 15075 7309
rect 15009 7304 19626 7306
rect 15009 7248 15014 7304
rect 15070 7248 19626 7304
rect 15009 7246 19626 7248
rect 15009 7243 15075 7246
rect 9305 7172 9371 7173
rect 9254 7108 9260 7172
rect 9324 7170 9371 7172
rect 14457 7170 14523 7173
rect 18965 7170 19031 7173
rect 9324 7168 9416 7170
rect 9366 7112 9416 7168
rect 9324 7110 9416 7112
rect 14457 7168 19031 7170
rect 14457 7112 14462 7168
rect 14518 7112 18970 7168
rect 19026 7112 19031 7168
rect 14457 7110 19031 7112
rect 9324 7108 9371 7110
rect 9305 7107 9371 7108
rect 14457 7107 14523 7110
rect 18965 7107 19031 7110
rect 3545 7104 3861 7105
rect 0 7034 800 7064
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 2681 7034 2747 7037
rect 0 7032 2747 7034
rect 0 6976 2686 7032
rect 2742 6976 2747 7032
rect 0 6974 2747 6976
rect 0 6944 800 6974
rect 2681 6971 2747 6974
rect 5349 7034 5415 7037
rect 9949 7034 10015 7037
rect 5349 7032 8586 7034
rect 5349 6976 5354 7032
rect 5410 6976 8586 7032
rect 5349 6974 8586 6976
rect 5349 6971 5415 6974
rect 5717 6898 5783 6901
rect 7741 6898 7807 6901
rect 5717 6896 7807 6898
rect 5717 6840 5722 6896
rect 5778 6840 7746 6896
rect 7802 6840 7807 6896
rect 5717 6838 7807 6840
rect 8526 6898 8586 6974
rect 9262 7032 10015 7034
rect 9262 6976 9954 7032
rect 10010 6976 10015 7032
rect 9262 6974 10015 6976
rect 9262 6898 9322 6974
rect 9949 6971 10015 6974
rect 15193 7034 15259 7037
rect 18505 7034 18571 7037
rect 15193 7032 18571 7034
rect 15193 6976 15198 7032
rect 15254 6976 18510 7032
rect 18566 6976 18571 7032
rect 15193 6974 18571 6976
rect 19566 7034 19626 7246
rect 21357 7034 21423 7037
rect 22200 7034 23000 7064
rect 19566 7032 23000 7034
rect 19566 6976 21362 7032
rect 21418 6976 23000 7032
rect 19566 6974 23000 6976
rect 15193 6971 15259 6974
rect 18505 6971 18571 6974
rect 21357 6971 21423 6974
rect 22200 6944 23000 6974
rect 8526 6838 9322 6898
rect 9489 6898 9555 6901
rect 19977 6898 20043 6901
rect 9489 6896 20043 6898
rect 9489 6840 9494 6896
rect 9550 6840 19982 6896
rect 20038 6840 20043 6896
rect 9489 6838 20043 6840
rect 5717 6835 5783 6838
rect 7741 6835 7807 6838
rect 9489 6835 9555 6838
rect 19977 6835 20043 6838
rect 2630 6700 2636 6764
rect 2700 6762 2706 6764
rect 3785 6762 3851 6765
rect 12525 6762 12591 6765
rect 2700 6760 3851 6762
rect 2700 6704 3790 6760
rect 3846 6704 3851 6760
rect 2700 6702 3851 6704
rect 2700 6700 2706 6702
rect 3785 6699 3851 6702
rect 5950 6760 12591 6762
rect 5950 6704 12530 6760
rect 12586 6704 12591 6760
rect 5950 6702 12591 6704
rect 0 6626 800 6656
rect 1485 6626 1551 6629
rect 5950 6626 6010 6702
rect 12525 6699 12591 6702
rect 14825 6762 14891 6765
rect 15142 6762 15148 6764
rect 14825 6760 15148 6762
rect 14825 6704 14830 6760
rect 14886 6704 15148 6760
rect 14825 6702 15148 6704
rect 14825 6699 14891 6702
rect 15142 6700 15148 6702
rect 15212 6700 15218 6764
rect 16573 6762 16639 6765
rect 16982 6762 16988 6764
rect 16573 6760 16988 6762
rect 16573 6704 16578 6760
rect 16634 6704 16988 6760
rect 16573 6702 16988 6704
rect 16573 6699 16639 6702
rect 16982 6700 16988 6702
rect 17052 6700 17058 6764
rect 19006 6700 19012 6764
rect 19076 6762 19082 6764
rect 19241 6762 19307 6765
rect 19076 6760 19307 6762
rect 19076 6704 19246 6760
rect 19302 6704 19307 6760
rect 19076 6702 19307 6704
rect 19076 6700 19082 6702
rect 19241 6699 19307 6702
rect 20713 6762 20779 6765
rect 20713 6760 22202 6762
rect 20713 6704 20718 6760
rect 20774 6704 22202 6760
rect 20713 6702 22202 6704
rect 20713 6699 20779 6702
rect 22142 6656 22202 6702
rect 0 6624 6010 6626
rect 0 6568 1490 6624
rect 1546 6568 6010 6624
rect 0 6566 6010 6568
rect 16941 6628 17007 6629
rect 16941 6624 16988 6628
rect 17052 6626 17058 6628
rect 16941 6568 16946 6624
rect 0 6536 800 6566
rect 1485 6563 1551 6566
rect 16941 6564 16988 6568
rect 17052 6566 17098 6626
rect 22142 6566 23000 6656
rect 17052 6564 17058 6566
rect 16941 6563 17007 6564
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 22200 6536 23000 6566
rect 21738 6495 22054 6496
rect 6862 6428 6868 6492
rect 6932 6490 6938 6492
rect 7557 6490 7623 6493
rect 8109 6490 8175 6493
rect 6932 6488 7623 6490
rect 6932 6432 7562 6488
rect 7618 6432 7623 6488
rect 6932 6430 7623 6432
rect 6932 6428 6938 6430
rect 7557 6427 7623 6430
rect 7790 6488 8175 6490
rect 7790 6432 8114 6488
rect 8170 6432 8175 6488
rect 7790 6430 8175 6432
rect 1577 6354 1643 6357
rect 2078 6354 2084 6356
rect 1577 6352 2084 6354
rect 1577 6296 1582 6352
rect 1638 6296 2084 6352
rect 1577 6294 2084 6296
rect 1577 6291 1643 6294
rect 2078 6292 2084 6294
rect 2148 6292 2154 6356
rect 6361 6354 6427 6357
rect 7790 6354 7850 6430
rect 8109 6427 8175 6430
rect 18045 6490 18111 6493
rect 18229 6490 18295 6493
rect 18045 6488 18295 6490
rect 18045 6432 18050 6488
rect 18106 6432 18234 6488
rect 18290 6432 18295 6488
rect 18045 6430 18295 6432
rect 18045 6427 18111 6430
rect 18229 6427 18295 6430
rect 6361 6352 7850 6354
rect 6361 6296 6366 6352
rect 6422 6296 7850 6352
rect 6361 6294 7850 6296
rect 8109 6354 8175 6357
rect 15285 6354 15351 6357
rect 19241 6354 19307 6357
rect 8109 6352 19307 6354
rect 8109 6296 8114 6352
rect 8170 6296 15290 6352
rect 15346 6296 19246 6352
rect 19302 6296 19307 6352
rect 8109 6294 19307 6296
rect 6361 6291 6427 6294
rect 8109 6291 8175 6294
rect 15285 6291 15351 6294
rect 19241 6291 19307 6294
rect 19609 6354 19675 6357
rect 20805 6354 20871 6357
rect 21081 6354 21147 6357
rect 19609 6352 21147 6354
rect 19609 6296 19614 6352
rect 19670 6296 20810 6352
rect 20866 6296 21086 6352
rect 21142 6296 21147 6352
rect 19609 6294 21147 6296
rect 19609 6291 19675 6294
rect 20805 6291 20871 6294
rect 21081 6291 21147 6294
rect 0 6218 800 6248
rect 2814 6218 2820 6220
rect 0 6158 2820 6218
rect 0 6128 800 6158
rect 2814 6156 2820 6158
rect 2884 6218 2890 6220
rect 3417 6218 3483 6221
rect 2884 6216 3483 6218
rect 2884 6160 3422 6216
rect 3478 6160 3483 6216
rect 2884 6158 3483 6160
rect 2884 6156 2890 6158
rect 3417 6155 3483 6158
rect 5165 6218 5231 6221
rect 17677 6218 17743 6221
rect 5165 6216 17743 6218
rect 5165 6160 5170 6216
rect 5226 6160 17682 6216
rect 17738 6160 17743 6216
rect 5165 6158 17743 6160
rect 5165 6155 5231 6158
rect 17677 6155 17743 6158
rect 18505 6218 18571 6221
rect 22200 6218 23000 6248
rect 18505 6216 23000 6218
rect 18505 6160 18510 6216
rect 18566 6160 23000 6216
rect 18505 6158 23000 6160
rect 18505 6155 18571 6158
rect 22200 6128 23000 6158
rect 15561 6082 15627 6085
rect 17953 6082 18019 6085
rect 15561 6080 18019 6082
rect 15561 6024 15566 6080
rect 15622 6024 17958 6080
rect 18014 6024 18019 6080
rect 15561 6022 18019 6024
rect 15561 6019 15627 6022
rect 17953 6019 18019 6022
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 4337 5946 4403 5949
rect 4470 5946 4476 5948
rect 4337 5944 4476 5946
rect 4337 5888 4342 5944
rect 4398 5888 4476 5944
rect 4337 5886 4476 5888
rect 4337 5883 4403 5886
rect 4470 5884 4476 5886
rect 4540 5884 4546 5948
rect 4613 5946 4679 5949
rect 7005 5946 7071 5949
rect 4613 5944 7071 5946
rect 4613 5888 4618 5944
rect 4674 5888 7010 5944
rect 7066 5888 7071 5944
rect 4613 5886 7071 5888
rect 4613 5883 4679 5886
rect 7005 5883 7071 5886
rect 9305 5946 9371 5949
rect 11697 5946 11763 5949
rect 9305 5944 11763 5946
rect 9305 5888 9310 5944
rect 9366 5888 11702 5944
rect 11758 5888 11763 5944
rect 9305 5886 11763 5888
rect 9305 5883 9371 5886
rect 11697 5883 11763 5886
rect 15285 5946 15351 5949
rect 18822 5946 18828 5948
rect 15285 5944 18828 5946
rect 15285 5888 15290 5944
rect 15346 5888 18828 5944
rect 15285 5886 18828 5888
rect 15285 5883 15351 5886
rect 18822 5884 18828 5886
rect 18892 5884 18898 5948
rect 0 5810 800 5840
rect 933 5810 999 5813
rect 0 5808 999 5810
rect 0 5752 938 5808
rect 994 5752 999 5808
rect 0 5750 999 5752
rect 0 5720 800 5750
rect 933 5747 999 5750
rect 1853 5810 1919 5813
rect 12157 5810 12223 5813
rect 1853 5808 12223 5810
rect 1853 5752 1858 5808
rect 1914 5752 12162 5808
rect 12218 5752 12223 5808
rect 1853 5750 12223 5752
rect 1853 5747 1919 5750
rect 12157 5747 12223 5750
rect 16849 5810 16915 5813
rect 18321 5810 18387 5813
rect 16849 5808 18387 5810
rect 16849 5752 16854 5808
rect 16910 5752 18326 5808
rect 18382 5752 18387 5808
rect 16849 5750 18387 5752
rect 16849 5747 16915 5750
rect 18321 5747 18387 5750
rect 18873 5810 18939 5813
rect 22200 5810 23000 5840
rect 18873 5808 23000 5810
rect 18873 5752 18878 5808
rect 18934 5752 23000 5808
rect 18873 5750 23000 5752
rect 18873 5747 18939 5750
rect 22200 5720 23000 5750
rect 1669 5674 1735 5677
rect 2998 5674 3004 5676
rect 1669 5672 3004 5674
rect 1669 5616 1674 5672
rect 1730 5616 3004 5672
rect 1669 5614 3004 5616
rect 1669 5611 1735 5614
rect 2998 5612 3004 5614
rect 3068 5612 3074 5676
rect 3969 5674 4035 5677
rect 6361 5674 6427 5677
rect 6729 5676 6795 5677
rect 3969 5672 6427 5674
rect 3969 5616 3974 5672
rect 4030 5616 6366 5672
rect 6422 5616 6427 5672
rect 3969 5614 6427 5616
rect 3969 5611 4035 5614
rect 6361 5611 6427 5614
rect 6678 5612 6684 5676
rect 6748 5674 6795 5676
rect 16113 5674 16179 5677
rect 19609 5674 19675 5677
rect 6748 5672 6840 5674
rect 6790 5616 6840 5672
rect 6748 5614 6840 5616
rect 16113 5672 19675 5674
rect 16113 5616 16118 5672
rect 16174 5616 19614 5672
rect 19670 5616 19675 5672
rect 16113 5614 19675 5616
rect 6748 5612 6795 5614
rect 6729 5611 6795 5612
rect 16113 5611 16179 5614
rect 19609 5611 19675 5614
rect 4153 5538 4219 5541
rect 5901 5538 5967 5541
rect 4153 5536 5967 5538
rect 4153 5480 4158 5536
rect 4214 5480 5906 5536
rect 5962 5480 5967 5536
rect 4153 5478 5967 5480
rect 4153 5475 4219 5478
rect 5901 5475 5967 5478
rect 19006 5476 19012 5540
rect 19076 5538 19082 5540
rect 19149 5538 19215 5541
rect 19076 5536 19215 5538
rect 19076 5480 19154 5536
rect 19210 5480 19215 5536
rect 19076 5478 19215 5480
rect 19076 5476 19082 5478
rect 19149 5475 19215 5478
rect 6144 5472 6460 5473
rect 0 5402 800 5432
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 17585 5402 17651 5405
rect 18137 5404 18203 5405
rect 17718 5402 17724 5404
rect 0 5342 2790 5402
rect 0 5312 800 5342
rect 2730 5266 2790 5342
rect 17585 5400 17724 5402
rect 17585 5344 17590 5400
rect 17646 5344 17724 5400
rect 17585 5342 17724 5344
rect 17585 5339 17651 5342
rect 17718 5340 17724 5342
rect 17788 5340 17794 5404
rect 18086 5340 18092 5404
rect 18156 5402 18203 5404
rect 21541 5402 21607 5405
rect 22200 5402 23000 5432
rect 18156 5400 18248 5402
rect 18198 5344 18248 5400
rect 18156 5342 18248 5344
rect 18646 5400 21607 5402
rect 18646 5344 21546 5400
rect 21602 5344 21607 5400
rect 18646 5342 21607 5344
rect 18156 5340 18203 5342
rect 18137 5339 18203 5340
rect 3325 5266 3391 5269
rect 10174 5266 10180 5268
rect 2730 5264 10180 5266
rect 2730 5208 3330 5264
rect 3386 5208 10180 5264
rect 2730 5206 10180 5208
rect 3325 5203 3391 5206
rect 10174 5204 10180 5206
rect 10244 5204 10250 5268
rect 14457 5266 14523 5269
rect 18646 5266 18706 5342
rect 21541 5339 21607 5342
rect 22142 5312 23000 5402
rect 14457 5264 18706 5266
rect 14457 5208 14462 5264
rect 14518 5208 18706 5264
rect 14457 5206 18706 5208
rect 18873 5266 18939 5269
rect 22142 5266 22202 5312
rect 18873 5264 22202 5266
rect 18873 5208 18878 5264
rect 18934 5208 22202 5264
rect 18873 5206 22202 5208
rect 14457 5203 14523 5206
rect 18873 5203 18939 5206
rect 5390 5068 5396 5132
rect 5460 5130 5466 5132
rect 21081 5130 21147 5133
rect 5460 5128 21147 5130
rect 5460 5072 21086 5128
rect 21142 5072 21147 5128
rect 5460 5070 21147 5072
rect 5460 5068 5466 5070
rect 21081 5067 21147 5070
rect 0 4994 800 5024
rect 933 4994 999 4997
rect 3417 4994 3483 4997
rect 0 4992 3483 4994
rect 0 4936 938 4992
rect 994 4936 3422 4992
rect 3478 4936 3483 4992
rect 0 4934 3483 4936
rect 0 4904 800 4934
rect 933 4931 999 4934
rect 3417 4931 3483 4934
rect 14917 4994 14983 4997
rect 18045 4994 18111 4997
rect 14917 4992 18111 4994
rect 14917 4936 14922 4992
rect 14978 4936 18050 4992
rect 18106 4936 18111 4992
rect 14917 4934 18111 4936
rect 14917 4931 14983 4934
rect 18045 4931 18111 4934
rect 19885 4994 19951 4997
rect 22200 4994 23000 5024
rect 19885 4992 23000 4994
rect 19885 4936 19890 4992
rect 19946 4936 23000 4992
rect 19885 4934 23000 4936
rect 19885 4931 19951 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 22200 4904 23000 4934
rect 19139 4863 19455 4864
rect 9806 4796 9812 4860
rect 9876 4858 9882 4860
rect 12014 4858 12020 4860
rect 9876 4798 12020 4858
rect 9876 4796 9882 4798
rect 12014 4796 12020 4798
rect 12084 4796 12090 4860
rect 3049 4722 3115 4725
rect 6453 4722 6519 4725
rect 16113 4722 16179 4725
rect 3049 4720 16179 4722
rect 3049 4664 3054 4720
rect 3110 4664 6458 4720
rect 6514 4664 16118 4720
rect 16174 4664 16179 4720
rect 3049 4662 16179 4664
rect 3049 4659 3115 4662
rect 6453 4659 6519 4662
rect 16113 4659 16179 4662
rect 16941 4722 17007 4725
rect 17493 4722 17559 4725
rect 16941 4720 17559 4722
rect 16941 4664 16946 4720
rect 17002 4664 17498 4720
rect 17554 4664 17559 4720
rect 16941 4662 17559 4664
rect 16941 4659 17007 4662
rect 17493 4659 17559 4662
rect 18137 4722 18203 4725
rect 18137 4720 21098 4722
rect 18137 4664 18142 4720
rect 18198 4664 21098 4720
rect 18137 4662 21098 4664
rect 18137 4659 18203 4662
rect 0 4586 800 4616
rect 2221 4586 2287 4589
rect 0 4584 2287 4586
rect 0 4528 2226 4584
rect 2282 4528 2287 4584
rect 0 4526 2287 4528
rect 0 4496 800 4526
rect 2221 4523 2287 4526
rect 2773 4586 2839 4589
rect 15285 4586 15351 4589
rect 2773 4584 15351 4586
rect 2773 4528 2778 4584
rect 2834 4528 15290 4584
rect 15346 4528 15351 4584
rect 2773 4526 15351 4528
rect 2773 4523 2839 4526
rect 15285 4523 15351 4526
rect 16297 4586 16363 4589
rect 21038 4586 21098 4662
rect 22200 4586 23000 4616
rect 16297 4584 20914 4586
rect 16297 4528 16302 4584
rect 16358 4528 20914 4584
rect 16297 4526 20914 4528
rect 21038 4526 23000 4586
rect 16297 4523 16363 4526
rect 4286 4388 4292 4452
rect 4356 4450 4362 4452
rect 4613 4450 4679 4453
rect 4356 4448 4679 4450
rect 4356 4392 4618 4448
rect 4674 4392 4679 4448
rect 4356 4390 4679 4392
rect 4356 4388 4362 4390
rect 4613 4387 4679 4390
rect 7465 4450 7531 4453
rect 8569 4450 8635 4453
rect 9121 4450 9187 4453
rect 7465 4448 9187 4450
rect 7465 4392 7470 4448
rect 7526 4392 8574 4448
rect 8630 4392 9126 4448
rect 9182 4392 9187 4448
rect 7465 4390 9187 4392
rect 7465 4387 7531 4390
rect 8569 4387 8635 4390
rect 9121 4387 9187 4390
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 3785 4314 3851 4317
rect 9949 4314 10015 4317
rect 3785 4312 6010 4314
rect 3785 4256 3790 4312
rect 3846 4256 6010 4312
rect 3785 4254 6010 4256
rect 3785 4251 3851 4254
rect 0 4178 800 4208
rect 2497 4178 2563 4181
rect 5717 4180 5783 4181
rect 5717 4178 5764 4180
rect 0 4176 2563 4178
rect 0 4120 2502 4176
rect 2558 4120 2563 4176
rect 0 4118 2563 4120
rect 5672 4176 5764 4178
rect 5672 4120 5722 4176
rect 5672 4118 5764 4120
rect 0 4088 800 4118
rect 2497 4115 2563 4118
rect 5717 4116 5764 4118
rect 5828 4116 5834 4180
rect 5950 4178 6010 4254
rect 6640 4312 10015 4314
rect 6640 4256 9954 4312
rect 10010 4256 10015 4312
rect 6640 4254 10015 4256
rect 6640 4178 6700 4254
rect 9949 4251 10015 4254
rect 11838 4254 16314 4314
rect 5950 4118 6700 4178
rect 9305 4178 9371 4181
rect 9622 4178 9628 4180
rect 9305 4176 9628 4178
rect 9305 4120 9310 4176
rect 9366 4120 9628 4176
rect 9305 4118 9628 4120
rect 5717 4115 5783 4116
rect 9305 4115 9371 4118
rect 9622 4116 9628 4118
rect 9692 4178 9698 4180
rect 11838 4178 11898 4254
rect 14774 4178 14780 4180
rect 9692 4118 11898 4178
rect 12390 4118 14780 4178
rect 9692 4116 9698 4118
rect 5574 3980 5580 4044
rect 5644 4042 5650 4044
rect 6085 4042 6151 4045
rect 5644 4040 6151 4042
rect 5644 3984 6090 4040
rect 6146 3984 6151 4040
rect 5644 3982 6151 3984
rect 5644 3980 5650 3982
rect 6085 3979 6151 3982
rect 7465 4042 7531 4045
rect 7598 4042 7604 4044
rect 7465 4040 7604 4042
rect 7465 3984 7470 4040
rect 7526 3984 7604 4040
rect 7465 3982 7604 3984
rect 7465 3979 7531 3982
rect 7598 3980 7604 3982
rect 7668 3980 7674 4044
rect 10358 4042 10364 4044
rect 7790 3982 10364 4042
rect 4613 3906 4679 3909
rect 4889 3906 4955 3909
rect 7790 3906 7850 3982
rect 10358 3980 10364 3982
rect 10428 3980 10434 4044
rect 11053 4042 11119 4045
rect 12390 4042 12450 4118
rect 14774 4116 14780 4118
rect 14844 4116 14850 4180
rect 16254 4178 16314 4254
rect 20621 4178 20687 4181
rect 16254 4176 20687 4178
rect 16254 4120 20626 4176
rect 20682 4120 20687 4176
rect 16254 4118 20687 4120
rect 20854 4178 20914 4526
rect 22200 4496 23000 4526
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 22200 4178 23000 4208
rect 20854 4118 23000 4178
rect 20621 4115 20687 4118
rect 22200 4088 23000 4118
rect 11053 4040 12450 4042
rect 11053 3984 11058 4040
rect 11114 3984 12450 4040
rect 11053 3982 12450 3984
rect 14273 4042 14339 4045
rect 14406 4042 14412 4044
rect 14273 4040 14412 4042
rect 14273 3984 14278 4040
rect 14334 3984 14412 4040
rect 14273 3982 14412 3984
rect 11053 3979 11119 3982
rect 14273 3979 14339 3982
rect 14406 3980 14412 3982
rect 14476 3980 14482 4044
rect 15142 3980 15148 4044
rect 15212 4042 15218 4044
rect 15929 4042 15995 4045
rect 20437 4044 20503 4045
rect 20437 4042 20484 4044
rect 15212 4040 15995 4042
rect 15212 3984 15934 4040
rect 15990 3984 15995 4040
rect 15212 3982 15995 3984
rect 20392 4040 20484 4042
rect 20392 3984 20442 4040
rect 20392 3982 20484 3984
rect 15212 3980 15218 3982
rect 15929 3979 15995 3982
rect 20437 3980 20484 3982
rect 20548 3980 20554 4044
rect 20437 3979 20503 3980
rect 4613 3904 7850 3906
rect 4613 3848 4618 3904
rect 4674 3848 4894 3904
rect 4950 3848 7850 3904
rect 4613 3846 7850 3848
rect 4613 3843 4679 3846
rect 4889 3843 4955 3846
rect 3545 3840 3861 3841
rect 0 3770 800 3800
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 2773 3770 2839 3773
rect 0 3768 2839 3770
rect 0 3712 2778 3768
rect 2834 3712 2839 3768
rect 0 3710 2839 3712
rect 0 3680 800 3710
rect 2773 3707 2839 3710
rect 19609 3770 19675 3773
rect 22200 3770 23000 3800
rect 19609 3768 23000 3770
rect 19609 3712 19614 3768
rect 19670 3712 23000 3768
rect 19609 3710 23000 3712
rect 19609 3707 19675 3710
rect 22200 3680 23000 3710
rect 1577 3634 1643 3637
rect 4613 3634 4679 3637
rect 1577 3632 4679 3634
rect 1577 3576 1582 3632
rect 1638 3576 4618 3632
rect 4674 3576 4679 3632
rect 1577 3574 4679 3576
rect 1577 3571 1643 3574
rect 4613 3571 4679 3574
rect 5993 3634 6059 3637
rect 6453 3634 6519 3637
rect 9806 3634 9812 3636
rect 5993 3632 9812 3634
rect 5993 3576 5998 3632
rect 6054 3576 6458 3632
rect 6514 3576 9812 3632
rect 5993 3574 9812 3576
rect 5993 3571 6059 3574
rect 6453 3571 6519 3574
rect 9806 3572 9812 3574
rect 9876 3572 9882 3636
rect 12525 3634 12591 3637
rect 16982 3634 16988 3636
rect 12525 3632 16988 3634
rect 12525 3576 12530 3632
rect 12586 3576 16988 3632
rect 12525 3574 16988 3576
rect 12525 3571 12591 3574
rect 16982 3572 16988 3574
rect 17052 3634 17058 3636
rect 19006 3634 19012 3636
rect 17052 3574 19012 3634
rect 17052 3572 17058 3574
rect 19006 3572 19012 3574
rect 19076 3634 19082 3636
rect 19241 3634 19307 3637
rect 19076 3632 19307 3634
rect 19076 3576 19246 3632
rect 19302 3576 19307 3632
rect 19076 3574 19307 3576
rect 19076 3572 19082 3574
rect 19241 3571 19307 3574
rect 4153 3498 4219 3501
rect 14825 3498 14891 3501
rect 4153 3496 14891 3498
rect 4153 3440 4158 3496
rect 4214 3440 14830 3496
rect 14886 3440 14891 3496
rect 4153 3438 14891 3440
rect 4153 3435 4219 3438
rect 14825 3435 14891 3438
rect 18045 3498 18111 3501
rect 18045 3496 22202 3498
rect 18045 3440 18050 3496
rect 18106 3440 22202 3496
rect 18045 3438 22202 3440
rect 18045 3435 18111 3438
rect 22142 3392 22202 3438
rect 0 3362 800 3392
rect 3969 3362 4035 3365
rect 0 3360 4035 3362
rect 0 3304 3974 3360
rect 4030 3304 4035 3360
rect 0 3302 4035 3304
rect 0 3272 800 3302
rect 3969 3299 4035 3302
rect 8201 3362 8267 3365
rect 11094 3362 11100 3364
rect 8201 3360 11100 3362
rect 8201 3304 8206 3360
rect 8262 3304 11100 3360
rect 8201 3302 11100 3304
rect 8201 3299 8267 3302
rect 11094 3300 11100 3302
rect 11164 3300 11170 3364
rect 22142 3302 23000 3392
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 22200 3272 23000 3302
rect 21738 3231 22054 3232
rect 6085 3090 6151 3093
rect 8477 3090 8543 3093
rect 9990 3090 9996 3092
rect 6085 3088 9996 3090
rect 6085 3032 6090 3088
rect 6146 3032 8482 3088
rect 8538 3032 9996 3088
rect 6085 3030 9996 3032
rect 6085 3027 6151 3030
rect 8477 3027 8543 3030
rect 9990 3028 9996 3030
rect 10060 3028 10066 3092
rect 10317 3090 10383 3093
rect 15929 3090 15995 3093
rect 17861 3090 17927 3093
rect 19149 3090 19215 3093
rect 19977 3092 20043 3093
rect 10317 3088 15995 3090
rect 10317 3032 10322 3088
rect 10378 3032 15934 3088
rect 15990 3032 15995 3088
rect 10317 3030 15995 3032
rect 10317 3027 10383 3030
rect 15929 3027 15995 3030
rect 16070 3088 19215 3090
rect 16070 3032 17866 3088
rect 17922 3032 19154 3088
rect 19210 3032 19215 3088
rect 16070 3030 19215 3032
rect 0 2954 800 2984
rect 2405 2954 2471 2957
rect 0 2952 2471 2954
rect 0 2896 2410 2952
rect 2466 2896 2471 2952
rect 0 2894 2471 2896
rect 0 2864 800 2894
rect 2405 2891 2471 2894
rect 4981 2954 5047 2957
rect 9029 2954 9095 2957
rect 4981 2952 9095 2954
rect 4981 2896 4986 2952
rect 5042 2896 9034 2952
rect 9090 2896 9095 2952
rect 4981 2894 9095 2896
rect 4981 2891 5047 2894
rect 9029 2891 9095 2894
rect 11973 2954 12039 2957
rect 14549 2954 14615 2957
rect 16070 2954 16130 3030
rect 17861 3027 17927 3030
rect 19149 3027 19215 3030
rect 19926 3028 19932 3092
rect 19996 3090 20043 3092
rect 19996 3088 20088 3090
rect 20038 3032 20088 3088
rect 19996 3030 20088 3032
rect 19996 3028 20043 3030
rect 19977 3027 20043 3028
rect 16297 2956 16363 2957
rect 11973 2952 16130 2954
rect 11973 2896 11978 2952
rect 12034 2896 14554 2952
rect 14610 2896 16130 2952
rect 11973 2894 16130 2896
rect 11973 2891 12039 2894
rect 14549 2891 14615 2894
rect 16246 2892 16252 2956
rect 16316 2954 16363 2956
rect 18597 2954 18663 2957
rect 22200 2954 23000 2984
rect 16316 2952 16408 2954
rect 16358 2896 16408 2952
rect 16316 2894 16408 2896
rect 18597 2952 23000 2954
rect 18597 2896 18602 2952
rect 18658 2896 23000 2952
rect 18597 2894 23000 2896
rect 16316 2892 16363 2894
rect 16297 2891 16363 2892
rect 18597 2891 18663 2894
rect 22200 2864 23000 2894
rect 8569 2820 8635 2821
rect 8518 2756 8524 2820
rect 8588 2818 8635 2820
rect 8588 2816 8680 2818
rect 8630 2760 8680 2816
rect 8588 2758 8680 2760
rect 8588 2756 8635 2758
rect 8569 2755 8635 2756
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 7649 2682 7715 2685
rect 7782 2682 7788 2684
rect 7649 2680 7788 2682
rect 7649 2624 7654 2680
rect 7710 2624 7788 2680
rect 7649 2622 7788 2624
rect 7649 2619 7715 2622
rect 7782 2620 7788 2622
rect 7852 2620 7858 2684
rect 9254 2620 9260 2684
rect 9324 2682 9330 2684
rect 10593 2682 10659 2685
rect 9324 2680 10659 2682
rect 9324 2624 10598 2680
rect 10654 2624 10659 2680
rect 9324 2622 10659 2624
rect 9324 2620 9330 2622
rect 10593 2619 10659 2622
rect 12249 2682 12315 2685
rect 13486 2682 13492 2684
rect 12249 2680 13492 2682
rect 12249 2624 12254 2680
rect 12310 2624 13492 2680
rect 12249 2622 13492 2624
rect 12249 2619 12315 2622
rect 13486 2620 13492 2622
rect 13556 2620 13562 2684
rect 0 2546 800 2576
rect 3969 2546 4035 2549
rect 0 2544 4035 2546
rect 0 2488 3974 2544
rect 4030 2488 4035 2544
rect 0 2486 4035 2488
rect 0 2456 800 2486
rect 3969 2483 4035 2486
rect 6361 2546 6427 2549
rect 8845 2546 8911 2549
rect 9438 2546 9444 2548
rect 6361 2544 9444 2546
rect 6361 2488 6366 2544
rect 6422 2488 8850 2544
rect 8906 2488 9444 2544
rect 6361 2486 9444 2488
rect 6361 2483 6427 2486
rect 8845 2483 8911 2486
rect 9438 2484 9444 2486
rect 9508 2484 9514 2548
rect 19241 2546 19307 2549
rect 22200 2546 23000 2576
rect 19241 2544 23000 2546
rect 19241 2488 19246 2544
rect 19302 2488 23000 2544
rect 19241 2486 23000 2488
rect 19241 2483 19307 2486
rect 22200 2456 23000 2486
rect 2221 2410 2287 2413
rect 13302 2410 13308 2412
rect 2221 2408 13308 2410
rect 2221 2352 2226 2408
rect 2282 2352 13308 2408
rect 2221 2350 13308 2352
rect 2221 2347 2287 2350
rect 13302 2348 13308 2350
rect 13372 2348 13378 2412
rect 6144 2208 6460 2209
rect 0 2138 800 2168
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 3969 2138 4035 2141
rect 22200 2138 23000 2168
rect 0 2136 4035 2138
rect 0 2080 3974 2136
rect 4030 2080 4035 2136
rect 0 2078 4035 2080
rect 0 2048 800 2078
rect 3969 2075 4035 2078
rect 22142 2048 23000 2138
rect 4429 2002 4495 2005
rect 14590 2002 14596 2004
rect 4429 2000 14596 2002
rect 4429 1944 4434 2000
rect 4490 1944 14596 2000
rect 4429 1942 14596 1944
rect 4429 1939 4495 1942
rect 14590 1940 14596 1942
rect 14660 1940 14666 2004
rect 17493 2002 17559 2005
rect 22142 2002 22202 2048
rect 17493 2000 22202 2002
rect 17493 1944 17498 2000
rect 17554 1944 22202 2000
rect 17493 1942 22202 1944
rect 17493 1939 17559 1942
rect 0 1730 800 1760
rect 2865 1730 2931 1733
rect 0 1728 2931 1730
rect 0 1672 2870 1728
rect 2926 1672 2931 1728
rect 0 1670 2931 1672
rect 0 1640 800 1670
rect 2865 1667 2931 1670
rect 18965 1730 19031 1733
rect 22200 1730 23000 1760
rect 18965 1728 23000 1730
rect 18965 1672 18970 1728
rect 19026 1672 23000 1728
rect 18965 1670 23000 1672
rect 18965 1667 19031 1670
rect 22200 1640 23000 1670
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 16252 19756 16316 19820
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3924 19348 3988 19412
rect 15148 19348 15212 19412
rect 16988 19408 17052 19412
rect 16988 19352 17002 19408
rect 17002 19352 17052 19408
rect 16988 19348 17052 19352
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 5580 18260 5644 18324
rect 8340 18260 8404 18324
rect 8156 17988 8220 18052
rect 12204 17988 12268 18052
rect 13492 17988 13556 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 10732 17852 10796 17916
rect 8156 17444 8220 17508
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 2636 16960 2700 16964
rect 2636 16904 2686 16960
rect 2686 16904 2700 16960
rect 2636 16900 2700 16904
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 5764 16628 5828 16692
rect 7972 16688 8036 16692
rect 7972 16632 7986 16688
rect 7986 16632 8036 16688
rect 7972 16628 8036 16632
rect 9996 16688 10060 16692
rect 9996 16632 10010 16688
rect 10010 16632 10060 16688
rect 9996 16628 10060 16632
rect 10364 16688 10428 16692
rect 10364 16632 10378 16688
rect 10378 16632 10428 16688
rect 10364 16628 10428 16632
rect 13124 16688 13188 16692
rect 13124 16632 13138 16688
rect 13138 16632 13188 16688
rect 13124 16628 13188 16632
rect 14412 16628 14476 16692
rect 17724 16688 17788 16692
rect 17724 16632 17774 16688
rect 17774 16632 17788 16688
rect 17724 16628 17788 16632
rect 20484 16628 20548 16692
rect 8524 16356 8588 16420
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 5396 16084 5460 16148
rect 6868 15948 6932 16012
rect 7236 15812 7300 15876
rect 14780 15812 14844 15876
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 7788 15540 7852 15604
rect 11100 15540 11164 15604
rect 14596 15540 14660 15604
rect 4108 15268 4172 15332
rect 4476 15268 4540 15332
rect 9444 15328 9508 15332
rect 9444 15272 9458 15328
rect 9458 15272 9508 15328
rect 9444 15268 9508 15272
rect 13308 15328 13372 15332
rect 13308 15272 13358 15328
rect 13358 15272 13372 15328
rect 13308 15268 13372 15272
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 8156 15056 8220 15060
rect 8156 15000 8206 15056
rect 8206 15000 8220 15056
rect 8156 14996 8220 15000
rect 14780 14860 14844 14924
rect 12388 14724 12452 14788
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 10180 14452 10244 14516
rect 19012 14452 19076 14516
rect 19932 14180 19996 14244
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 11836 13908 11900 13972
rect 7420 13772 7484 13836
rect 7604 13832 7668 13836
rect 7604 13776 7618 13832
rect 7618 13776 7668 13832
rect 7604 13772 7668 13776
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 7052 13500 7116 13564
rect 2820 13364 2884 13428
rect 6868 13364 6932 13428
rect 3372 13228 3436 13292
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 4476 13016 4540 13020
rect 4476 12960 4526 13016
rect 4526 12960 4540 13016
rect 4476 12956 4540 12960
rect 16252 12820 16316 12884
rect 3004 12608 3068 12612
rect 3004 12552 3054 12608
rect 3054 12552 3068 12608
rect 3004 12548 3068 12552
rect 6684 12608 6748 12612
rect 6684 12552 6698 12608
rect 6698 12552 6748 12608
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 6684 12548 6748 12552
rect 10732 12548 10796 12612
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 12020 12472 12084 12476
rect 12020 12416 12034 12472
rect 12034 12416 12084 12472
rect 12020 12412 12084 12416
rect 7972 12276 8036 12340
rect 12020 12276 12084 12340
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 4108 11596 4172 11660
rect 5212 11596 5276 11660
rect 5948 11460 6012 11524
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 4476 11188 4540 11252
rect 18092 11188 18156 11252
rect 6684 11052 6748 11116
rect 9628 11052 9692 11116
rect 12020 11112 12084 11116
rect 12020 11056 12034 11112
rect 12034 11056 12084 11112
rect 12020 11052 12084 11056
rect 16252 11052 16316 11116
rect 7052 10976 7116 10980
rect 7052 10920 7102 10976
rect 7102 10920 7116 10976
rect 7052 10916 7116 10920
rect 10732 10976 10796 10980
rect 10732 10920 10782 10976
rect 10782 10920 10796 10976
rect 10732 10916 10796 10920
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 3924 10508 3988 10572
rect 7236 10508 7300 10572
rect 12388 10372 12452 10436
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 5396 10296 5460 10300
rect 5396 10240 5446 10296
rect 5446 10240 5460 10296
rect 5396 10236 5460 10240
rect 7420 10296 7484 10300
rect 7420 10240 7470 10296
rect 7470 10240 7484 10296
rect 7420 10236 7484 10240
rect 2084 9964 2148 10028
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 5948 9148 6012 9212
rect 11836 8876 11900 8940
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 4292 8468 4356 8532
rect 5396 8332 5460 8396
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 13124 8060 13188 8124
rect 12204 7924 12268 7988
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 8340 7516 8404 7580
rect 3372 7440 3436 7444
rect 3372 7384 3386 7440
rect 3386 7384 3436 7440
rect 3372 7380 3436 7384
rect 9260 7168 9324 7172
rect 9260 7112 9310 7168
rect 9310 7112 9324 7168
rect 9260 7108 9324 7112
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 2636 6700 2700 6764
rect 15148 6700 15212 6764
rect 16988 6700 17052 6764
rect 19012 6700 19076 6764
rect 16988 6624 17052 6628
rect 16988 6568 17002 6624
rect 17002 6568 17052 6624
rect 16988 6564 17052 6568
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 6868 6428 6932 6492
rect 2084 6292 2148 6356
rect 2820 6156 2884 6220
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 4476 5884 4540 5948
rect 18828 5884 18892 5948
rect 3004 5612 3068 5676
rect 6684 5672 6748 5676
rect 6684 5616 6734 5672
rect 6734 5616 6748 5672
rect 6684 5612 6748 5616
rect 19012 5476 19076 5540
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 17724 5340 17788 5404
rect 18092 5400 18156 5404
rect 18092 5344 18142 5400
rect 18142 5344 18156 5400
rect 18092 5340 18156 5344
rect 10180 5204 10244 5268
rect 5396 5068 5460 5132
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 9812 4796 9876 4860
rect 12020 4796 12084 4860
rect 4292 4388 4356 4452
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 5764 4176 5828 4180
rect 5764 4120 5778 4176
rect 5778 4120 5828 4176
rect 5764 4116 5828 4120
rect 9628 4116 9692 4180
rect 5580 3980 5644 4044
rect 7604 3980 7668 4044
rect 10364 3980 10428 4044
rect 14780 4116 14844 4180
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 14412 3980 14476 4044
rect 15148 3980 15212 4044
rect 20484 4040 20548 4044
rect 20484 3984 20498 4040
rect 20498 3984 20548 4040
rect 20484 3980 20548 3984
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 9812 3572 9876 3636
rect 16988 3572 17052 3636
rect 19012 3572 19076 3636
rect 11100 3300 11164 3364
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 9996 3028 10060 3092
rect 19932 3088 19996 3092
rect 19932 3032 19982 3088
rect 19982 3032 19996 3088
rect 19932 3028 19996 3032
rect 16252 2952 16316 2956
rect 16252 2896 16302 2952
rect 16302 2896 16316 2952
rect 16252 2892 16316 2896
rect 8524 2816 8588 2820
rect 8524 2760 8574 2816
rect 8574 2760 8588 2816
rect 8524 2756 8588 2760
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 7788 2620 7852 2684
rect 9260 2620 9324 2684
rect 13492 2620 13556 2684
rect 9444 2484 9508 2548
rect 13308 2348 13372 2412
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
rect 14596 1940 14660 2004
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 3923 19412 3989 19413
rect 3923 19348 3924 19412
rect 3988 19348 3989 19412
rect 3923 19347 3989 19348
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 2635 16964 2701 16965
rect 2635 16900 2636 16964
rect 2700 16900 2701 16964
rect 2635 16899 2701 16900
rect 2083 10028 2149 10029
rect 2083 9964 2084 10028
rect 2148 9964 2149 10028
rect 2083 9963 2149 9964
rect 2086 6357 2146 9963
rect 2638 6765 2698 16899
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 2819 13428 2885 13429
rect 2819 13364 2820 13428
rect 2884 13364 2885 13428
rect 2819 13363 2885 13364
rect 2635 6764 2701 6765
rect 2635 6700 2636 6764
rect 2700 6700 2701 6764
rect 2635 6699 2701 6700
rect 2083 6356 2149 6357
rect 2083 6292 2084 6356
rect 2148 6292 2149 6356
rect 2083 6291 2149 6292
rect 2822 6221 2882 13363
rect 3371 13292 3437 13293
rect 3371 13228 3372 13292
rect 3436 13228 3437 13292
rect 3371 13227 3437 13228
rect 3003 12612 3069 12613
rect 3003 12548 3004 12612
rect 3068 12548 3069 12612
rect 3003 12547 3069 12548
rect 2819 6220 2885 6221
rect 2819 6156 2820 6220
rect 2884 6156 2885 6220
rect 2819 6155 2885 6156
rect 3006 5677 3066 12547
rect 3374 7445 3434 13227
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3926 10573 3986 19347
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 5579 18324 5645 18325
rect 5579 18260 5580 18324
rect 5644 18260 5645 18324
rect 5579 18259 5645 18260
rect 5395 16148 5461 16149
rect 5395 16084 5396 16148
rect 5460 16084 5461 16148
rect 5395 16083 5461 16084
rect 4107 15332 4173 15333
rect 4107 15268 4108 15332
rect 4172 15268 4173 15332
rect 4107 15267 4173 15268
rect 4475 15332 4541 15333
rect 4475 15268 4476 15332
rect 4540 15268 4541 15332
rect 4475 15267 4541 15268
rect 4110 11661 4170 15267
rect 4478 13021 4538 15267
rect 4475 13020 4541 13021
rect 4475 12956 4476 13020
rect 4540 12956 4541 13020
rect 4475 12955 4541 12956
rect 4107 11660 4173 11661
rect 4107 11596 4108 11660
rect 4172 11596 4173 11660
rect 4107 11595 4173 11596
rect 5211 11660 5277 11661
rect 5211 11596 5212 11660
rect 5276 11596 5277 11660
rect 5211 11595 5277 11596
rect 4475 11252 4541 11253
rect 4475 11188 4476 11252
rect 4540 11188 4541 11252
rect 4475 11187 4541 11188
rect 3923 10572 3989 10573
rect 3923 10508 3924 10572
rect 3988 10508 3989 10572
rect 3923 10507 3989 10508
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 4291 8532 4357 8533
rect 4291 8468 4292 8532
rect 4356 8468 4357 8532
rect 4291 8467 4357 8468
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3371 7444 3437 7445
rect 3371 7380 3372 7444
rect 3436 7380 3437 7444
rect 3371 7379 3437 7380
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3003 5676 3069 5677
rect 3003 5612 3004 5676
rect 3068 5612 3069 5676
rect 3003 5611 3069 5612
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 4294 4453 4354 8467
rect 4478 5949 4538 11187
rect 5214 9890 5274 11595
rect 5398 10301 5458 16083
rect 5395 10300 5461 10301
rect 5395 10236 5396 10300
rect 5460 10236 5461 10300
rect 5395 10235 5461 10236
rect 5214 9830 5458 9890
rect 5398 8397 5458 9830
rect 5395 8396 5461 8397
rect 5395 8332 5396 8396
rect 5460 8332 5461 8396
rect 5395 8331 5461 8332
rect 4475 5948 4541 5949
rect 4475 5884 4476 5948
rect 4540 5884 4541 5948
rect 4475 5883 4541 5884
rect 5398 5133 5458 8331
rect 5395 5132 5461 5133
rect 5395 5068 5396 5132
rect 5460 5068 5461 5132
rect 5395 5067 5461 5068
rect 4291 4452 4357 4453
rect 4291 4388 4292 4452
rect 4356 4388 4357 4452
rect 4291 4387 4357 4388
rect 5582 4045 5642 18259
rect 6142 17440 6462 18464
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8339 18324 8405 18325
rect 8339 18260 8340 18324
rect 8404 18260 8405 18324
rect 8339 18259 8405 18260
rect 8155 18052 8221 18053
rect 8155 17988 8156 18052
rect 8220 17988 8221 18052
rect 8155 17987 8221 17988
rect 8158 17509 8218 17987
rect 8155 17508 8221 17509
rect 8155 17444 8156 17508
rect 8220 17444 8221 17508
rect 8155 17443 8221 17444
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 5763 16692 5829 16693
rect 5763 16628 5764 16692
rect 5828 16628 5829 16692
rect 5763 16627 5829 16628
rect 5766 4181 5826 16627
rect 6142 16352 6462 17376
rect 7971 16692 8037 16693
rect 7971 16628 7972 16692
rect 8036 16628 8037 16692
rect 7971 16627 8037 16628
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6867 16012 6933 16013
rect 6867 15948 6868 16012
rect 6932 15948 6933 16012
rect 6867 15947 6933 15948
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6870 13429 6930 15947
rect 7235 15876 7301 15877
rect 7235 15812 7236 15876
rect 7300 15812 7301 15876
rect 7235 15811 7301 15812
rect 7051 13564 7117 13565
rect 7051 13500 7052 13564
rect 7116 13500 7117 13564
rect 7051 13499 7117 13500
rect 6867 13428 6933 13429
rect 6867 13364 6868 13428
rect 6932 13364 6933 13428
rect 6867 13363 6933 13364
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6683 12612 6749 12613
rect 6683 12548 6684 12612
rect 6748 12548 6749 12612
rect 6683 12547 6749 12548
rect 6686 12450 6746 12547
rect 6686 12390 6930 12450
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 5947 11524 6013 11525
rect 5947 11460 5948 11524
rect 6012 11460 6013 11524
rect 5947 11459 6013 11460
rect 5950 9213 6010 11459
rect 6142 10912 6462 11936
rect 6683 11116 6749 11117
rect 6683 11052 6684 11116
rect 6748 11052 6749 11116
rect 6683 11051 6749 11052
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 5947 9212 6013 9213
rect 5947 9148 5948 9212
rect 6012 9148 6013 9212
rect 5947 9147 6013 9148
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6686 5677 6746 11051
rect 6870 6493 6930 12390
rect 7054 10981 7114 13499
rect 7051 10980 7117 10981
rect 7051 10916 7052 10980
rect 7116 10916 7117 10980
rect 7051 10915 7117 10916
rect 7238 10573 7298 15811
rect 7787 15604 7853 15605
rect 7787 15540 7788 15604
rect 7852 15540 7853 15604
rect 7787 15539 7853 15540
rect 7419 13836 7485 13837
rect 7419 13772 7420 13836
rect 7484 13772 7485 13836
rect 7419 13771 7485 13772
rect 7603 13836 7669 13837
rect 7603 13772 7604 13836
rect 7668 13772 7669 13836
rect 7603 13771 7669 13772
rect 7235 10572 7301 10573
rect 7235 10508 7236 10572
rect 7300 10508 7301 10572
rect 7235 10507 7301 10508
rect 7422 10301 7482 13771
rect 7419 10300 7485 10301
rect 7419 10236 7420 10300
rect 7484 10236 7485 10300
rect 7419 10235 7485 10236
rect 6867 6492 6933 6493
rect 6867 6428 6868 6492
rect 6932 6428 6933 6492
rect 6867 6427 6933 6428
rect 6683 5676 6749 5677
rect 6683 5612 6684 5676
rect 6748 5612 6749 5676
rect 6683 5611 6749 5612
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 5763 4180 5829 4181
rect 5763 4116 5764 4180
rect 5828 4116 5829 4180
rect 5763 4115 5829 4116
rect 5579 4044 5645 4045
rect 5579 3980 5580 4044
rect 5644 3980 5645 4044
rect 5579 3979 5645 3980
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 3296 6462 4320
rect 7606 4045 7666 13771
rect 7603 4044 7669 4045
rect 7603 3980 7604 4044
rect 7668 3980 7669 4044
rect 7603 3979 7669 3980
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 7790 2685 7850 15539
rect 7974 12341 8034 16627
rect 8158 15061 8218 17443
rect 8155 15060 8221 15061
rect 8155 14996 8156 15060
rect 8220 14996 8221 15060
rect 8155 14995 8221 14996
rect 7971 12340 8037 12341
rect 7971 12276 7972 12340
rect 8036 12276 8037 12340
rect 7971 12275 8037 12276
rect 8342 7581 8402 18259
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 10731 17916 10797 17917
rect 10731 17852 10732 17916
rect 10796 17852 10797 17916
rect 10731 17851 10797 17852
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8523 16420 8589 16421
rect 8523 16356 8524 16420
rect 8588 16356 8589 16420
rect 8523 16355 8589 16356
rect 8339 7580 8405 7581
rect 8339 7516 8340 7580
rect 8404 7516 8405 7580
rect 8339 7515 8405 7516
rect 8526 2821 8586 16355
rect 8741 15808 9061 16832
rect 9995 16692 10061 16693
rect 9995 16628 9996 16692
rect 10060 16628 10061 16692
rect 9995 16627 10061 16628
rect 10363 16692 10429 16693
rect 10363 16628 10364 16692
rect 10428 16628 10429 16692
rect 10363 16627 10429 16628
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 9443 15332 9509 15333
rect 9443 15268 9444 15332
rect 9508 15268 9509 15332
rect 9443 15267 9509 15268
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 9259 7172 9325 7173
rect 9259 7108 9260 7172
rect 9324 7108 9325 7172
rect 9259 7107 9325 7108
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8523 2820 8589 2821
rect 8523 2756 8524 2820
rect 8588 2756 8589 2820
rect 8523 2755 8589 2756
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 7787 2684 7853 2685
rect 7787 2620 7788 2684
rect 7852 2620 7853 2684
rect 7787 2619 7853 2620
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 2128 9061 2688
rect 9262 2685 9322 7107
rect 9259 2684 9325 2685
rect 9259 2620 9260 2684
rect 9324 2620 9325 2684
rect 9259 2619 9325 2620
rect 9446 2549 9506 15267
rect 9627 11116 9693 11117
rect 9627 11052 9628 11116
rect 9692 11052 9693 11116
rect 9627 11051 9693 11052
rect 9630 4181 9690 11051
rect 9811 4860 9877 4861
rect 9811 4796 9812 4860
rect 9876 4796 9877 4860
rect 9811 4795 9877 4796
rect 9627 4180 9693 4181
rect 9627 4116 9628 4180
rect 9692 4116 9693 4180
rect 9627 4115 9693 4116
rect 9814 3637 9874 4795
rect 9811 3636 9877 3637
rect 9811 3572 9812 3636
rect 9876 3572 9877 3636
rect 9811 3571 9877 3572
rect 9998 3093 10058 16627
rect 10179 14516 10245 14517
rect 10179 14452 10180 14516
rect 10244 14452 10245 14516
rect 10179 14451 10245 14452
rect 10182 5269 10242 14451
rect 10179 5268 10245 5269
rect 10179 5204 10180 5268
rect 10244 5204 10245 5268
rect 10179 5203 10245 5204
rect 10366 4045 10426 16627
rect 10734 12613 10794 17851
rect 11340 17440 11660 18464
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16251 19820 16317 19821
rect 16251 19756 16252 19820
rect 16316 19756 16317 19820
rect 16251 19755 16317 19756
rect 15147 19412 15213 19413
rect 15147 19348 15148 19412
rect 15212 19348 15213 19412
rect 15147 19347 15213 19348
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 12203 18052 12269 18053
rect 12203 17988 12204 18052
rect 12268 17988 12269 18052
rect 12203 17987 12269 17988
rect 13491 18052 13557 18053
rect 13491 17988 13492 18052
rect 13556 17988 13557 18052
rect 13491 17987 13557 17988
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11099 15604 11165 15605
rect 11099 15540 11100 15604
rect 11164 15540 11165 15604
rect 11099 15539 11165 15540
rect 10731 12612 10797 12613
rect 10731 12548 10732 12612
rect 10796 12548 10797 12612
rect 10731 12547 10797 12548
rect 10734 10981 10794 12547
rect 10731 10980 10797 10981
rect 10731 10916 10732 10980
rect 10796 10916 10797 10980
rect 10731 10915 10797 10916
rect 10363 4044 10429 4045
rect 10363 3980 10364 4044
rect 10428 3980 10429 4044
rect 10363 3979 10429 3980
rect 11102 3365 11162 15539
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11835 13972 11901 13973
rect 11835 13908 11836 13972
rect 11900 13908 11901 13972
rect 11835 13907 11901 13908
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11838 8941 11898 13907
rect 12019 12476 12085 12477
rect 12019 12412 12020 12476
rect 12084 12412 12085 12476
rect 12019 12411 12085 12412
rect 12022 12341 12082 12411
rect 12019 12340 12085 12341
rect 12019 12276 12020 12340
rect 12084 12276 12085 12340
rect 12019 12275 12085 12276
rect 12019 11116 12085 11117
rect 12019 11052 12020 11116
rect 12084 11052 12085 11116
rect 12019 11051 12085 11052
rect 11835 8940 11901 8941
rect 11835 8876 11836 8940
rect 11900 8876 11901 8940
rect 11835 8875 11901 8876
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 12022 4861 12082 11051
rect 12206 7989 12266 17987
rect 13123 16692 13189 16693
rect 13123 16628 13124 16692
rect 13188 16628 13189 16692
rect 13123 16627 13189 16628
rect 12387 14788 12453 14789
rect 12387 14724 12388 14788
rect 12452 14724 12453 14788
rect 12387 14723 12453 14724
rect 12390 10437 12450 14723
rect 12387 10436 12453 10437
rect 12387 10372 12388 10436
rect 12452 10372 12453 10436
rect 12387 10371 12453 10372
rect 13126 8125 13186 16627
rect 13307 15332 13373 15333
rect 13307 15268 13308 15332
rect 13372 15268 13373 15332
rect 13307 15267 13373 15268
rect 13123 8124 13189 8125
rect 13123 8060 13124 8124
rect 13188 8060 13189 8124
rect 13123 8059 13189 8060
rect 12203 7988 12269 7989
rect 12203 7924 12204 7988
rect 12268 7924 12269 7988
rect 12203 7923 12269 7924
rect 12019 4860 12085 4861
rect 12019 4796 12020 4860
rect 12084 4796 12085 4860
rect 12019 4795 12085 4796
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11099 3364 11165 3365
rect 11099 3300 11100 3364
rect 11164 3300 11165 3364
rect 11099 3299 11165 3300
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 9995 3092 10061 3093
rect 9995 3028 9996 3092
rect 10060 3028 10061 3092
rect 9995 3027 10061 3028
rect 9443 2548 9509 2549
rect 9443 2484 9444 2548
rect 9508 2484 9509 2548
rect 9443 2483 9509 2484
rect 11340 2208 11660 3232
rect 13310 2413 13370 15267
rect 13494 2685 13554 17987
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 14411 16692 14477 16693
rect 14411 16628 14412 16692
rect 14476 16628 14477 16692
rect 14411 16627 14477 16628
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 14414 4045 14474 16627
rect 14779 15876 14845 15877
rect 14779 15812 14780 15876
rect 14844 15812 14845 15876
rect 14779 15811 14845 15812
rect 14595 15604 14661 15605
rect 14595 15540 14596 15604
rect 14660 15540 14661 15604
rect 14595 15539 14661 15540
rect 14411 4044 14477 4045
rect 14411 3980 14412 4044
rect 14476 3980 14477 4044
rect 14411 3979 14477 3980
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13491 2684 13557 2685
rect 13491 2620 13492 2684
rect 13556 2620 13557 2684
rect 13491 2619 13557 2620
rect 13307 2412 13373 2413
rect 13307 2348 13308 2412
rect 13372 2348 13373 2412
rect 13307 2347 13373 2348
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 2128 14259 2688
rect 14598 2005 14658 15539
rect 14782 14925 14842 15811
rect 14779 14924 14845 14925
rect 14779 14860 14780 14924
rect 14844 14860 14845 14924
rect 14779 14859 14845 14860
rect 14782 4181 14842 14859
rect 15150 6765 15210 19347
rect 16254 12885 16314 19755
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 16987 19412 17053 19413
rect 16987 19348 16988 19412
rect 17052 19348 17053 19412
rect 16987 19347 17053 19348
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16251 12884 16317 12885
rect 16251 12820 16252 12884
rect 16316 12820 16317 12884
rect 16251 12819 16317 12820
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16251 11116 16317 11117
rect 16251 11052 16252 11116
rect 16316 11052 16317 11116
rect 16251 11051 16317 11052
rect 15147 6764 15213 6765
rect 15147 6700 15148 6764
rect 15212 6700 15213 6764
rect 15147 6699 15213 6700
rect 14779 4180 14845 4181
rect 14779 4116 14780 4180
rect 14844 4116 14845 4180
rect 14779 4115 14845 4116
rect 15150 4045 15210 6699
rect 15147 4044 15213 4045
rect 15147 3980 15148 4044
rect 15212 3980 15213 4044
rect 15147 3979 15213 3980
rect 16254 2957 16314 11051
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16990 6765 17050 19347
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 17723 16692 17789 16693
rect 17723 16628 17724 16692
rect 17788 16628 17789 16692
rect 17723 16627 17789 16628
rect 16987 6764 17053 6765
rect 16987 6700 16988 6764
rect 17052 6700 17053 6764
rect 16987 6699 17053 6700
rect 16987 6628 17053 6629
rect 16987 6564 16988 6628
rect 17052 6564 17053 6628
rect 16987 6563 17053 6564
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16990 3637 17050 6563
rect 17726 5405 17786 16627
rect 19137 15808 19457 16832
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 20483 16692 20549 16693
rect 20483 16628 20484 16692
rect 20548 16628 20549 16692
rect 20483 16627 20549 16628
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19011 14516 19077 14517
rect 19011 14452 19012 14516
rect 19076 14452 19077 14516
rect 19011 14451 19077 14452
rect 18091 11252 18157 11253
rect 18091 11188 18092 11252
rect 18156 11188 18157 11252
rect 18091 11187 18157 11188
rect 18094 5405 18154 11187
rect 19014 6765 19074 14451
rect 19137 13632 19457 14656
rect 19931 14244 19997 14245
rect 19931 14180 19932 14244
rect 19996 14180 19997 14244
rect 19931 14179 19997 14180
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19011 6764 19077 6765
rect 19011 6700 19012 6764
rect 19076 6700 19077 6764
rect 19011 6699 19077 6700
rect 19014 6490 19074 6699
rect 18830 6430 19074 6490
rect 18830 5949 18890 6430
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 18827 5948 18893 5949
rect 18827 5884 18828 5948
rect 18892 5884 18893 5948
rect 18827 5883 18893 5884
rect 19011 5540 19077 5541
rect 19011 5476 19012 5540
rect 19076 5476 19077 5540
rect 19011 5475 19077 5476
rect 17723 5404 17789 5405
rect 17723 5340 17724 5404
rect 17788 5340 17789 5404
rect 17723 5339 17789 5340
rect 18091 5404 18157 5405
rect 18091 5340 18092 5404
rect 18156 5340 18157 5404
rect 18091 5339 18157 5340
rect 19014 3637 19074 5475
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 16987 3636 17053 3637
rect 16987 3572 16988 3636
rect 17052 3572 17053 3636
rect 16987 3571 17053 3572
rect 19011 3636 19077 3637
rect 19011 3572 19012 3636
rect 19076 3572 19077 3636
rect 19011 3571 19077 3572
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16251 2956 16317 2957
rect 16251 2892 16252 2956
rect 16316 2892 16317 2956
rect 16251 2891 16317 2892
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 2752 19457 3776
rect 19934 3093 19994 14179
rect 20486 4045 20546 16627
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 20483 4044 20549 4045
rect 20483 3980 20484 4044
rect 20548 3980 20549 4044
rect 20483 3979 20549 3980
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 19931 3092 19997 3093
rect 19931 3028 19932 3092
rect 19996 3028 19997 3092
rect 19931 3027 19997 3028
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
rect 14595 2004 14661 2005
rect 14595 1940 14596 2004
rect 14660 1940 14661 2004
rect 14595 1939 14661 1940
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2944 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1649977179
transform 1 0 5888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1649977179
transform -1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1649977179
transform -1 0 2116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1649977179
transform 1 0 5336 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1649977179
transform -1 0 3864 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1649977179
transform -1 0 5152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1649977179
transform -1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1649977179
transform -1 0 3496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1649977179
transform -1 0 4324 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform -1 0 3956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1649977179
transform 1 0 4508 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1649977179
transform 1 0 18032 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform 1 0 17940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform 1 0 18400 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1649977179
transform 1 0 11960 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1649977179
transform -1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform -1 0 16100 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform 1 0 12328 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform 1 0 15824 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform -1 0 14536 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform -1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 13524 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 10212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 9384 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 5428 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 12420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 6440 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 11868 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 4416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 6624 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 6072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 6532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 5980 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 8096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 3128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 4048 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 9476 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 6440 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 12972 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 8004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 8188 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 8372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 15088 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 12880 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 14628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 14536 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 17020 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 15456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 15640 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 17112 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 11224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 14352 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 12696 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 11592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 9476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 3680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 10580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 9108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 11684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 6808 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 12604 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 12052 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 9016 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 5612 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform 1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 8280 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 8464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 8372 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 12788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 5060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 14076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 12420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1649977179
transform -1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 11776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13156 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10396 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12880 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10580 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10948 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10580 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13340 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17112 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17296 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 14812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1649977179
transform -1 0 18492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18676 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 18492 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13800 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 11500 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1649977179
transform 1 0 17204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 12144 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15272 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14720 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10948 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13432 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 13708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.delay_buf_A
timestamp 1649977179
transform 1 0 11776 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 14444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 18768 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15088 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12052 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 11592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11960 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 19412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15640 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 14444 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20700 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 17020 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14628 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16008 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 17296 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 12604 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 6072 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 12788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10672 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 11868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 12972 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12052 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5888 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 9844 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9108 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6900 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7268 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6532 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9476 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10764 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 8280 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 6808 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8096 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 6624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4416 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9200 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11316 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12696 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12788 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13064 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform -1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 18676 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 15364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 17112 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7360 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6992 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 6624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 5336 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 5520 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 5704 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1649977179
transform -1 0 4784 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1649977179
transform 1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5244 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 3404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_4__A0
timestamp 1649977179
transform -1 0 11684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 5612 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 6716 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1649977179
transform -1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7452 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9200 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 6992 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 7360 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 8648 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 4232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 4600 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7268 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 6072 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 11868 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 4324 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 4048 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8372 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8004 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 8740 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 5888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 5520 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 17572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 14536 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3772 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 4416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 17480 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 17112 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1649977179
transform 1 0 16744 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 14168 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7452 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9844 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1649977179
transform -1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1649977179
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1649977179
transform 1 0 18032 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 18400 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6716 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 7452 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6624 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8004 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 8832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14260 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14536 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 15916 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 14996 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 14076 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 16468 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 11684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 8648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 14536 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 16468 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 18032 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__S
timestamp 1649977179
transform -1 0 12604 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 14628 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 12328 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1649977179
transform -1 0 13248 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1649977179
transform 1 0 12696 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 13984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1649977179
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1649977179
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1649977179
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_122
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_135
timestamp 1649977179
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_179
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1649977179
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_201
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_207
timestamp 1649977179
transform 1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_211
timestamp 1649977179
transform 1 0 20516 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_20
timestamp 1649977179
transform 1 0 2944 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_25
timestamp 1649977179
transform 1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_30
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1649977179
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_47
timestamp 1649977179
transform 1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_60
timestamp 1649977179
transform 1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_65
timestamp 1649977179
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_89
timestamp 1649977179
transform 1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_100
timestamp 1649977179
transform 1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_104
timestamp 1649977179
transform 1 0 10672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_109
timestamp 1649977179
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1649977179
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1649977179
transform 1 0 13984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_146
timestamp 1649977179
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_153
timestamp 1649977179
transform 1 0 15180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1649977179
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_179
timestamp 1649977179
transform 1 0 17572 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_191
timestamp 1649977179
transform 1 0 18676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_202
timestamp 1649977179
transform 1 0 19688 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_216
timestamp 1649977179
transform 1 0 20976 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_38
timestamp 1649977179
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_50
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_54
timestamp 1649977179
transform 1 0 6072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_64
timestamp 1649977179
transform 1 0 6992 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1649977179
transform 1 0 10488 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_120
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_125
timestamp 1649977179
transform 1 0 12604 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_130
timestamp 1649977179
transform 1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1649977179
transform 1 0 14352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_164
timestamp 1649977179
transform 1 0 16192 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_169
timestamp 1649977179
transform 1 0 16652 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_174
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1649977179
transform 1 0 18308 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1649977179
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1649977179
transform 1 0 19596 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_211
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1649977179
transform 1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_24
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_28
timestamp 1649977179
transform 1 0 3680 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_33
timestamp 1649977179
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_49
timestamp 1649977179
transform 1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_67
timestamp 1649977179
transform 1 0 7268 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp 1649977179
transform 1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_77
timestamp 1649977179
transform 1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1649977179
transform 1 0 8648 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_87
timestamp 1649977179
transform 1 0 9108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1649977179
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1649977179
transform 1 0 13156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_154
timestamp 1649977179
transform 1 0 15272 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_159
timestamp 1649977179
transform 1 0 15732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_178
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_185
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_203
timestamp 1649977179
transform 1 0 19780 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1649977179
transform 1 0 20240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1649977179
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_31
timestamp 1649977179
transform 1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_42
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_64
timestamp 1649977179
transform 1 0 6992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_70
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_75
timestamp 1649977179
transform 1 0 8004 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_99
timestamp 1649977179
transform 1 0 10212 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_103
timestamp 1649977179
transform 1 0 10580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_108
timestamp 1649977179
transform 1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_126
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_130
timestamp 1649977179
transform 1 0 13064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_134
timestamp 1649977179
transform 1 0 13432 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_157
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_164
timestamp 1649977179
transform 1 0 16192 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_169
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_175
timestamp 1649977179
transform 1 0 17204 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1649977179
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_199
timestamp 1649977179
transform 1 0 19412 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_205
timestamp 1649977179
transform 1 0 19964 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_217
timestamp 1649977179
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_20
timestamp 1649977179
transform 1 0 2944 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_25
timestamp 1649977179
transform 1 0 3404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_30
timestamp 1649977179
transform 1 0 3864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_35
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_40
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1649977179
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_67
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_78
timestamp 1649977179
transform 1 0 8280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_103
timestamp 1649977179
transform 1 0 10580 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1649977179
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1649977179
transform 1 0 11960 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_136
timestamp 1649977179
transform 1 0 13616 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_140
timestamp 1649977179
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_146
timestamp 1649977179
transform 1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_151
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1649977179
transform 1 0 15456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_180
timestamp 1649977179
transform 1 0 17664 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_185
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_191
timestamp 1649977179
transform 1 0 18676 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_196
timestamp 1649977179
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_214
timestamp 1649977179
transform 1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1649977179
transform 1 0 21436 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1649977179
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_58
timestamp 1649977179
transform 1 0 6440 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_63
timestamp 1649977179
transform 1 0 6900 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_68
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_72
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1649977179
transform 1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_106
timestamp 1649977179
transform 1 0 10856 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1649977179
transform 1 0 12512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_128
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_143
timestamp 1649977179
transform 1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_166
timestamp 1649977179
transform 1 0 16376 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_171
timestamp 1649977179
transform 1 0 16836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1649977179
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_22
timestamp 1649977179
transform 1 0 3128 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_40
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_45
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_49
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_64
timestamp 1649977179
transform 1 0 6992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_78
timestamp 1649977179
transform 1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_82
timestamp 1649977179
transform 1 0 8648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_86
timestamp 1649977179
transform 1 0 9016 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_115
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 1649977179
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_122
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_126
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_145
timestamp 1649977179
transform 1 0 14444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_186
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_192
timestamp 1649977179
transform 1 0 18768 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_198
timestamp 1649977179
transform 1 0 19320 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_209
timestamp 1649977179
transform 1 0 20332 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1649977179
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_38
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_42
timestamp 1649977179
transform 1 0 4968 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_52
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_56
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1649977179
transform 1 0 7176 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_103
timestamp 1649977179
transform 1 0 10580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_124
timestamp 1649977179
transform 1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_132
timestamp 1649977179
transform 1 0 13248 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_152
timestamp 1649977179
transform 1 0 15088 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_156
timestamp 1649977179
transform 1 0 15456 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_169
timestamp 1649977179
transform 1 0 16652 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_174
timestamp 1649977179
transform 1 0 17112 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_185
timestamp 1649977179
transform 1 0 18124 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_213
timestamp 1649977179
transform 1 0 20700 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_14
timestamp 1649977179
transform 1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_20
timestamp 1649977179
transform 1 0 2944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_25
timestamp 1649977179
transform 1 0 3404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_47
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1649977179
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_75
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1649977179
transform 1 0 8372 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1649977179
transform 1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_87
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1649977179
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_115
timestamp 1649977179
transform 1 0 11684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1649977179
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1649977179
transform 1 0 12420 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_133
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_141
timestamp 1649977179
transform 1 0 14076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp 1649977179
transform 1 0 14444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1649977179
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_171
timestamp 1649977179
transform 1 0 16836 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_175
timestamp 1649977179
transform 1 0 17204 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1649977179
transform 1 0 17572 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_190
timestamp 1649977179
transform 1 0 18584 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_210
timestamp 1649977179
transform 1 0 20424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_14
timestamp 1649977179
transform 1 0 2392 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_20
timestamp 1649977179
transform 1 0 2944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1649977179
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1649977179
transform 1 0 4048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 1649977179
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_40
timestamp 1649977179
transform 1 0 4784 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_50
timestamp 1649977179
transform 1 0 5704 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_54
timestamp 1649977179
transform 1 0 6072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_67
timestamp 1649977179
transform 1 0 7268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_78
timestamp 1649977179
transform 1 0 8280 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_87
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_106
timestamp 1649977179
transform 1 0 10856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_110
timestamp 1649977179
transform 1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_114
timestamp 1649977179
transform 1 0 11592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_117
timestamp 1649977179
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_132
timestamp 1649977179
transform 1 0 13248 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1649977179
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_157
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_160
timestamp 1649977179
transform 1 0 15824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_164
timestamp 1649977179
transform 1 0 16192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_168
timestamp 1649977179
transform 1 0 16560 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_187
timestamp 1649977179
transform 1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1649977179
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_214
timestamp 1649977179
transform 1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_13
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_24
timestamp 1649977179
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_29
timestamp 1649977179
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_33
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_38
timestamp 1649977179
transform 1 0 4600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_49
timestamp 1649977179
transform 1 0 5612 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1649977179
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_63
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1649977179
transform 1 0 8280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_88
timestamp 1649977179
transform 1 0 9200 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp 1649977179
transform 1 0 10856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_116
timestamp 1649977179
transform 1 0 11776 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_134
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_138
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_142
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_148
timestamp 1649977179
transform 1 0 14720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_152
timestamp 1649977179
transform 1 0 15088 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_156
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_160
timestamp 1649977179
transform 1 0 15824 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_185
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_189
timestamp 1649977179
transform 1 0 18492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_204
timestamp 1649977179
transform 1 0 19872 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_215
timestamp 1649977179
transform 1 0 20884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_13
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_19
timestamp 1649977179
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1649977179
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_38
timestamp 1649977179
transform 1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1649977179
transform 1 0 5704 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_54
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1649977179
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_62
timestamp 1649977179
transform 1 0 6808 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1649977179
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_76
timestamp 1649977179
transform 1 0 8096 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1649977179
transform 1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_115
timestamp 1649977179
transform 1 0 11684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_158
timestamp 1649977179
transform 1 0 15640 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_162
timestamp 1649977179
transform 1 0 16008 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_179
timestamp 1649977179
transform 1 0 17572 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_185
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1649977179
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_201
timestamp 1649977179
transform 1 0 19596 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_212
timestamp 1649977179
transform 1 0 20608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_216
timestamp 1649977179
transform 1 0 20976 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_5
timestamp 1649977179
transform 1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1649977179
transform 1 0 2576 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_33
timestamp 1649977179
transform 1 0 4140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_38
timestamp 1649977179
transform 1 0 4600 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_49
timestamp 1649977179
transform 1 0 5612 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1649977179
transform 1 0 6808 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1649977179
transform 1 0 8188 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1649977179
transform 1 0 8648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp 1649977179
transform 1 0 9016 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_104
timestamp 1649977179
transform 1 0 10672 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1649977179
transform 1 0 13248 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_136
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1649977179
transform 1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_159
timestamp 1649977179
transform 1 0 15732 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_182
timestamp 1649977179
transform 1 0 17848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_186
timestamp 1649977179
transform 1 0 18216 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_203
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_209
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_21
timestamp 1649977179
transform 1 0 3036 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_31
timestamp 1649977179
transform 1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_42
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_54
timestamp 1649977179
transform 1 0 6072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1649977179
transform 1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_101
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp 1649977179
transform 1 0 10764 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_110
timestamp 1649977179
transform 1 0 11224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_114
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_119
timestamp 1649977179
transform 1 0 12052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_143
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_147
timestamp 1649977179
transform 1 0 14628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1649977179
transform 1 0 14996 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_169
timestamp 1649977179
transform 1 0 16652 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_187
timestamp 1649977179
transform 1 0 18308 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_191
timestamp 1649977179
transform 1 0 18676 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_203
timestamp 1649977179
transform 1 0 19780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 1649977179
transform 1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_29
timestamp 1649977179
transform 1 0 3772 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_33
timestamp 1649977179
transform 1 0 4140 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_43
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_59
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_65
timestamp 1649977179
transform 1 0 7084 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_73
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_84
timestamp 1649977179
transform 1 0 8832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_103
timestamp 1649977179
transform 1 0 10580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1649977179
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_116
timestamp 1649977179
transform 1 0 11776 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_124
timestamp 1649977179
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_128
timestamp 1649977179
transform 1 0 12880 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_147
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_151
timestamp 1649977179
transform 1 0 14996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_155
timestamp 1649977179
transform 1 0 15364 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1649977179
transform 1 0 16008 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1649977179
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_171
timestamp 1649977179
transform 1 0 16836 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1649977179
transform 1 0 17204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_212
timestamp 1649977179
transform 1 0 20608 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_216
timestamp 1649977179
transform 1 0 20976 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_14
timestamp 1649977179
transform 1 0 2392 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp 1649977179
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_33
timestamp 1649977179
transform 1 0 4140 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_46
timestamp 1649977179
transform 1 0 5336 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_58
timestamp 1649977179
transform 1 0 6440 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_63
timestamp 1649977179
transform 1 0 6900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_74
timestamp 1649977179
transform 1 0 7912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_78
timestamp 1649977179
transform 1 0 8280 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_103
timestamp 1649977179
transform 1 0 10580 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_107
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_111
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_131
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_146
timestamp 1649977179
transform 1 0 14536 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_150
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_156
timestamp 1649977179
transform 1 0 15456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_160
timestamp 1649977179
transform 1 0 15824 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_164
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_168
timestamp 1649977179
transform 1 0 16560 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_173
timestamp 1649977179
transform 1 0 17020 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_181
timestamp 1649977179
transform 1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_185
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_214
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_13
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_24
timestamp 1649977179
transform 1 0 3312 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_28
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_38
timestamp 1649977179
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_47
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_59
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_72
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_76
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_80
timestamp 1649977179
transform 1 0 8464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_121
timestamp 1649977179
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_129
timestamp 1649977179
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_148
timestamp 1649977179
transform 1 0 14720 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_185
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_189
timestamp 1649977179
transform 1 0 18492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_197
timestamp 1649977179
transform 1 0 19228 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_208
timestamp 1649977179
transform 1 0 20240 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1649977179
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_13
timestamp 1649977179
transform 1 0 2300 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_38
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_42
timestamp 1649977179
transform 1 0 4968 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1649977179
transform 1 0 5888 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_57
timestamp 1649977179
transform 1 0 6348 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_69
timestamp 1649977179
transform 1 0 7452 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_73
timestamp 1649977179
transform 1 0 7820 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_103
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_107
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_111
timestamp 1649977179
transform 1 0 11316 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_115
timestamp 1649977179
transform 1 0 11684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_119
timestamp 1649977179
transform 1 0 12052 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_123
timestamp 1649977179
transform 1 0 12420 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1649977179
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1649977179
transform 1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_175
timestamp 1649977179
transform 1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_200
timestamp 1649977179
transform 1 0 19504 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_211
timestamp 1649977179
transform 1 0 20516 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1649977179
transform 1 0 20884 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_14
timestamp 1649977179
transform 1 0 2392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_25
timestamp 1649977179
transform 1 0 3404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_30
timestamp 1649977179
transform 1 0 3864 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_35
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_62
timestamp 1649977179
transform 1 0 6808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_74
timestamp 1649977179
transform 1 0 7912 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1649977179
transform 1 0 8280 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_103
timestamp 1649977179
transform 1 0 10580 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1649977179
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_135
timestamp 1649977179
transform 1 0 13524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 1649977179
transform 1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1649977179
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_148
timestamp 1649977179
transform 1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_171
timestamp 1649977179
transform 1 0 16836 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_175
timestamp 1649977179
transform 1 0 17204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_178
timestamp 1649977179
transform 1 0 17480 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1649977179
transform 1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1649977179
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_209
timestamp 1649977179
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1649977179
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_20
timestamp 1649977179
transform 1 0 2944 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1649977179
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1649977179
transform 1 0 4048 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_36
timestamp 1649977179
transform 1 0 4416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1649977179
transform 1 0 5612 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_60
timestamp 1649977179
transform 1 0 6624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_64
timestamp 1649977179
transform 1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_75
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_79
timestamp 1649977179
transform 1 0 8372 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_101
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_105
timestamp 1649977179
transform 1 0 10764 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_113
timestamp 1649977179
transform 1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_117
timestamp 1649977179
transform 1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1649977179
transform 1 0 12604 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_129
timestamp 1649977179
transform 1 0 12972 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1649977179
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1649977179
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_143
timestamp 1649977179
transform 1 0 14260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_147
timestamp 1649977179
transform 1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_151
timestamp 1649977179
transform 1 0 14996 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1649977179
transform 1 0 15272 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_158
timestamp 1649977179
transform 1 0 15640 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_176
timestamp 1649977179
transform 1 0 17296 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_199
timestamp 1649977179
transform 1 0 19412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_207
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_218
timestamp 1649977179
transform 1 0 21160 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_222
timestamp 1649977179
transform 1 0 21528 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1649977179
transform 1 0 2208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_17
timestamp 1649977179
transform 1 0 2668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_22
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_40
timestamp 1649977179
transform 1 0 4784 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1649977179
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_59
timestamp 1649977179
transform 1 0 6532 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_63
timestamp 1649977179
transform 1 0 6900 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1649977179
transform 1 0 7176 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_70
timestamp 1649977179
transform 1 0 7544 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 1649977179
transform 1 0 9568 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_115
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1649977179
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_122
timestamp 1649977179
transform 1 0 12328 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_140
timestamp 1649977179
transform 1 0 13984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1649977179
transform 1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_174
timestamp 1649977179
transform 1 0 17112 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_178
timestamp 1649977179
transform 1 0 17480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_182
timestamp 1649977179
transform 1 0 17848 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_186
timestamp 1649977179
transform 1 0 18216 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_190
timestamp 1649977179
transform 1 0 18584 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_194
timestamp 1649977179
transform 1 0 18952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_198
timestamp 1649977179
transform 1 0 19320 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_216
timestamp 1649977179
transform 1 0 20976 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_13
timestamp 1649977179
transform 1 0 2300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_18
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_22
timestamp 1649977179
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_38
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_42
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_48
timestamp 1649977179
transform 1 0 5520 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1649977179
transform 1 0 6624 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 1649977179
transform 1 0 7636 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_75
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1649977179
transform 1 0 12144 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_176
timestamp 1649977179
transform 1 0 17296 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1649977179
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_12
timestamp 1649977179
transform 1 0 2208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1649977179
transform 1 0 3220 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_31
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1649977179
transform 1 0 6808 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_73
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_77
timestamp 1649977179
transform 1 0 8188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_85
timestamp 1649977179
transform 1 0 8924 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_89
timestamp 1649977179
transform 1 0 9292 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1649977179
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_119
timestamp 1649977179
transform 1 0 12052 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_123
timestamp 1649977179
transform 1 0 12420 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_126
timestamp 1649977179
transform 1 0 12696 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1649977179
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_171
timestamp 1649977179
transform 1 0 16836 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_175
timestamp 1649977179
transform 1 0 17204 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_178
timestamp 1649977179
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_197
timestamp 1649977179
transform 1 0 19228 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1649977179
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_20
timestamp 1649977179
transform 1 0 2944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1649977179
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_38
timestamp 1649977179
transform 1 0 4600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_51
timestamp 1649977179
transform 1 0 5796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_63
timestamp 1649977179
transform 1 0 6900 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_74
timestamp 1649977179
transform 1 0 7912 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1649977179
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_105
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_113
timestamp 1649977179
transform 1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_117
timestamp 1649977179
transform 1 0 11868 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1649977179
transform 1 0 12604 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1649977179
transform 1 0 12972 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_143
timestamp 1649977179
transform 1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_147
timestamp 1649977179
transform 1 0 14628 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_151
timestamp 1649977179
transform 1 0 14996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_155
timestamp 1649977179
transform 1 0 15364 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_172
timestamp 1649977179
transform 1 0 16928 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_176
timestamp 1649977179
transform 1 0 17296 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 1649977179
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1649977179
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 1649977179
transform 1 0 2300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_18
timestamp 1649977179
transform 1 0 2760 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_22
timestamp 1649977179
transform 1 0 3128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_33
timestamp 1649977179
transform 1 0 4140 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_37
timestamp 1649977179
transform 1 0 4508 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1649977179
transform 1 0 4784 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_44
timestamp 1649977179
transform 1 0 5152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_48
timestamp 1649977179
transform 1 0 5520 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_61
timestamp 1649977179
transform 1 0 6716 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_72
timestamp 1649977179
transform 1 0 7728 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_83
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_87
timestamp 1649977179
transform 1 0 9108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_91
timestamp 1649977179
transform 1 0 9476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_95
timestamp 1649977179
transform 1 0 9844 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_99
timestamp 1649977179
transform 1 0 10212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1649977179
transform 1 0 10580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1649977179
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_119
timestamp 1649977179
transform 1 0 12052 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1649977179
transform 1 0 12420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_127
timestamp 1649977179
transform 1 0 12788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1649977179
transform 1 0 13156 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_135
timestamp 1649977179
transform 1 0 13524 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_140
timestamp 1649977179
transform 1 0 13984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_144
timestamp 1649977179
transform 1 0 14352 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1649977179
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_152
timestamp 1649977179
transform 1 0 15088 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_157
timestamp 1649977179
transform 1 0 15548 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1649977179
transform 1 0 16008 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_171
timestamp 1649977179
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_176
timestamp 1649977179
transform 1 0 17296 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_180
timestamp 1649977179
transform 1 0 17664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_186
timestamp 1649977179
transform 1 0 18216 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_190
timestamp 1649977179
transform 1 0 18584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_195
timestamp 1649977179
transform 1 0 19044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_200
timestamp 1649977179
transform 1 0 19504 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_206
timestamp 1649977179
transform 1 0 20056 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_14
timestamp 1649977179
transform 1 0 2392 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_21
timestamp 1649977179
transform 1 0 3036 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1649977179
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_34
timestamp 1649977179
transform 1 0 4232 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_38
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_49
timestamp 1649977179
transform 1 0 5612 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1649977179
transform 1 0 6256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_60
timestamp 1649977179
transform 1 0 6624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1649977179
transform 1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_75
timestamp 1649977179
transform 1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1649977179
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_94
timestamp 1649977179
transform 1 0 9752 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1649977179
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1649977179
transform 1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_106
timestamp 1649977179
transform 1 0 10856 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_110
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_123
timestamp 1649977179
transform 1 0 12420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1649977179
transform 1 0 12788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_131
timestamp 1649977179
transform 1 0 13156 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_135
timestamp 1649977179
transform 1 0 13524 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_147
timestamp 1649977179
transform 1 0 14628 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_159
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_163
timestamp 1649977179
transform 1 0 16100 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1649977179
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_172
timestamp 1649977179
transform 1 0 16928 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1649977179
transform 1 0 17296 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_187
timestamp 1649977179
transform 1 0 18308 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1649977179
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_199
timestamp 1649977179
transform 1 0 19412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1649977179
transform 1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1649977179
transform 1 0 2116 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_22
timestamp 1649977179
transform 1 0 3128 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_33
timestamp 1649977179
transform 1 0 4140 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_37
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_43
timestamp 1649977179
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_66
timestamp 1649977179
transform 1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_79
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_83
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_94
timestamp 1649977179
transform 1 0 9752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_106
timestamp 1649977179
transform 1 0 10856 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1649977179
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_115
timestamp 1649977179
transform 1 0 11684 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_127
timestamp 1649977179
transform 1 0 12788 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1649977179
transform 1 0 13248 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 1649977179
transform 1 0 14260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_154
timestamp 1649977179
transform 1 0 15272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_171
timestamp 1649977179
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_175
timestamp 1649977179
transform 1 0 17204 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_185
timestamp 1649977179
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_198
timestamp 1649977179
transform 1 0 19320 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1649977179
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_13
timestamp 1649977179
transform 1 0 2300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_18
timestamp 1649977179
transform 1 0 2760 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp 1649977179
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_40
timestamp 1649977179
transform 1 0 4784 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_52
timestamp 1649977179
transform 1 0 5888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_57
timestamp 1649977179
transform 1 0 6348 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1649977179
transform 1 0 6900 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1649977179
transform 1 0 7268 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_71
timestamp 1649977179
transform 1 0 7636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_87
timestamp 1649977179
transform 1 0 9108 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_91
timestamp 1649977179
transform 1 0 9476 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1649977179
transform 1 0 10488 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_113
timestamp 1649977179
transform 1 0 11500 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_118
timestamp 1649977179
transform 1 0 11960 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_129
timestamp 1649977179
transform 1 0 12972 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_134
timestamp 1649977179
transform 1 0 13432 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1649977179
transform 1 0 14444 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1649977179
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_154
timestamp 1649977179
transform 1 0 15272 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_169
timestamp 1649977179
transform 1 0 16652 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1649977179
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_185
timestamp 1649977179
transform 1 0 18124 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_207
timestamp 1649977179
transform 1 0 20148 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1649977179
transform 1 0 20884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_12
timestamp 1649977179
transform 1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1649977179
transform 1 0 2668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_22
timestamp 1649977179
transform 1 0 3128 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_26
timestamp 1649977179
transform 1 0 3496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_30
timestamp 1649977179
transform 1 0 3864 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_34
timestamp 1649977179
transform 1 0 4232 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_44
timestamp 1649977179
transform 1 0 5152 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_48
timestamp 1649977179
transform 1 0 5520 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1649977179
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_67
timestamp 1649977179
transform 1 0 7268 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_80
timestamp 1649977179
transform 1 0 8464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_84
timestamp 1649977179
transform 1 0 8832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_88
timestamp 1649977179
transform 1 0 9200 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1649977179
transform 1 0 10396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1649977179
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1649977179
transform 1 0 12144 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_124
timestamp 1649977179
transform 1 0 12512 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_128
timestamp 1649977179
transform 1 0 12880 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_139
timestamp 1649977179
transform 1 0 13892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_150
timestamp 1649977179
transform 1 0 14904 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1649977179
transform 1 0 17480 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1649977179
transform 1 0 18676 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_195
timestamp 1649977179
transform 1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_200
timestamp 1649977179
transform 1 0 19504 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1649977179
transform 1 0 20424 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1649977179
transform 1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1649977179
transform 1 0 2668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_22
timestamp 1649977179
transform 1 0 3128 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1649977179
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_31
timestamp 1649977179
transform 1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_35
timestamp 1649977179
transform 1 0 4324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_46
timestamp 1649977179
transform 1 0 5336 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_50
timestamp 1649977179
transform 1 0 5704 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_54
timestamp 1649977179
transform 1 0 6072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_58
timestamp 1649977179
transform 1 0 6440 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_62
timestamp 1649977179
transform 1 0 6808 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_66
timestamp 1649977179
transform 1 0 7176 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_70
timestamp 1649977179
transform 1 0 7544 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_87
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_91
timestamp 1649977179
transform 1 0 9476 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_95 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9844 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_106
timestamp 1649977179
transform 1 0 10856 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_110
timestamp 1649977179
transform 1 0 11224 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_113
timestamp 1649977179
transform 1 0 11500 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_117
timestamp 1649977179
transform 1 0 11868 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_124
timestamp 1649977179
transform 1 0 12512 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_128
timestamp 1649977179
transform 1 0 12880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_132
timestamp 1649977179
transform 1 0 13248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_146
timestamp 1649977179
transform 1 0 14536 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_157
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1649977179
transform 1 0 16100 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_167
timestamp 1649977179
transform 1 0 16468 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_174
timestamp 1649977179
transform 1 0 17112 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_179
timestamp 1649977179
transform 1 0 17572 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_184
timestamp 1649977179
transform 1 0 18032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_203
timestamp 1649977179
transform 1 0 19780 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_208
timestamp 1649977179
transform 1 0 20240 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_18
timestamp 1649977179
transform 1 0 2760 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_22
timestamp 1649977179
transform 1 0 3128 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_32
timestamp 1649977179
transform 1 0 4048 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1649977179
transform 1 0 4416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_40
timestamp 1649977179
transform 1 0 4784 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1649977179
transform 1 0 6808 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_73
timestamp 1649977179
transform 1 0 7820 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1649977179
transform 1 0 8188 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_82
timestamp 1649977179
transform 1 0 8648 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_86
timestamp 1649977179
transform 1 0 9016 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_90
timestamp 1649977179
transform 1 0 9384 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_94
timestamp 1649977179
transform 1 0 9752 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_97
timestamp 1649977179
transform 1 0 10028 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_122
timestamp 1649977179
transform 1 0 12328 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_127
timestamp 1649977179
transform 1 0 12788 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_143
timestamp 1649977179
transform 1 0 14260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_147
timestamp 1649977179
transform 1 0 14628 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_158
timestamp 1649977179
transform 1 0 15640 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1649977179
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_178
timestamp 1649977179
transform 1 0 17480 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_191
timestamp 1649977179
transform 1 0 18676 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_195
timestamp 1649977179
transform 1 0 19044 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1649977179
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_210
timestamp 1649977179
transform 1 0 20424 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1649977179
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_18
timestamp 1649977179
transform 1 0 2760 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1649977179
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_38
timestamp 1649977179
transform 1 0 4600 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_43
timestamp 1649977179
transform 1 0 5060 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_50
timestamp 1649977179
transform 1 0 5704 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_54
timestamp 1649977179
transform 1 0 6072 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_58
timestamp 1649977179
transform 1 0 6440 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_63
timestamp 1649977179
transform 1 0 6900 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_67
timestamp 1649977179
transform 1 0 7268 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1649977179
transform 1 0 7636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_88
timestamp 1649977179
transform 1 0 9200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1649977179
transform 1 0 9660 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_104
timestamp 1649977179
transform 1 0 10672 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_115
timestamp 1649977179
transform 1 0 11684 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_127
timestamp 1649977179
transform 1 0 12788 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1649977179
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1649977179
transform 1 0 14352 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1649977179
transform 1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_160
timestamp 1649977179
transform 1 0 15824 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1649977179
transform 1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_182
timestamp 1649977179
transform 1 0 17848 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_187
timestamp 1649977179
transform 1 0 18308 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1649977179
transform 1 0 20056 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_210
timestamp 1649977179
transform 1 0 20424 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1649977179
transform 1 0 20884 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1649977179
transform 1 0 1748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1649977179
transform 1 0 2300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_18
timestamp 1649977179
transform 1 0 2760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_23
timestamp 1649977179
transform 1 0 3220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_31
timestamp 1649977179
transform 1 0 3956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_35
timestamp 1649977179
transform 1 0 4324 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_43
timestamp 1649977179
transform 1 0 5060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_47
timestamp 1649977179
transform 1 0 5428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_67
timestamp 1649977179
transform 1 0 7268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp 1649977179
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_83
timestamp 1649977179
transform 1 0 8740 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_90
timestamp 1649977179
transform 1 0 9384 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_101
timestamp 1649977179
transform 1 0 10396 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_106
timestamp 1649977179
transform 1 0 10856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_118
timestamp 1649977179
transform 1 0 11960 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_122
timestamp 1649977179
transform 1 0 12328 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_129
timestamp 1649977179
transform 1 0 12972 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_133
timestamp 1649977179
transform 1 0 13340 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_146
timestamp 1649977179
transform 1 0 14536 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_151
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1649977179
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_159
timestamp 1649977179
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1649977179
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_172
timestamp 1649977179
transform 1 0 16928 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_180
timestamp 1649977179
transform 1 0 17664 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_184
timestamp 1649977179
transform 1 0 18032 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_189
timestamp 1649977179
transform 1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _056_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18676 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1649977179
transform 1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1649977179
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1649977179
transform 1 0 2760 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1649977179
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 2392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform 1 0 2852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 2944 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 2392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 2852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 2944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform 1 0 20608 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform -1 0 19504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform -1 0 19964 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform -1 0 20332 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform 1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform -1 0 19228 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 19044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform -1 0 20424 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform -1 0 18032 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 15272 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 16376 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 18952 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 17572 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 19504 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 12788 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 18952 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 16928 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 17112 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 4324 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform -1 0 3404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 8648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 15272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 10212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 16192 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform 1 0 21160 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform -1 0 15456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform -1 0 5244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform -1 0 5428 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform -1 0 5796 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform 1 0 3772 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1649977179
transform 1 0 2668 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1649977179
transform -1 0 2300 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 3496 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1649977179
transform -1 0 2300 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 1932 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 3128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform 1 0 2576 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1649977179
transform -1 0 2300 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1649977179
transform -1 0 2300 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform 1 0 20516 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 19320 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1649977179
transform 1 0 20516 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 21436 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 18952 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1649977179
transform -1 0 21436 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1649977179
transform 1 0 20516 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 21160 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 18768 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1649977179
transform 1 0 20516 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform -1 0 21436 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform -1 0 21436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform -1 0 18952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 21436 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform -1 0 21436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform -1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1649977179
transform 1 0 9200 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform -1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform 1 0 10764 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform 1 0 12328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform -1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform -1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform -1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1649977179
transform -1 0 6072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1649977179
transform -1 0 8004 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1649977179
transform -1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform -1 0 8004 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1649977179
transform -1 0 6072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1649977179
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1649977179
transform 1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1649977179
transform 1 0 3128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1649977179
transform 1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1649977179
transform -1 0 2300 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1649977179
transform -1 0 3220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1649977179
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1649977179
transform -1 0 17572 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1649977179
transform -1 0 13800 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1649977179
transform -1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1649977179
transform 1 0 14720 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1649977179
transform -1 0 16376 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1649977179
transform -1 0 16376 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1649977179
transform -1 0 18676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1649977179
transform -1 0 16376 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  mem_bottom_track_1.delay_buf_2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12788 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14628 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14720 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_bottom_track_3.delay_buf_2
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16376 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13156 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10488 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_bottom_track_5.delay_buf_2
timestamp 1649977179
transform -1 0 5612 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10948 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13432 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10580 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_bottom_track_7.delay_buf_2
timestamp 1649977179
transform 1 0 7820 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12696 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10580 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10856 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13984 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9016 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10764 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10580 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9200 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10764 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9384 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9752 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14352 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16928 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14812 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17296 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 17296 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14904 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15640 0 1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 19780 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10672 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13616 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12512 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10488 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11868 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10948 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10580 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15640 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 12144 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_left_track_17.delay_buf_2
timestamp 1649977179
transform -1 0 5888 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16100 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14444 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_left_track_25.delay_buf_2
timestamp 1649977179
transform -1 0 11500 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14720 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13708 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10764 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16376 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13248 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_right_track_0.delay_buf
timestamp 1649977179
transform 1 0 11960 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14628 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18216 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17480 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20424 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18952 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17020 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 20792 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17572 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 20976 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 20884 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_right_track_16.delay_buf_2
timestamp 1649977179
transform -1 0 17480 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19228 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13892 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  mem_right_track_24.delay_buf_2
timestamp 1649977179
transform -1 0 12420 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18308 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21068 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3312 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2116 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l1_in_3__172 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2300 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2484 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3312 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4968 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1649977179
transform -1 0 5520 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l1_in_3__182
timestamp 1649977179
transform 1 0 6532 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6164 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6440 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5980 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5152 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform -1 0 5612 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2576 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l1_in_3__155
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4416 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4968 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_7.mux_l1_in_3__156
timestamp 1649977179
transform 1 0 6624 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1649977179
transform 1 0 5612 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5060 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5704 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6072 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7728 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8740 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_1__157
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8648 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9660 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_11.mux_l2_in_1__173
timestamp 1649977179
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8648 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10396 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_13.mux_l1_in_1__174
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7360 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7728 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_15.mux_l1_in_1__175
timestamp 1649977179
transform 1 0 6072 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1649977179
transform -1 0 5888 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7452 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7176 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l1_in_1__176
timestamp 1649977179
transform -1 0 5060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 5612 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7636 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10396 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_19.mux_l1_in_1__177
timestamp 1649977179
transform 1 0 13156 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12144 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10856 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_21.mux_l1_in_1__178
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13800 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14260 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10672 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_23.mux_l1_in_1__179
timestamp 1649977179
transform 1 0 13432 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13064 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11684 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17664 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_1__180
timestamp 1649977179
transform 1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16284 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16652 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20056 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_27.mux_l2_in_0__181
timestamp 1649977179
transform -1 0 16376 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17020 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7084 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4968 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4508 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_3__158
timestamp 1649977179
transform 1 0 6072 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3956 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4232 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4600 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6440 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7360 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3128 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2760 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_3__161
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5060 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2668 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2484 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform -1 0 3220 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1649977179
transform 1 0 1564 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1649977179
transform 1 0 1656 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3312 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 2392 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_3__163
timestamp 1649977179
transform 1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 1656 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 1564 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2392 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7636 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4048 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l2_in_3__164
timestamp 1649977179
transform 1 0 4784 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4600 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6440 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5152 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l1_in_3__159
timestamp 1649977179
transform 1 0 3312 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1649977179
transform -1 0 3496 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2300 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6992 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6900 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l1_in_3__160
timestamp 1649977179
transform 1 0 5244 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4784 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6256 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 3404 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l2_in_1__162
timestamp 1649977179
transform 1 0 5428 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4968 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4508 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2760 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20608 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20516 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 20240 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19780 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19688 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3404 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_3__165
timestamp 1649977179
transform 1 0 18216 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17848 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19504 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 17756 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 18124 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18768 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8280 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8648 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1649977179
transform -1 0 11040 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_3__167
timestamp 1649977179
transform 1 0 10580 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15088 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13248 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 18124 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20056 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 19872 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 20608 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1649977179
transform -1 0 20332 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1649977179
transform 1 0 20240 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1649977179
transform -1 0 13984 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1649977179
transform 1 0 20608 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20424 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 20332 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1649977179
transform -1 0 17664 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_3__170
timestamp 1649977179
transform -1 0 19504 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 20240 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19596 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 18308 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 19320 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20424 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20424 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8372 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 7820 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l2_in_3__171
timestamp 1649977179
transform -1 0 14628 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19320 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 14904 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 18676 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19780 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11592 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8096 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15732 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l1_in_3__166
timestamp 1649977179
transform 1 0 15456 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1649977179
transform -1 0 15824 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12328 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15088 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13892 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18216 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15548 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1649977179
transform 1 0 16008 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l1_in_3__168
timestamp 1649977179
transform -1 0 16100 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16652 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15640 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10304 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16376 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l2_in_1__169
timestamp 1649977179
transform -1 0 18952 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 20056 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19504 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output89 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 17296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 2300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform -1 0 2300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform -1 0 2300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform -1 0 20148 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 21068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform 1 0 20516 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform 1 0 21068 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 20516 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 19964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform 1 0 19688 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 20516 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1649977179
transform 1 0 17204 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform -1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform 1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform 1 0 19596 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  repeater151
timestamp 1649977179
transform -1 0 21436 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater152
timestamp 1649977179
transform 1 0 17756 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater153
timestamp 1649977179
transform -1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater154
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 406 592
<< labels >>
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 0 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 1 nsew signal tristate
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_42_
port 4 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_43_
port 5 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_44_
port 6 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_45_
port 7 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_46_
port 8 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_47_
port 9 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_48_
port 10 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_49_
port 11 nsew signal input
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 ccff_head
port 12 nsew signal input
flabel metal2 s 17222 22200 17278 23000 0 FreeSans 224 90 0 0 ccff_tail
port 13 nsew signal tristate
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 14 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 15 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 16 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 17 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 18 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 19 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 20 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 21 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 22 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 23 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 24 nsew signal input
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 25 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 26 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 27 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 28 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 29 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 30 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 31 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 32 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 33 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 34 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 35 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 36 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 37 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 38 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 39 nsew signal tristate
flabel metal3 s 0 19184 800 19304 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 40 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 41 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 42 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 43 nsew signal tristate
flabel metal3 s 0 20816 800 20936 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 44 nsew signal tristate
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 45 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 46 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 47 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 48 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 49 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 50 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 51 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 52 nsew signal tristate
flabel metal3 s 0 16736 800 16856 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 53 nsew signal tristate
flabel metal3 s 22200 4904 23000 5024 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 54 nsew signal input
flabel metal3 s 22200 8984 23000 9104 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 55 nsew signal input
flabel metal3 s 22200 9392 23000 9512 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 56 nsew signal input
flabel metal3 s 22200 9800 23000 9920 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 57 nsew signal input
flabel metal3 s 22200 10208 23000 10328 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 58 nsew signal input
flabel metal3 s 22200 10616 23000 10736 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 59 nsew signal input
flabel metal3 s 22200 11024 23000 11144 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 60 nsew signal input
flabel metal3 s 22200 11432 23000 11552 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 61 nsew signal input
flabel metal3 s 22200 11840 23000 11960 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 62 nsew signal input
flabel metal3 s 22200 12248 23000 12368 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 63 nsew signal input
flabel metal3 s 22200 12656 23000 12776 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 64 nsew signal input
flabel metal3 s 22200 5312 23000 5432 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 65 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 66 nsew signal input
flabel metal3 s 22200 6128 23000 6248 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 67 nsew signal input
flabel metal3 s 22200 6536 23000 6656 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 68 nsew signal input
flabel metal3 s 22200 6944 23000 7064 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 69 nsew signal input
flabel metal3 s 22200 7352 23000 7472 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 70 nsew signal input
flabel metal3 s 22200 7760 23000 7880 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 71 nsew signal input
flabel metal3 s 22200 8168 23000 8288 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 72 nsew signal input
flabel metal3 s 22200 8576 23000 8696 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 73 nsew signal input
flabel metal3 s 22200 13064 23000 13184 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 74 nsew signal tristate
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 75 nsew signal tristate
flabel metal3 s 22200 17552 23000 17672 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 76 nsew signal tristate
flabel metal3 s 22200 17960 23000 18080 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 77 nsew signal tristate
flabel metal3 s 22200 18368 23000 18488 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 78 nsew signal tristate
flabel metal3 s 22200 18776 23000 18896 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 79 nsew signal tristate
flabel metal3 s 22200 19184 23000 19304 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 80 nsew signal tristate
flabel metal3 s 22200 19592 23000 19712 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 81 nsew signal tristate
flabel metal3 s 22200 20000 23000 20120 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 82 nsew signal tristate
flabel metal3 s 22200 20408 23000 20528 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 83 nsew signal tristate
flabel metal3 s 22200 20816 23000 20936 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 84 nsew signal tristate
flabel metal3 s 22200 13472 23000 13592 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 85 nsew signal tristate
flabel metal3 s 22200 13880 23000 14000 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 86 nsew signal tristate
flabel metal3 s 22200 14288 23000 14408 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 87 nsew signal tristate
flabel metal3 s 22200 14696 23000 14816 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 88 nsew signal tristate
flabel metal3 s 22200 15104 23000 15224 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 89 nsew signal tristate
flabel metal3 s 22200 15512 23000 15632 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 90 nsew signal tristate
flabel metal3 s 22200 15920 23000 16040 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 91 nsew signal tristate
flabel metal3 s 22200 16328 23000 16448 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 92 nsew signal tristate
flabel metal3 s 22200 16736 23000 16856 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 93 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 94 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 95 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 96 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 97 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 98 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 99 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 100 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 101 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 102 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 103 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 104 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 105 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 106 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 107 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 108 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 109 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 110 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 111 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 112 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 113 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 114 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 115 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 116 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 117 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 118 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 119 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 120 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 121 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 122 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 123 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 124 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 125 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 126 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 127 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 128 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 129 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 130 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 131 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 132 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 133 nsew signal tristate
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 left_bottom_grid_pin_34_
port 134 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 left_bottom_grid_pin_35_
port 135 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 left_bottom_grid_pin_36_
port 136 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 left_bottom_grid_pin_37_
port 137 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_bottom_grid_pin_38_
port 138 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_bottom_grid_pin_39_
port 139 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 left_bottom_grid_pin_40_
port 140 nsew signal input
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 left_bottom_grid_pin_41_
port 141 nsew signal input
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 left_top_grid_pin_1_
port 142 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 prog_clk_0_S_in
port 143 nsew signal input
flabel metal3 s 22200 1640 23000 1760 0 FreeSans 480 0 0 0 right_bottom_grid_pin_34_
port 144 nsew signal input
flabel metal3 s 22200 2048 23000 2168 0 FreeSans 480 0 0 0 right_bottom_grid_pin_35_
port 145 nsew signal input
flabel metal3 s 22200 2456 23000 2576 0 FreeSans 480 0 0 0 right_bottom_grid_pin_36_
port 146 nsew signal input
flabel metal3 s 22200 2864 23000 2984 0 FreeSans 480 0 0 0 right_bottom_grid_pin_37_
port 147 nsew signal input
flabel metal3 s 22200 3272 23000 3392 0 FreeSans 480 0 0 0 right_bottom_grid_pin_38_
port 148 nsew signal input
flabel metal3 s 22200 3680 23000 3800 0 FreeSans 480 0 0 0 right_bottom_grid_pin_39_
port 149 nsew signal input
flabel metal3 s 22200 4088 23000 4208 0 FreeSans 480 0 0 0 right_bottom_grid_pin_40_
port 150 nsew signal input
flabel metal3 s 22200 4496 23000 4616 0 FreeSans 480 0 0 0 right_bottom_grid_pin_41_
port 151 nsew signal input
flabel metal3 s 22200 21224 23000 21344 0 FreeSans 480 0 0 0 right_top_grid_pin_1_
port 152 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
