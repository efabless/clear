magic
tech sky130A
magscale 1 2
timestamp 1625786300
<< locali >>
rect 11713 21335 11747 21505
rect 23581 19363 23615 20213
rect 17049 14875 17083 15113
rect 23581 13855 23615 14773
rect 17785 13719 17819 13821
rect 16497 11543 16531 11781
rect 14289 10455 14323 10557
rect 16497 10455 16531 10761
rect 11713 9435 11747 9605
rect 13645 9435 13679 9605
rect 13921 7735 13955 7973
rect 23581 3043 23615 3893
rect 23581 1411 23615 2329
<< viali >>
rect 3709 22185 3743 22219
rect 5181 22185 5215 22219
rect 7849 22185 7883 22219
rect 8217 22185 8251 22219
rect 8493 22185 8527 22219
rect 12173 22185 12207 22219
rect 15669 22185 15703 22219
rect 18889 22185 18923 22219
rect 4077 22117 4111 22151
rect 4445 22117 4479 22151
rect 5641 22117 5675 22151
rect 10793 22117 10827 22151
rect 13737 22117 13771 22151
rect 15577 22117 15611 22151
rect 17417 22117 17451 22151
rect 17923 22117 17957 22151
rect 20453 22117 20487 22151
rect 22201 22117 22235 22151
rect 22937 22117 22971 22151
rect 1409 22049 1443 22083
rect 1593 22049 1627 22083
rect 1961 22049 1995 22083
rect 2329 22049 2363 22083
rect 2697 22049 2731 22083
rect 2881 22049 2915 22083
rect 3065 22049 3099 22083
rect 3525 22049 3559 22083
rect 4261 22049 4295 22083
rect 4813 22049 4847 22083
rect 4997 22049 5031 22083
rect 5365 22049 5399 22083
rect 6001 22049 6035 22083
rect 6093 22049 6127 22083
rect 6745 22049 6779 22083
rect 7021 22049 7055 22083
rect 7389 22049 7423 22083
rect 8677 22049 8711 22083
rect 9229 22049 9263 22083
rect 9873 22049 9907 22083
rect 10057 22049 10091 22083
rect 11621 22049 11655 22083
rect 12081 22049 12115 22083
rect 12357 22049 12391 22083
rect 12725 22049 12759 22083
rect 12817 22049 12851 22083
rect 13093 22049 13127 22083
rect 14381 22049 14415 22083
rect 14565 22049 14599 22083
rect 15025 22049 15059 22083
rect 15393 22049 15427 22083
rect 15853 22049 15887 22083
rect 16129 22049 16163 22083
rect 16497 22049 16531 22083
rect 16589 22049 16623 22083
rect 17049 22049 17083 22083
rect 17233 22049 17267 22083
rect 18061 22049 18095 22083
rect 18705 22049 18739 22083
rect 19165 22049 19199 22083
rect 19533 22049 19567 22083
rect 19901 22049 19935 22083
rect 20085 22049 20119 22083
rect 20269 22049 20303 22083
rect 20821 22049 20855 22083
rect 20913 22049 20947 22083
rect 21097 22049 21131 22083
rect 21465 22049 21499 22083
rect 21649 22049 21683 22083
rect 21833 22049 21867 22083
rect 23121 22049 23155 22083
rect 1777 21981 1811 22015
rect 2513 21981 2547 22015
rect 7573 21981 7607 22015
rect 7757 21981 7791 22015
rect 8401 21981 8435 22015
rect 8971 21981 9005 22015
rect 9781 21981 9815 22015
rect 10517 21981 10551 22015
rect 10701 21981 10735 22015
rect 10885 21981 10919 22015
rect 13829 21981 13863 22015
rect 13921 21981 13955 22015
rect 18153 21981 18187 22015
rect 19717 21981 19751 22015
rect 22385 21981 22419 22015
rect 2145 21913 2179 21947
rect 3893 21913 3927 21947
rect 4721 21913 4755 21947
rect 5825 21913 5859 21947
rect 11437 21913 11471 21947
rect 13369 21913 13403 21947
rect 14841 21913 14875 21947
rect 18521 21913 18555 21947
rect 19349 21913 19383 21947
rect 3341 21845 3375 21879
rect 5549 21845 5583 21879
rect 6285 21845 6319 21879
rect 6561 21845 6595 21879
rect 6837 21845 6871 21879
rect 7205 21845 7239 21879
rect 11253 21845 11287 21879
rect 11897 21845 11931 21879
rect 12541 21845 12575 21879
rect 13001 21845 13035 21879
rect 13277 21845 13311 21879
rect 14197 21845 14231 21879
rect 14749 21845 14783 21879
rect 15209 21845 15243 21879
rect 15945 21845 15979 21879
rect 16773 21845 16807 21879
rect 16865 21845 16899 21879
rect 20637 21845 20671 21879
rect 21925 21845 21959 21879
rect 1869 21641 1903 21675
rect 2145 21641 2179 21675
rect 4077 21641 4111 21675
rect 6469 21641 6503 21675
rect 6745 21641 6779 21675
rect 6929 21641 6963 21675
rect 9229 21641 9263 21675
rect 9413 21641 9447 21675
rect 10977 21641 11011 21675
rect 16129 21641 16163 21675
rect 16773 21641 16807 21675
rect 19441 21641 19475 21675
rect 2513 21573 2547 21607
rect 3985 21573 4019 21607
rect 11345 21573 11379 21607
rect 14657 21573 14691 21607
rect 16221 21573 16255 21607
rect 19717 21573 19751 21607
rect 22753 21573 22787 21607
rect 5917 21505 5951 21539
rect 8309 21505 8343 21539
rect 10793 21505 10827 21539
rect 11713 21505 11747 21539
rect 11805 21505 11839 21539
rect 18797 21505 18831 21539
rect 19901 21505 19935 21539
rect 23121 21505 23155 21539
rect 1593 21437 1627 21471
rect 1685 21437 1719 21471
rect 2053 21437 2087 21471
rect 2329 21437 2363 21471
rect 2605 21437 2639 21471
rect 4261 21437 4295 21471
rect 4445 21437 4479 21471
rect 6653 21437 6687 21471
rect 8053 21437 8087 21471
rect 8493 21437 8527 21471
rect 11061 21437 11095 21471
rect 11529 21437 11563 21471
rect 2872 21369 2906 21403
rect 4712 21369 4746 21403
rect 6101 21369 6135 21403
rect 6285 21369 6319 21403
rect 8953 21369 8987 21403
rect 10548 21369 10582 21403
rect 13277 21437 13311 21471
rect 14749 21437 14783 21471
rect 16405 21437 16439 21471
rect 16957 21437 16991 21471
rect 18521 21437 18555 21471
rect 20085 21437 20119 21471
rect 22937 21437 22971 21471
rect 12072 21369 12106 21403
rect 13522 21369 13556 21403
rect 14994 21369 15028 21403
rect 16497 21369 16531 21403
rect 17224 21369 17258 21403
rect 19349 21369 19383 21403
rect 22569 21369 22603 21403
rect 5825 21301 5859 21335
rect 11253 21301 11287 21335
rect 11713 21301 11747 21335
rect 13185 21301 13219 21335
rect 18337 21301 18371 21335
rect 20729 21301 20763 21335
rect 21373 21301 21407 21335
rect 21925 21301 21959 21335
rect 22201 21301 22235 21335
rect 1961 21097 1995 21131
rect 3525 21097 3559 21131
rect 5273 21097 5307 21131
rect 8309 21097 8343 21131
rect 8585 21097 8619 21131
rect 9137 21097 9171 21131
rect 10793 21097 10827 21131
rect 11069 21097 11103 21131
rect 11529 21097 11563 21131
rect 13369 21097 13403 21131
rect 13737 21097 13771 21131
rect 13921 21097 13955 21131
rect 15761 21097 15795 21131
rect 18797 21097 18831 21131
rect 19073 21097 19107 21131
rect 19625 21097 19659 21131
rect 21189 21097 21223 21131
rect 21741 21097 21775 21131
rect 22293 21097 22327 21131
rect 1501 21029 1535 21063
rect 4160 21029 4194 21063
rect 5632 21029 5666 21063
rect 9588 21029 9622 21063
rect 11345 21029 11379 21063
rect 13277 21029 13311 21063
rect 14013 21029 14047 21063
rect 14648 21029 14682 21063
rect 16120 21029 16154 21063
rect 22569 21029 22603 21063
rect 1777 20961 1811 20995
rect 2053 20961 2087 20995
rect 2320 20961 2354 20995
rect 3709 20961 3743 20995
rect 3893 20961 3927 20995
rect 5365 20961 5399 20995
rect 7093 20961 7127 20995
rect 8493 20961 8527 20995
rect 8769 20961 8803 20995
rect 12642 20961 12676 20995
rect 12909 20961 12943 20995
rect 17592 20961 17626 20995
rect 19257 20961 19291 20995
rect 19349 20961 19383 20995
rect 20729 20961 20763 20995
rect 21005 20961 21039 20995
rect 21281 20961 21315 20995
rect 21557 20961 21591 20995
rect 21833 20961 21867 20995
rect 22201 20961 22235 20995
rect 22937 20961 22971 20995
rect 6837 20893 6871 20927
rect 8861 20893 8895 20927
rect 9321 20893 9355 20927
rect 13185 20893 13219 20927
rect 14381 20893 14415 20927
rect 15853 20893 15887 20927
rect 17325 20893 17359 20927
rect 1685 20825 1719 20859
rect 3433 20825 3467 20859
rect 20821 20825 20855 20859
rect 21465 20825 21499 20859
rect 22017 20825 22051 20859
rect 22753 20825 22787 20859
rect 6745 20757 6779 20791
rect 8217 20757 8251 20791
rect 10701 20757 10735 20791
rect 17233 20757 17267 20791
rect 18705 20757 18739 20791
rect 23029 20757 23063 20791
rect 2973 20553 3007 20587
rect 7021 20553 7055 20587
rect 8677 20553 8711 20587
rect 9229 20553 9263 20587
rect 11345 20553 11379 20587
rect 13185 20553 13219 20587
rect 13921 20553 13955 20587
rect 16681 20553 16715 20587
rect 17325 20553 17359 20587
rect 19625 20553 19659 20587
rect 21741 20553 21775 20587
rect 22017 20553 22051 20587
rect 20729 20485 20763 20519
rect 3249 20417 3283 20451
rect 4077 20417 4111 20451
rect 4905 20417 4939 20451
rect 5733 20417 5767 20451
rect 7205 20417 7239 20451
rect 10885 20417 10919 20451
rect 14473 20417 14507 20451
rect 14841 20417 14875 20451
rect 15761 20417 15795 20451
rect 18889 20417 18923 20451
rect 20177 20417 20211 20451
rect 1593 20349 1627 20383
rect 3433 20349 3467 20383
rect 4261 20349 4295 20383
rect 6929 20349 6963 20383
rect 7472 20349 7506 20383
rect 8861 20349 8895 20383
rect 10609 20349 10643 20383
rect 13093 20349 13127 20383
rect 13369 20349 13403 20383
rect 14289 20349 14323 20383
rect 14381 20349 14415 20383
rect 15853 20349 15887 20383
rect 16589 20349 16623 20383
rect 17141 20349 17175 20383
rect 18705 20349 18739 20383
rect 21005 20349 21039 20383
rect 21281 20349 21315 20383
rect 21557 20349 21591 20383
rect 21833 20349 21867 20383
rect 22477 20349 22511 20383
rect 1860 20281 1894 20315
rect 3341 20281 3375 20315
rect 4997 20281 5031 20315
rect 5825 20281 5859 20315
rect 9137 20281 9171 20315
rect 10342 20281 10376 20315
rect 10793 20281 10827 20315
rect 12826 20281 12860 20315
rect 13645 20281 13679 20315
rect 15117 20281 15151 20315
rect 15945 20281 15979 20315
rect 18438 20281 18472 20315
rect 19165 20281 19199 20315
rect 19993 20281 20027 20315
rect 22845 20281 22879 20315
rect 3801 20213 3835 20247
rect 4169 20213 4203 20247
rect 4629 20213 4663 20247
rect 5089 20213 5123 20247
rect 5457 20213 5491 20247
rect 5917 20213 5951 20247
rect 6285 20213 6319 20247
rect 6653 20213 6687 20247
rect 6745 20213 6779 20247
rect 8585 20213 8619 20247
rect 10885 20213 10919 20247
rect 11713 20213 11747 20247
rect 15025 20213 15059 20247
rect 15485 20213 15519 20247
rect 16313 20213 16347 20247
rect 16405 20213 16439 20247
rect 19073 20213 19107 20247
rect 19533 20213 19567 20247
rect 20085 20213 20119 20247
rect 20453 20213 20487 20247
rect 20913 20213 20947 20247
rect 21189 20213 21223 20247
rect 21465 20213 21499 20247
rect 22293 20213 22327 20247
rect 23581 20213 23615 20247
rect 1593 20009 1627 20043
rect 3709 20009 3743 20043
rect 3893 20009 3927 20043
rect 4261 20009 4295 20043
rect 5457 20009 5491 20043
rect 5825 20009 5859 20043
rect 6377 20009 6411 20043
rect 7113 20009 7147 20043
rect 8769 20009 8803 20043
rect 11161 20009 11195 20043
rect 11989 20009 12023 20043
rect 12449 20009 12483 20043
rect 12909 20009 12943 20043
rect 13277 20009 13311 20043
rect 13737 20009 13771 20043
rect 15301 20009 15335 20043
rect 15945 20009 15979 20043
rect 16405 20009 16439 20043
rect 16773 20009 16807 20043
rect 22661 20009 22695 20043
rect 4353 19941 4387 19975
rect 5917 19941 5951 19975
rect 8248 19941 8282 19975
rect 9934 19941 9968 19975
rect 14749 19941 14783 19975
rect 15577 19941 15611 19975
rect 16313 19941 16347 19975
rect 17325 19941 17359 19975
rect 18714 19941 18748 19975
rect 22937 19941 22971 19975
rect 2717 19873 2751 19907
rect 3249 19873 3283 19907
rect 3525 19873 3559 19907
rect 5089 19873 5123 19907
rect 6561 19873 6595 19907
rect 11529 19873 11563 19907
rect 12265 19873 12299 19907
rect 14841 19873 14875 19907
rect 15485 19873 15519 19907
rect 15761 19873 15795 19907
rect 16865 19873 16899 19907
rect 19993 19873 20027 19907
rect 20729 19873 20763 19907
rect 21272 19873 21306 19907
rect 22477 19873 22511 19907
rect 2973 19805 3007 19839
rect 4537 19805 4571 19839
rect 4905 19805 4939 19839
rect 4997 19805 5031 19839
rect 5733 19805 5767 19839
rect 8493 19805 8527 19839
rect 9689 19805 9723 19839
rect 11621 19805 11655 19839
rect 11713 19805 11747 19839
rect 12725 19805 12759 19839
rect 12817 19805 12851 19839
rect 13553 19805 13587 19839
rect 13645 19805 13679 19839
rect 14657 19805 14691 19839
rect 16129 19805 16163 19839
rect 18981 19805 19015 19839
rect 19809 19805 19843 19839
rect 19901 19805 19935 19839
rect 21005 19805 21039 19839
rect 3433 19737 3467 19771
rect 6285 19737 6319 19771
rect 14105 19737 14139 19771
rect 17141 19737 17175 19771
rect 20913 19737 20947 19771
rect 23121 19737 23155 19771
rect 3157 19669 3191 19703
rect 6745 19669 6779 19703
rect 9229 19669 9263 19703
rect 11069 19669 11103 19703
rect 15209 19669 15243 19703
rect 17049 19669 17083 19703
rect 17601 19669 17635 19703
rect 20361 19669 20395 19703
rect 20637 19669 20671 19703
rect 22385 19669 22419 19703
rect 3985 19465 4019 19499
rect 5825 19465 5859 19499
rect 9321 19465 9355 19499
rect 11529 19465 11563 19499
rect 13093 19465 13127 19499
rect 19809 19465 19843 19499
rect 21557 19465 21591 19499
rect 3341 19329 3375 19363
rect 4629 19329 4663 19363
rect 5457 19329 5491 19363
rect 6561 19329 6595 19363
rect 6745 19329 6779 19363
rect 7944 19329 7978 19363
rect 10241 19329 10275 19363
rect 10609 19329 10643 19363
rect 13277 19329 13311 19363
rect 14105 19329 14139 19363
rect 15393 19329 15427 19363
rect 16221 19329 16255 19363
rect 19257 19329 19291 19363
rect 22017 19329 22051 19363
rect 22845 19329 22879 19363
rect 23581 19329 23615 19363
rect 1685 19261 1719 19295
rect 5641 19261 5675 19295
rect 5917 19261 5951 19295
rect 6837 19261 6871 19295
rect 7481 19261 7515 19295
rect 8217 19261 8251 19295
rect 11345 19261 11379 19295
rect 11713 19261 11747 19295
rect 14381 19261 14415 19295
rect 18070 19261 18104 19295
rect 18337 19261 18371 19295
rect 19901 19261 19935 19295
rect 21373 19261 21407 19295
rect 21833 19261 21867 19295
rect 22569 19261 22603 19295
rect 1952 19193 1986 19227
rect 3525 19193 3559 19227
rect 4445 19193 4479 19227
rect 5181 19193 5215 19227
rect 10057 19193 10091 19227
rect 11980 19193 12014 19227
rect 13553 19193 13587 19227
rect 14289 19193 14323 19227
rect 20168 19193 20202 19227
rect 21649 19193 21683 19227
rect 22661 19193 22695 19227
rect 3065 19125 3099 19159
rect 3433 19125 3467 19159
rect 3893 19125 3927 19159
rect 4353 19125 4387 19159
rect 4813 19125 4847 19159
rect 5273 19125 5307 19159
rect 6101 19125 6135 19159
rect 7205 19125 7239 19159
rect 7947 19125 7981 19159
rect 9505 19125 9539 19159
rect 9689 19125 9723 19159
rect 10149 19125 10183 19159
rect 10793 19125 10827 19159
rect 10885 19125 10919 19159
rect 11253 19125 11287 19159
rect 13461 19125 13495 19159
rect 13921 19125 13955 19159
rect 14749 19125 14783 19159
rect 14841 19125 14875 19159
rect 15209 19125 15243 19159
rect 15301 19125 15335 19159
rect 15669 19125 15703 19159
rect 16037 19125 16071 19159
rect 16129 19125 16163 19159
rect 16773 19125 16807 19159
rect 16957 19125 16991 19159
rect 19349 19125 19383 19159
rect 19441 19125 19475 19159
rect 21281 19125 21315 19159
rect 22201 19125 22235 19159
rect 23029 19125 23063 19159
rect 1777 18921 1811 18955
rect 4169 18921 4203 18955
rect 4629 18921 4663 18955
rect 4997 18921 5031 18955
rect 5273 18921 5307 18955
rect 8585 18921 8619 18955
rect 8953 18921 8987 18955
rect 11069 18921 11103 18955
rect 11529 18921 11563 18955
rect 13277 18921 13311 18955
rect 14197 18921 14231 18955
rect 14565 18921 14599 18955
rect 14841 18921 14875 18955
rect 22477 18921 22511 18955
rect 4261 18853 4295 18887
rect 5641 18853 5675 18887
rect 7858 18853 7892 18887
rect 8493 18853 8527 18887
rect 11437 18853 11471 18887
rect 16497 18853 16531 18887
rect 18797 18853 18831 18887
rect 18981 18853 19015 18887
rect 21364 18853 21398 18887
rect 2890 18785 2924 18819
rect 3157 18785 3191 18819
rect 4813 18785 4847 18819
rect 6101 18785 6135 18819
rect 9873 18785 9907 18819
rect 12164 18785 12198 18819
rect 13829 18785 13863 18819
rect 14381 18785 14415 18819
rect 14657 18785 14691 18819
rect 15189 18785 15223 18819
rect 17004 18785 17038 18819
rect 17417 18785 17451 18819
rect 19892 18785 19926 18819
rect 4077 18717 4111 18751
rect 5733 18717 5767 18751
rect 5917 18717 5951 18751
rect 8125 18717 8159 18751
rect 8309 18717 8343 18751
rect 9137 18717 9171 18751
rect 9460 18717 9494 18751
rect 9643 18717 9677 18751
rect 11621 18717 11655 18751
rect 11897 18717 11931 18751
rect 13645 18717 13679 18751
rect 13737 18717 13771 18751
rect 14933 18717 14967 18751
rect 16681 18717 16715 18751
rect 17144 18717 17178 18751
rect 18705 18717 18739 18751
rect 19625 18717 19659 18751
rect 21097 18717 21131 18751
rect 10977 18649 11011 18683
rect 16313 18649 16347 18683
rect 19257 18649 19291 18683
rect 6285 18581 6319 18615
rect 6745 18581 6779 18615
rect 18521 18581 18555 18615
rect 21005 18581 21039 18615
rect 2237 18377 2271 18411
rect 4721 18377 4755 18411
rect 7205 18377 7239 18411
rect 9689 18377 9723 18411
rect 13921 18377 13955 18411
rect 14749 18377 14783 18411
rect 18245 18377 18279 18411
rect 20361 18377 20395 18411
rect 3709 18309 3743 18343
rect 11713 18309 11747 18343
rect 16405 18309 16439 18343
rect 18429 18309 18463 18343
rect 1593 18241 1627 18275
rect 4353 18241 4387 18275
rect 4813 18241 4847 18275
rect 8309 18241 8343 18275
rect 8582 18241 8616 18275
rect 9597 18241 9631 18275
rect 11066 18241 11100 18275
rect 13093 18241 13127 18275
rect 14473 18241 14507 18275
rect 16129 18241 16163 18275
rect 17601 18241 17635 18275
rect 18705 18241 18739 18275
rect 22845 18241 22879 18275
rect 1685 18173 1719 18207
rect 3350 18173 3384 18207
rect 3610 18173 3644 18207
rect 4169 18173 4203 18207
rect 4537 18173 4571 18207
rect 5080 18173 5114 18207
rect 9045 18173 9079 18207
rect 10793 18173 10827 18207
rect 11529 18173 11563 18207
rect 15862 18173 15896 18207
rect 16221 18173 16255 18207
rect 17877 18173 17911 18207
rect 18613 18173 18647 18207
rect 18972 18173 19006 18207
rect 20177 18173 20211 18207
rect 20637 18173 20671 18207
rect 20904 18173 20938 18207
rect 22569 18173 22603 18207
rect 1777 18105 1811 18139
rect 12848 18105 12882 18139
rect 2145 18037 2179 18071
rect 4077 18037 4111 18071
rect 6193 18037 6227 18071
rect 6929 18037 6963 18071
rect 8578 18037 8612 18071
rect 9229 18037 9263 18071
rect 11062 18037 11096 18071
rect 13185 18037 13219 18071
rect 14289 18037 14323 18071
rect 14381 18037 14415 18071
rect 17233 18037 17267 18071
rect 17417 18037 17451 18071
rect 17785 18037 17819 18071
rect 20085 18037 20119 18071
rect 22017 18037 22051 18071
rect 22201 18037 22235 18071
rect 22661 18037 22695 18071
rect 3893 17833 3927 17867
rect 4813 17833 4847 17867
rect 9597 17833 9631 17867
rect 12265 17833 12299 17867
rect 13553 17833 13587 17867
rect 15761 17833 15795 17867
rect 17509 17833 17543 17867
rect 19625 17833 19659 17867
rect 22937 17833 22971 17867
rect 2412 17765 2446 17799
rect 5948 17765 5982 17799
rect 8042 17765 8076 17799
rect 11170 17765 11204 17799
rect 14626 17765 14660 17799
rect 16966 17765 17000 17799
rect 21640 17765 21674 17799
rect 4261 17697 4295 17731
rect 6193 17697 6227 17731
rect 6653 17697 6687 17731
rect 9505 17697 9539 17731
rect 12357 17697 12391 17731
rect 13185 17697 13219 17731
rect 14381 17697 14415 17731
rect 17325 17697 17359 17731
rect 17601 17697 17635 17731
rect 18328 17697 18362 17731
rect 20738 17697 20772 17731
rect 21097 17697 21131 17731
rect 23029 17697 23063 17731
rect 2145 17629 2179 17663
rect 4353 17629 4387 17663
rect 4537 17629 4571 17663
rect 8309 17629 8343 17663
rect 9689 17629 9723 17663
rect 11437 17629 11471 17663
rect 12173 17629 12207 17663
rect 12909 17629 12943 17663
rect 13093 17629 13127 17663
rect 17233 17629 17267 17663
rect 18061 17629 18095 17663
rect 21005 17629 21039 17663
rect 21373 17629 21407 17663
rect 3525 17561 3559 17595
rect 6929 17561 6963 17595
rect 9137 17561 9171 17595
rect 10057 17561 10091 17595
rect 15853 17561 15887 17595
rect 17785 17561 17819 17595
rect 19441 17561 19475 17595
rect 22753 17561 22787 17595
rect 6469 17493 6503 17527
rect 8953 17493 8987 17527
rect 12725 17493 12759 17527
rect 13737 17493 13771 17527
rect 17877 17493 17911 17527
rect 21281 17493 21315 17527
rect 1777 17289 1811 17323
rect 3249 17289 3283 17323
rect 6469 17289 6503 17323
rect 8217 17289 8251 17323
rect 13369 17289 13403 17323
rect 14933 17289 14967 17323
rect 16589 17289 16623 17323
rect 19073 17289 19107 17323
rect 19993 17289 20027 17323
rect 21005 17289 21039 17323
rect 10057 17221 10091 17255
rect 14841 17221 14875 17255
rect 17417 17221 17451 17255
rect 22017 17221 22051 17255
rect 4813 17153 4847 17187
rect 7021 17153 7055 17187
rect 7665 17153 7699 17187
rect 10701 17153 10735 17187
rect 16313 17153 16347 17187
rect 19257 17153 19291 17187
rect 20453 17153 20487 17187
rect 20545 17153 20579 17187
rect 21557 17153 21591 17187
rect 22661 17153 22695 17187
rect 22753 17153 22787 17187
rect 2901 17085 2935 17119
rect 3157 17085 3191 17119
rect 4362 17085 4396 17119
rect 4629 17085 4663 17119
rect 5080 17085 5114 17119
rect 8309 17085 8343 17119
rect 8565 17085 8599 17119
rect 9781 17085 9815 17119
rect 10425 17085 10459 17119
rect 11253 17085 11287 17119
rect 11989 17085 12023 17119
rect 12256 17085 12290 17119
rect 13461 17085 13495 17119
rect 13717 17085 13751 17119
rect 16046 17085 16080 17119
rect 16773 17085 16807 17119
rect 17325 17085 17359 17119
rect 17601 17085 17635 17119
rect 17700 17085 17734 17119
rect 19533 17085 19567 17119
rect 20361 17085 20395 17119
rect 21373 17085 21407 17119
rect 21833 17085 21867 17119
rect 22569 17085 22603 17119
rect 6929 17017 6963 17051
rect 7757 17017 7791 17051
rect 17049 17017 17083 17051
rect 17960 17017 17994 17051
rect 19441 17017 19475 17051
rect 21465 17017 21499 17051
rect 6193 16949 6227 16983
rect 6837 16949 6871 16983
rect 7849 16949 7883 16983
rect 9689 16949 9723 16983
rect 9965 16949 9999 16983
rect 10517 16949 10551 16983
rect 11437 16949 11471 16983
rect 17141 16949 17175 16983
rect 19901 16949 19935 16983
rect 22201 16949 22235 16983
rect 2973 16745 3007 16779
rect 4813 16745 4847 16779
rect 7021 16745 7055 16779
rect 7481 16745 7515 16779
rect 9137 16745 9171 16779
rect 9689 16745 9723 16779
rect 12541 16745 12575 16779
rect 15035 16745 15069 16779
rect 15945 16745 15979 16779
rect 17601 16745 17635 16779
rect 20821 16745 20855 16779
rect 5948 16677 5982 16711
rect 6469 16677 6503 16711
rect 8616 16677 8650 16711
rect 11406 16677 11440 16711
rect 13645 16677 13679 16711
rect 14565 16677 14599 16711
rect 17150 16677 17184 16711
rect 21732 16677 21766 16711
rect 1593 16609 1627 16643
rect 1860 16609 1894 16643
rect 4445 16609 4479 16643
rect 4721 16609 4755 16643
rect 6929 16609 6963 16643
rect 9597 16609 9631 16643
rect 10813 16609 10847 16643
rect 13001 16609 13035 16643
rect 13185 16609 13219 16643
rect 15485 16609 15519 16643
rect 15577 16609 15611 16643
rect 17417 16609 17451 16643
rect 18725 16609 18759 16643
rect 19073 16609 19107 16643
rect 19257 16609 19291 16643
rect 19993 16609 20027 16643
rect 20085 16609 20119 16643
rect 21465 16609 21499 16643
rect 23121 16609 23155 16643
rect 6193 16541 6227 16575
rect 6837 16541 6871 16575
rect 8861 16541 8895 16575
rect 11069 16541 11103 16575
rect 11161 16541 11195 16575
rect 12909 16541 12943 16575
rect 14473 16541 14507 16575
rect 14657 16541 14691 16575
rect 15393 16541 15427 16575
rect 18981 16541 19015 16575
rect 20269 16541 20303 16575
rect 20913 16541 20947 16575
rect 21005 16541 21039 16575
rect 7389 16473 7423 16507
rect 19625 16473 19659 16507
rect 20453 16473 20487 16507
rect 4261 16405 4295 16439
rect 4537 16405 4571 16439
rect 6377 16405 6411 16439
rect 9413 16405 9447 16439
rect 16037 16405 16071 16439
rect 19441 16405 19475 16439
rect 22845 16405 22879 16439
rect 22937 16405 22971 16439
rect 3433 16201 3467 16235
rect 6285 16201 6319 16235
rect 8401 16201 8435 16235
rect 14381 16201 14415 16235
rect 16773 16201 16807 16235
rect 18981 16201 19015 16235
rect 20177 16201 20211 16235
rect 21005 16201 21039 16235
rect 21833 16201 21867 16235
rect 22937 16201 22971 16235
rect 4721 16133 4755 16167
rect 4077 16065 4111 16099
rect 5365 16065 5399 16099
rect 5733 16065 5767 16099
rect 6469 16065 6503 16099
rect 8953 16065 8987 16099
rect 9413 16065 9447 16099
rect 9876 16065 9910 16099
rect 10149 16065 10183 16099
rect 11897 16065 11931 16099
rect 13737 16065 13771 16099
rect 14657 16065 14691 16099
rect 14933 16065 14967 16099
rect 15439 16065 15473 16099
rect 19533 16065 19567 16099
rect 20453 16065 20487 16099
rect 20545 16065 20579 16099
rect 21281 16065 21315 16099
rect 22385 16065 22419 16099
rect 22477 16065 22511 16099
rect 2053 15997 2087 16031
rect 4261 15997 4295 16031
rect 6929 15997 6963 16031
rect 12173 15997 12207 16031
rect 15669 15997 15703 16031
rect 16957 15997 16991 16031
rect 17509 15997 17543 16031
rect 17601 15997 17635 16031
rect 17868 15997 17902 16031
rect 19165 15997 19199 16031
rect 19717 15997 19751 16031
rect 21465 15997 21499 16031
rect 22569 15997 22603 16031
rect 1593 15929 1627 15963
rect 2298 15929 2332 15963
rect 5089 15929 5123 15963
rect 6653 15929 6687 15963
rect 6837 15929 6871 15963
rect 7196 15929 7230 15963
rect 12440 15929 12474 15963
rect 13921 15929 13955 15963
rect 21373 15929 21407 15963
rect 1501 15861 1535 15895
rect 4169 15861 4203 15895
rect 4629 15861 4663 15895
rect 5181 15861 5215 15895
rect 5825 15861 5859 15895
rect 5917 15861 5951 15895
rect 8309 15861 8343 15895
rect 8769 15861 8803 15895
rect 8861 15861 8895 15895
rect 9321 15861 9355 15895
rect 9879 15861 9913 15895
rect 11253 15861 11287 15895
rect 11345 15861 11379 15895
rect 12081 15861 12115 15895
rect 13553 15861 13587 15895
rect 14013 15861 14047 15895
rect 14841 15861 14875 15895
rect 15399 15861 15433 15895
rect 17141 15861 17175 15895
rect 17325 15861 17359 15895
rect 19349 15861 19383 15895
rect 19809 15861 19843 15895
rect 20637 15861 20671 15895
rect 6745 15657 6779 15691
rect 8217 15657 8251 15691
rect 8493 15657 8527 15691
rect 9413 15657 9447 15691
rect 9873 15657 9907 15691
rect 10333 15657 10367 15691
rect 12173 15657 12207 15691
rect 12731 15657 12765 15691
rect 14105 15657 14139 15691
rect 15853 15657 15887 15691
rect 17509 15657 17543 15691
rect 18981 15657 19015 15691
rect 19625 15657 19659 15691
rect 22753 15657 22787 15691
rect 7082 15589 7116 15623
rect 9505 15589 9539 15623
rect 15494 15589 15528 15623
rect 16966 15589 17000 15623
rect 18644 15589 18678 15623
rect 20738 15589 20772 15623
rect 21548 15589 21582 15623
rect 1501 15521 1535 15555
rect 1768 15521 1802 15555
rect 3341 15521 3375 15555
rect 3893 15521 3927 15555
rect 4160 15521 4194 15555
rect 5365 15521 5399 15555
rect 5632 15521 5666 15555
rect 8309 15521 8343 15555
rect 8585 15521 8619 15555
rect 11060 15521 11094 15555
rect 13001 15521 13035 15555
rect 15761 15521 15795 15555
rect 17417 15521 17451 15555
rect 19165 15521 19199 15555
rect 19441 15521 19475 15555
rect 21005 15521 21039 15555
rect 22937 15521 22971 15555
rect 3065 15453 3099 15487
rect 3249 15453 3283 15487
rect 6837 15453 6871 15487
rect 9321 15453 9355 15487
rect 10149 15453 10183 15487
rect 10241 15453 10275 15487
rect 10793 15453 10827 15487
rect 12265 15453 12299 15487
rect 12728 15453 12762 15487
rect 17233 15453 17267 15487
rect 18889 15453 18923 15487
rect 21281 15453 21315 15487
rect 8769 15385 8803 15419
rect 14381 15385 14415 15419
rect 2881 15317 2915 15351
rect 3709 15317 3743 15351
rect 5273 15317 5307 15351
rect 10701 15317 10735 15351
rect 19257 15317 19291 15351
rect 21097 15317 21131 15351
rect 22661 15317 22695 15351
rect 4905 15113 4939 15147
rect 4997 15113 5031 15147
rect 6469 15113 6503 15147
rect 8309 15113 8343 15147
rect 9229 15113 9263 15147
rect 10057 15113 10091 15147
rect 11713 15113 11747 15147
rect 14473 15113 14507 15147
rect 15761 15113 15795 15147
rect 17049 15113 17083 15147
rect 18153 15113 18187 15147
rect 21281 15113 21315 15147
rect 11529 15045 11563 15079
rect 3525 14977 3559 15011
rect 5457 14977 5491 15011
rect 5641 14977 5675 15011
rect 7021 14977 7055 15011
rect 7389 14977 7423 15011
rect 7573 14977 7607 15011
rect 8677 14977 8711 15011
rect 9505 14977 9539 15011
rect 9597 14977 9631 15011
rect 10149 14977 10183 15011
rect 12265 14977 12299 15011
rect 13093 14977 13127 15011
rect 15209 14977 15243 15011
rect 16221 14977 16255 15011
rect 16313 14977 16347 15011
rect 2053 14909 2087 14943
rect 5365 14909 5399 14943
rect 6837 14909 6871 14943
rect 7665 14909 7699 14943
rect 8125 14909 8159 14943
rect 8861 14909 8895 14943
rect 9689 14909 9723 14943
rect 12541 14909 12575 14943
rect 13360 14909 13394 14943
rect 15485 14909 15519 14943
rect 18429 14977 18463 15011
rect 22293 14977 22327 15011
rect 22477 14977 22511 15011
rect 17233 14909 17267 14943
rect 18061 14909 18095 14943
rect 18337 14909 18371 14943
rect 19901 14909 19935 14943
rect 21557 14909 21591 14943
rect 22569 14909 22603 14943
rect 2298 14841 2332 14875
rect 3792 14841 3826 14875
rect 6929 14841 6963 14875
rect 8769 14841 8803 14875
rect 10394 14841 10428 14875
rect 12725 14841 12759 14875
rect 15025 14841 15059 14875
rect 16129 14841 16163 14875
rect 16589 14841 16623 14875
rect 17049 14841 17083 14875
rect 17601 14841 17635 14875
rect 18696 14841 18730 14875
rect 20146 14841 20180 14875
rect 3433 14773 3467 14807
rect 8033 14773 8067 14807
rect 12081 14773 12115 14807
rect 12173 14773 12207 14807
rect 12909 14773 12943 14807
rect 14565 14773 14599 14807
rect 14933 14773 14967 14807
rect 15669 14773 15703 14807
rect 19809 14773 19843 14807
rect 21373 14773 21407 14807
rect 22017 14773 22051 14807
rect 22937 14773 22971 14807
rect 23581 14773 23615 14807
rect 4077 14569 4111 14603
rect 6009 14569 6043 14603
rect 6929 14569 6963 14603
rect 12541 14569 12575 14603
rect 13829 14569 13863 14603
rect 14197 14569 14231 14603
rect 14381 14569 14415 14603
rect 19993 14569 20027 14603
rect 20361 14569 20395 14603
rect 20821 14569 20855 14603
rect 22753 14569 22787 14603
rect 2890 14501 2924 14535
rect 4896 14501 4930 14535
rect 7450 14501 7484 14535
rect 11161 14501 11195 14535
rect 11253 14501 11287 14535
rect 12081 14501 12115 14535
rect 18337 14501 18371 14535
rect 18521 14501 18555 14535
rect 3157 14433 3191 14467
rect 3893 14433 3927 14467
rect 6193 14433 6227 14467
rect 7113 14433 7147 14467
rect 8769 14433 8803 14467
rect 9137 14433 9171 14467
rect 10537 14433 10571 14467
rect 12909 14433 12943 14467
rect 14565 14433 14599 14467
rect 14749 14433 14783 14467
rect 15292 14433 15326 14467
rect 16764 14433 16798 14467
rect 18613 14433 18647 14467
rect 18797 14433 18831 14467
rect 19165 14433 19199 14467
rect 19257 14433 19291 14467
rect 22405 14433 22439 14467
rect 22661 14433 22695 14467
rect 22937 14433 22971 14467
rect 4629 14365 4663 14399
rect 6745 14365 6779 14399
rect 7205 14365 7239 14399
rect 10793 14365 10827 14399
rect 11069 14365 11103 14399
rect 11805 14365 11839 14399
rect 11989 14365 12023 14399
rect 13001 14365 13035 14399
rect 13185 14365 13219 14399
rect 13645 14365 13679 14399
rect 13737 14365 13771 14399
rect 15025 14365 15059 14399
rect 16497 14365 16531 14399
rect 19809 14365 19843 14399
rect 19901 14365 19935 14399
rect 20637 14365 20671 14399
rect 20729 14365 20763 14399
rect 8953 14297 8987 14331
rect 9413 14297 9447 14331
rect 12449 14297 12483 14331
rect 18981 14297 19015 14331
rect 21189 14297 21223 14331
rect 1777 14229 1811 14263
rect 8585 14229 8619 14263
rect 9321 14229 9355 14263
rect 11621 14229 11655 14263
rect 14933 14229 14967 14263
rect 16405 14229 16439 14263
rect 17877 14229 17911 14263
rect 18061 14229 18095 14263
rect 19441 14229 19475 14263
rect 21281 14229 21315 14263
rect 1409 14025 1443 14059
rect 3617 14025 3651 14059
rect 3709 14025 3743 14059
rect 4721 14025 4755 14059
rect 6009 14025 6043 14059
rect 9689 14025 9723 14059
rect 11713 14025 11747 14059
rect 13277 14025 13311 14059
rect 13553 14025 13587 14059
rect 15761 14025 15795 14059
rect 19257 14025 19291 14059
rect 19717 14025 19751 14059
rect 22201 14025 22235 14059
rect 5733 13957 5767 13991
rect 9597 13957 9631 13991
rect 14289 13957 14323 13991
rect 16129 13957 16163 13991
rect 2973 13889 3007 13923
rect 3157 13889 3191 13923
rect 4169 13889 4203 13923
rect 4353 13889 4387 13923
rect 5181 13889 5215 13923
rect 9045 13889 9079 13923
rect 10149 13889 10183 13923
rect 10333 13889 10367 13923
rect 11161 13889 11195 13923
rect 13093 13889 13127 13923
rect 16589 13889 16623 13923
rect 16681 13889 16715 13923
rect 17417 13889 17451 13923
rect 17509 13889 17543 13923
rect 20453 13889 20487 13923
rect 22753 13889 22787 13923
rect 2533 13821 2567 13855
rect 2789 13821 2823 13855
rect 4077 13821 4111 13855
rect 4537 13821 4571 13855
rect 5273 13821 5307 13855
rect 5825 13821 5859 13855
rect 8502 13821 8536 13855
rect 8769 13821 8803 13855
rect 9137 13821 9171 13855
rect 10977 13821 11011 13855
rect 12826 13821 12860 13855
rect 13737 13821 13771 13855
rect 15577 13821 15611 13855
rect 15853 13821 15887 13855
rect 17785 13821 17819 13855
rect 17877 13821 17911 13855
rect 19441 13821 19475 13855
rect 19533 13821 19567 13855
rect 20637 13821 20671 13855
rect 20904 13821 20938 13855
rect 22661 13821 22695 13855
rect 23581 13821 23615 13855
rect 3249 13753 3283 13787
rect 9229 13753 9263 13787
rect 11345 13753 11379 13787
rect 13369 13753 13403 13787
rect 16589 13753 16623 13787
rect 18144 13753 18178 13787
rect 20177 13753 20211 13787
rect 20269 13753 20303 13787
rect 22569 13753 22603 13787
rect 5365 13685 5399 13719
rect 7389 13685 7423 13719
rect 10057 13685 10091 13719
rect 10517 13685 10551 13719
rect 10885 13685 10919 13719
rect 16957 13685 16991 13719
rect 17325 13685 17359 13719
rect 17785 13685 17819 13719
rect 19809 13685 19843 13719
rect 22017 13685 22051 13719
rect 23029 13685 23063 13719
rect 3341 13481 3375 13515
rect 3893 13481 3927 13515
rect 6193 13481 6227 13515
rect 6561 13481 6595 13515
rect 8769 13481 8803 13515
rect 9413 13481 9447 13515
rect 9873 13481 9907 13515
rect 10149 13481 10183 13515
rect 12449 13481 12483 13515
rect 17417 13481 17451 13515
rect 7656 13413 7690 13447
rect 9505 13413 9539 13447
rect 13952 13413 13986 13447
rect 14648 13413 14682 13447
rect 17754 13413 17788 13447
rect 18981 13413 19015 13447
rect 4261 13345 4295 13379
rect 4988 13345 5022 13379
rect 7205 13345 7239 13379
rect 9965 13345 9999 13379
rect 10609 13345 10643 13379
rect 11325 13345 11359 13379
rect 12541 13345 12575 13379
rect 14197 13345 14231 13379
rect 14381 13345 14415 13379
rect 16037 13345 16071 13379
rect 16304 13345 16338 13379
rect 19165 13345 19199 13379
rect 19349 13345 19383 13379
rect 19809 13345 19843 13379
rect 19993 13345 20027 13379
rect 22385 13345 22419 13379
rect 3065 13277 3099 13311
rect 3249 13277 3283 13311
rect 4353 13277 4387 13311
rect 4445 13277 4479 13311
rect 4721 13277 4755 13311
rect 6653 13277 6687 13311
rect 6745 13277 6779 13311
rect 7389 13277 7423 13311
rect 9321 13277 9355 13311
rect 10701 13277 10735 13311
rect 10885 13277 10919 13311
rect 11069 13277 11103 13311
rect 17509 13277 17543 13311
rect 20320 13277 20354 13311
rect 20499 13277 20533 13311
rect 20729 13277 20763 13311
rect 22477 13277 22511 13311
rect 22569 13277 22603 13311
rect 22845 13277 22879 13311
rect 3709 13209 3743 13243
rect 12725 13209 12759 13243
rect 22017 13209 22051 13243
rect 6101 13141 6135 13175
rect 7021 13141 7055 13175
rect 10241 13141 10275 13175
rect 12817 13141 12851 13175
rect 15761 13141 15795 13175
rect 18889 13141 18923 13175
rect 19625 13141 19659 13175
rect 21833 13141 21867 13175
rect 3985 12937 4019 12971
rect 5549 12937 5583 12971
rect 6469 12937 6503 12971
rect 7941 12937 7975 12971
rect 10793 12937 10827 12971
rect 14749 12937 14783 12971
rect 16497 12937 16531 12971
rect 20269 12937 20303 12971
rect 5457 12869 5491 12903
rect 20361 12869 20395 12903
rect 22845 12869 22879 12903
rect 6009 12801 6043 12835
rect 6101 12801 6135 12835
rect 10057 12801 10091 12835
rect 11345 12801 11379 12835
rect 13277 12801 13311 12835
rect 16221 12801 16255 12835
rect 17141 12801 17175 12835
rect 17233 12801 17267 12835
rect 19809 12801 19843 12835
rect 22385 12801 22419 12835
rect 2605 12733 2639 12767
rect 4077 12733 4111 12767
rect 5917 12733 5951 12767
rect 7582 12733 7616 12767
rect 7849 12733 7883 12767
rect 9054 12733 9088 12767
rect 9321 12733 9355 12767
rect 11161 12733 11195 12767
rect 13369 12733 13403 12767
rect 15954 12733 15988 12767
rect 16313 12733 16347 12767
rect 16589 12733 16623 12767
rect 17325 12733 17359 12767
rect 17785 12733 17819 12767
rect 18052 12733 18086 12767
rect 20085 12733 20119 12767
rect 21485 12733 21519 12767
rect 21741 12733 21775 12767
rect 2872 12665 2906 12699
rect 4344 12665 4378 12699
rect 13032 12665 13066 12699
rect 13636 12665 13670 12699
rect 19717 12665 19751 12699
rect 22293 12665 22327 12699
rect 9413 12597 9447 12631
rect 9781 12597 9815 12631
rect 9873 12597 9907 12631
rect 11253 12597 11287 12631
rect 11897 12597 11931 12631
rect 14841 12597 14875 12631
rect 16773 12597 16807 12631
rect 17693 12597 17727 12631
rect 19165 12597 19199 12631
rect 19257 12597 19291 12631
rect 19625 12597 19659 12631
rect 21833 12597 21867 12631
rect 22385 12597 22419 12631
rect 3617 12393 3651 12427
rect 5273 12393 5307 12427
rect 6745 12393 6779 12427
rect 8309 12393 8343 12427
rect 9413 12393 9447 12427
rect 9873 12393 9907 12427
rect 10241 12393 10275 12427
rect 11989 12393 12023 12427
rect 13737 12393 13771 12427
rect 16681 12393 16715 12427
rect 17877 12393 17911 12427
rect 19165 12393 19199 12427
rect 19625 12393 19659 12427
rect 19993 12393 20027 12427
rect 4160 12325 4194 12359
rect 5632 12325 5666 12359
rect 7196 12325 7230 12359
rect 17325 12325 17359 12359
rect 18797 12325 18831 12359
rect 3249 12257 3283 12291
rect 5365 12257 5399 12291
rect 8585 12257 8619 12291
rect 8677 12257 8711 12291
rect 9505 12257 9539 12291
rect 10057 12257 10091 12291
rect 10333 12257 10367 12291
rect 10876 12257 10910 12291
rect 12265 12257 12299 12291
rect 14749 12257 14783 12291
rect 15209 12257 15243 12291
rect 15485 12257 15519 12291
rect 16313 12257 16347 12291
rect 17969 12257 18003 12291
rect 19257 12257 19291 12291
rect 21750 12257 21784 12291
rect 22017 12257 22051 12291
rect 22569 12257 22603 12291
rect 22753 12257 22787 12291
rect 22845 12257 22879 12291
rect 2973 12189 3007 12223
rect 3157 12189 3191 12223
rect 3893 12189 3927 12223
rect 6929 12189 6963 12223
rect 9321 12189 9355 12223
rect 10609 12189 10643 12223
rect 14841 12189 14875 12223
rect 15025 12189 15059 12223
rect 16037 12189 16071 12223
rect 16221 12189 16255 12223
rect 17233 12189 17267 12223
rect 17417 12189 17451 12223
rect 17693 12189 17727 12223
rect 18613 12189 18647 12223
rect 18705 12189 18739 12223
rect 20085 12189 20119 12223
rect 20177 12189 20211 12223
rect 22109 12189 22143 12223
rect 8861 12121 8895 12155
rect 15393 12121 15427 12155
rect 16865 12121 16899 12155
rect 8401 12053 8435 12087
rect 10517 12053 10551 12087
rect 14381 12053 14415 12087
rect 15669 12053 15703 12087
rect 15853 12053 15887 12087
rect 18337 12053 18371 12087
rect 19441 12053 19475 12087
rect 20453 12053 20487 12087
rect 20637 12053 20671 12087
rect 3433 11849 3467 11883
rect 10885 11849 10919 11883
rect 12081 11849 12115 11883
rect 15025 11849 15059 11883
rect 17693 11849 17727 11883
rect 18061 11849 18095 11883
rect 22017 11849 22051 11883
rect 22201 11849 22235 11883
rect 3801 11781 3835 11815
rect 11161 11781 11195 11815
rect 14933 11781 14967 11815
rect 16497 11781 16531 11815
rect 17969 11781 18003 11815
rect 10241 11713 10275 11747
rect 13461 11713 13495 11747
rect 2053 11645 2087 11679
rect 3985 11645 4019 11679
rect 7021 11645 7055 11679
rect 8585 11645 8619 11679
rect 10977 11645 11011 11679
rect 13194 11645 13228 11679
rect 13553 11645 13587 11679
rect 16138 11645 16172 11679
rect 16405 11645 16439 11679
rect 2320 11577 2354 11611
rect 7288 11577 7322 11611
rect 8852 11577 8886 11611
rect 13820 11577 13854 11611
rect 17049 11713 17083 11747
rect 17233 11713 17267 11747
rect 20640 11713 20674 11747
rect 20913 11713 20947 11747
rect 22753 11713 22787 11747
rect 16773 11645 16807 11679
rect 17325 11645 17359 11679
rect 17785 11645 17819 11679
rect 19185 11645 19219 11679
rect 19441 11645 19475 11679
rect 20177 11645 20211 11679
rect 22569 11645 22603 11679
rect 19533 11577 19567 11611
rect 8401 11509 8435 11543
rect 9965 11509 9999 11543
rect 10425 11509 10459 11543
rect 10517 11509 10551 11543
rect 16497 11509 16531 11543
rect 16589 11509 16623 11543
rect 19901 11509 19935 11543
rect 20643 11509 20677 11543
rect 22661 11509 22695 11543
rect 2789 11305 2823 11339
rect 6837 11305 6871 11339
rect 8585 11305 8619 11339
rect 9781 11305 9815 11339
rect 11253 11305 11287 11339
rect 14197 11305 14231 11339
rect 14749 11305 14783 11339
rect 16773 11305 16807 11339
rect 17141 11305 17175 11339
rect 17601 11305 17635 11339
rect 17969 11305 18003 11339
rect 7972 11237 8006 11271
rect 10894 11237 10928 11271
rect 15660 11237 15694 11271
rect 18306 11237 18340 11271
rect 20922 11237 20956 11271
rect 21526 11237 21560 11271
rect 1409 11169 1443 11203
rect 1676 11169 1710 11203
rect 8769 11169 8803 11203
rect 12366 11169 12400 11203
rect 13084 11169 13118 11203
rect 14841 11169 14875 11203
rect 17233 11169 17267 11203
rect 17785 11169 17819 11203
rect 21189 11169 21223 11203
rect 21281 11169 21315 11203
rect 8217 11101 8251 11135
rect 11161 11101 11195 11135
rect 12633 11101 12667 11135
rect 12817 11101 12851 11135
rect 15025 11101 15059 11135
rect 15393 11101 15427 11135
rect 16957 11101 16991 11135
rect 18061 11101 18095 11135
rect 19625 11101 19659 11135
rect 22753 11101 22787 11135
rect 14381 11033 14415 11067
rect 19809 11033 19843 11067
rect 19441 10965 19475 10999
rect 22661 10965 22695 10999
rect 9137 10761 9171 10795
rect 10609 10761 10643 10795
rect 11713 10761 11747 10795
rect 12817 10761 12851 10795
rect 15025 10761 15059 10795
rect 16497 10761 16531 10795
rect 22017 10761 22051 10795
rect 8585 10625 8619 10659
rect 12173 10625 12207 10659
rect 12265 10625 12299 10659
rect 8318 10557 8352 10591
rect 8953 10557 8987 10591
rect 9229 10557 9263 10591
rect 9496 10557 9530 10591
rect 11345 10557 11379 10591
rect 14197 10557 14231 10591
rect 14289 10557 14323 10591
rect 14565 10557 14599 10591
rect 14749 10557 14783 10591
rect 16405 10557 16439 10591
rect 10793 10489 10827 10523
rect 12081 10489 12115 10523
rect 13952 10489 13986 10523
rect 16160 10489 16194 10523
rect 16773 10693 16807 10727
rect 22845 10693 22879 10727
rect 18705 10625 18739 10659
rect 19763 10625 19797 10659
rect 21465 10625 21499 10659
rect 16589 10557 16623 10591
rect 18429 10557 18463 10591
rect 18981 10557 19015 10591
rect 19257 10557 19291 10591
rect 19993 10557 20027 10591
rect 18184 10489 18218 10523
rect 21649 10489 21683 10523
rect 22293 10489 22327 10523
rect 22569 10489 22603 10523
rect 7205 10421 7239 10455
rect 14289 10421 14323 10455
rect 14381 10421 14415 10455
rect 14933 10421 14967 10455
rect 16497 10421 16531 10455
rect 17049 10421 17083 10455
rect 18797 10421 18831 10455
rect 19165 10421 19199 10455
rect 19723 10421 19757 10455
rect 21097 10421 21131 10455
rect 21557 10421 21591 10455
rect 22385 10421 22419 10455
rect 7573 10217 7607 10251
rect 9597 10217 9631 10251
rect 9689 10217 9723 10251
rect 10057 10217 10091 10251
rect 11529 10217 11563 10251
rect 15761 10217 15795 10251
rect 19257 10217 19291 10251
rect 22477 10217 22511 10251
rect 8708 10149 8742 10183
rect 10416 10149 10450 10183
rect 13829 10149 13863 10183
rect 16874 10149 16908 10183
rect 19870 10149 19904 10183
rect 10149 10081 10183 10115
rect 12929 10081 12963 10115
rect 14473 10081 14507 10115
rect 15025 10081 15059 10115
rect 17417 10081 17451 10115
rect 21353 10081 21387 10115
rect 23121 10081 23155 10115
rect 8953 10013 8987 10047
rect 9413 10013 9447 10047
rect 13185 10013 13219 10047
rect 13645 10013 13679 10047
rect 13737 10013 13771 10047
rect 17141 10013 17175 10047
rect 17740 10013 17774 10047
rect 17923 10013 17957 10047
rect 18153 10013 18187 10047
rect 19625 10013 19659 10047
rect 21097 10013 21131 10047
rect 22845 10013 22879 10047
rect 11805 9877 11839 9911
rect 14197 9877 14231 9911
rect 15669 9877 15703 9911
rect 17325 9877 17359 9911
rect 21005 9877 21039 9911
rect 16037 9673 16071 9707
rect 22201 9673 22235 9707
rect 8677 9605 8711 9639
rect 11529 9605 11563 9639
rect 11713 9605 11747 9639
rect 11805 9605 11839 9639
rect 13645 9605 13679 9639
rect 16497 9605 16531 9639
rect 16773 9605 16807 9639
rect 18613 9605 18647 9639
rect 22017 9605 22051 9639
rect 8125 9537 8159 9571
rect 8217 9537 8251 9571
rect 10977 9537 11011 9571
rect 9873 9469 9907 9503
rect 11161 9469 11195 9503
rect 13185 9537 13219 9571
rect 14013 9537 14047 9571
rect 14105 9537 14139 9571
rect 16221 9537 16255 9571
rect 19257 9537 19291 9571
rect 19625 9537 19659 9571
rect 19809 9537 19843 9571
rect 22753 9537 22787 9571
rect 14657 9469 14691 9503
rect 16313 9469 16347 9503
rect 16589 9469 16623 9503
rect 17141 9469 17175 9503
rect 17233 9469 17267 9503
rect 19901 9469 19935 9503
rect 20637 9469 20671 9503
rect 8309 9401 8343 9435
rect 11713 9401 11747 9435
rect 12918 9401 12952 9435
rect 13461 9401 13495 9435
rect 13645 9401 13679 9435
rect 14902 9401 14936 9435
rect 17500 9401 17534 9435
rect 20545 9401 20579 9435
rect 20904 9401 20938 9435
rect 22569 9401 22603 9435
rect 10057 9333 10091 9367
rect 11069 9333 11103 9367
rect 13369 9333 13403 9367
rect 14197 9333 14231 9367
rect 14565 9333 14599 9367
rect 16957 9333 16991 9367
rect 18705 9333 18739 9367
rect 19073 9333 19107 9367
rect 19165 9333 19199 9367
rect 20269 9333 20303 9367
rect 22661 9333 22695 9367
rect 23121 9333 23155 9367
rect 1593 9129 1627 9163
rect 13093 9129 13127 9163
rect 13461 9129 13495 9163
rect 14381 9129 14415 9163
rect 19901 9129 19935 9163
rect 20361 9129 20395 9163
rect 22937 9129 22971 9163
rect 13553 9061 13587 9095
rect 15494 9061 15528 9095
rect 17724 9061 17758 9095
rect 1409 8993 1443 9027
rect 1685 8993 1719 9027
rect 9137 8993 9171 9027
rect 9393 8993 9427 9027
rect 10977 8993 11011 9027
rect 11713 8993 11747 9027
rect 11980 8993 12014 9027
rect 15761 8993 15795 9027
rect 16037 8993 16071 9027
rect 16497 8993 16531 9027
rect 19174 8993 19208 9027
rect 19993 8993 20027 9027
rect 20913 8993 20947 9027
rect 21097 8993 21131 9027
rect 21189 8993 21223 9027
rect 21824 8993 21858 9027
rect 10793 8925 10827 8959
rect 10885 8925 10919 8959
rect 13369 8925 13403 8959
rect 17969 8925 18003 8959
rect 19441 8925 19475 8959
rect 19717 8925 19751 8959
rect 20453 8925 20487 8959
rect 21557 8925 21591 8959
rect 10517 8789 10551 8823
rect 11345 8789 11379 8823
rect 13921 8789 13955 8823
rect 15853 8789 15887 8823
rect 16313 8789 16347 8823
rect 16589 8789 16623 8823
rect 18061 8789 18095 8823
rect 1777 8585 1811 8619
rect 8861 8585 8895 8619
rect 11069 8585 11103 8619
rect 11529 8585 11563 8619
rect 14105 8585 14139 8619
rect 22017 8585 22051 8619
rect 16681 8517 16715 8551
rect 16957 8517 16991 8551
rect 17233 8517 17267 8551
rect 10425 8449 10459 8483
rect 10609 8449 10643 8483
rect 13737 8449 13771 8483
rect 16129 8449 16163 8483
rect 17693 8449 17727 8483
rect 17877 8449 17911 8483
rect 18800 8449 18834 8483
rect 22753 8449 22787 8483
rect 1961 8381 1995 8415
rect 2145 8381 2179 8415
rect 10241 8381 10275 8415
rect 10701 8381 10735 8415
rect 11345 8381 11379 8415
rect 13093 8381 13127 8415
rect 13553 8381 13587 8415
rect 15229 8381 15263 8415
rect 15485 8381 15519 8415
rect 17141 8381 17175 8415
rect 18061 8381 18095 8415
rect 18337 8381 18371 8415
rect 19073 8381 19107 8415
rect 20637 8381 20671 8415
rect 9996 8313 10030 8347
rect 12848 8313 12882 8347
rect 15577 8313 15611 8347
rect 16221 8313 16255 8347
rect 16405 8313 16439 8347
rect 17601 8313 17635 8347
rect 20545 8313 20579 8347
rect 20904 8313 20938 8347
rect 22661 8313 22695 8347
rect 11713 8245 11747 8279
rect 13185 8245 13219 8279
rect 13645 8245 13679 8279
rect 15853 8245 15887 8279
rect 18803 8245 18837 8279
rect 20177 8245 20211 8279
rect 22201 8245 22235 8279
rect 22569 8245 22603 8279
rect 9137 8041 9171 8075
rect 10885 8041 10919 8075
rect 11345 8041 11379 8075
rect 11621 8041 11655 8075
rect 12449 8041 12483 8075
rect 13277 8041 13311 8075
rect 13737 8041 13771 8075
rect 16405 8041 16439 8075
rect 16963 8041 16997 8075
rect 18337 8041 18371 8075
rect 18613 8041 18647 8075
rect 19441 8041 19475 8075
rect 10272 7973 10306 8007
rect 13369 7973 13403 8007
rect 13921 7973 13955 8007
rect 14473 7973 14507 8007
rect 18981 7973 19015 8007
rect 7389 7905 7423 7939
rect 8217 7905 8251 7939
rect 10977 7905 11011 7939
rect 11437 7905 11471 7939
rect 11897 7905 11931 7939
rect 12541 7905 12575 7939
rect 8493 7837 8527 7871
rect 10517 7837 10551 7871
rect 10701 7837 10735 7871
rect 12357 7837 12391 7871
rect 13185 7837 13219 7871
rect 12909 7769 12943 7803
rect 14013 7905 14047 7939
rect 14888 7905 14922 7939
rect 15301 7905 15335 7939
rect 17233 7905 17267 7939
rect 19073 7905 19107 7939
rect 19809 7905 19843 7939
rect 21833 7905 21867 7939
rect 22477 7905 22511 7939
rect 22661 7905 22695 7939
rect 14565 7837 14599 7871
rect 15028 7837 15062 7871
rect 16497 7837 16531 7871
rect 17003 7837 17037 7871
rect 18889 7837 18923 7871
rect 19901 7837 19935 7871
rect 20224 7837 20258 7871
rect 20407 7837 20441 7871
rect 20637 7837 20671 7871
rect 22385 7837 22419 7871
rect 23121 7837 23155 7871
rect 21741 7769 21775 7803
rect 12081 7701 12115 7735
rect 13921 7701 13955 7735
rect 14197 7701 14231 7735
rect 22017 7701 22051 7735
rect 10517 7497 10551 7531
rect 11989 7497 12023 7531
rect 13645 7497 13679 7531
rect 18061 7497 18095 7531
rect 18337 7497 18371 7531
rect 21741 7497 21775 7531
rect 22845 7497 22879 7531
rect 11897 7429 11931 7463
rect 21833 7429 21867 7463
rect 10793 7361 10827 7395
rect 12633 7361 12667 7395
rect 13001 7361 13035 7395
rect 13093 7361 13127 7395
rect 14197 7361 14231 7395
rect 14381 7361 14415 7395
rect 15117 7361 15151 7395
rect 15761 7361 15795 7395
rect 17417 7361 17451 7395
rect 17601 7361 17635 7395
rect 22385 7361 22419 7395
rect 9137 7293 9171 7327
rect 9404 7293 9438 7327
rect 11713 7293 11747 7327
rect 13185 7293 13219 7327
rect 14473 7293 14507 7327
rect 16221 7293 16255 7327
rect 16405 7293 16439 7327
rect 16497 7293 16531 7327
rect 17785 7293 17819 7327
rect 18245 7293 18279 7327
rect 19461 7293 19495 7327
rect 19717 7293 19751 7327
rect 20361 7293 20395 7327
rect 22017 7293 22051 7327
rect 23029 7293 23063 7327
rect 10885 7225 10919 7259
rect 12449 7225 12483 7259
rect 13829 7225 13863 7259
rect 14013 7225 14047 7259
rect 19901 7225 19935 7259
rect 20085 7225 20119 7259
rect 20269 7225 20303 7259
rect 20628 7225 20662 7259
rect 22293 7225 22327 7259
rect 10977 7157 11011 7191
rect 11345 7157 11379 7191
rect 12357 7157 12391 7191
rect 13553 7157 13587 7191
rect 14841 7157 14875 7191
rect 15209 7157 15243 7191
rect 15301 7157 15335 7191
rect 15669 7157 15703 7191
rect 16957 7157 16991 7191
rect 17325 7157 17359 7191
rect 22385 7157 22419 7191
rect 10977 6953 11011 6987
rect 11437 6953 11471 6987
rect 12265 6953 12299 6987
rect 13093 6953 13127 6987
rect 17233 6953 17267 6987
rect 20453 6953 20487 6987
rect 10272 6885 10306 6919
rect 11805 6817 11839 6851
rect 12633 6817 12667 6851
rect 13461 6817 13495 6851
rect 14013 6817 14047 6851
rect 14648 6817 14682 6851
rect 16109 6817 16143 6851
rect 18438 6817 18472 6851
rect 18797 6817 18831 6851
rect 19349 6817 19383 6851
rect 19809 6817 19843 6851
rect 20913 6817 20947 6851
rect 22762 6817 22796 6851
rect 10517 6749 10551 6783
rect 10701 6749 10735 6783
rect 10885 6749 10919 6783
rect 11897 6749 11931 6783
rect 11989 6749 12023 6783
rect 12725 6749 12759 6783
rect 12909 6749 12943 6783
rect 13553 6749 13587 6783
rect 13645 6749 13679 6783
rect 14381 6749 14415 6783
rect 15853 6749 15887 6783
rect 18705 6749 18739 6783
rect 19073 6749 19107 6783
rect 20269 6749 20303 6783
rect 20361 6749 20395 6783
rect 23029 6749 23063 6783
rect 11345 6681 11379 6715
rect 17325 6681 17359 6715
rect 19993 6681 20027 6715
rect 21097 6681 21131 6715
rect 9137 6613 9171 6647
rect 14197 6613 14231 6647
rect 15761 6613 15795 6647
rect 20821 6613 20855 6647
rect 21189 6613 21223 6647
rect 21649 6613 21683 6647
rect 10057 6409 10091 6443
rect 11529 6409 11563 6443
rect 13093 6409 13127 6443
rect 14565 6409 14599 6443
rect 16037 6409 16071 6443
rect 16589 6409 16623 6443
rect 18337 6409 18371 6443
rect 18521 6409 18555 6443
rect 19349 6409 19383 6443
rect 10149 6273 10183 6307
rect 18797 6273 18831 6307
rect 21465 6273 21499 6307
rect 8677 6205 8711 6239
rect 8944 6205 8978 6239
rect 11713 6205 11747 6239
rect 13185 6205 13219 6239
rect 14657 6205 14691 6239
rect 14913 6205 14947 6239
rect 16129 6205 16163 6239
rect 16957 6205 16991 6239
rect 19441 6205 19475 6239
rect 21281 6205 21315 6239
rect 22293 6205 22327 6239
rect 10416 6137 10450 6171
rect 11980 6137 12014 6171
rect 13430 6137 13464 6171
rect 17202 6137 17236 6171
rect 18889 6137 18923 6171
rect 19708 6137 19742 6171
rect 21741 6137 21775 6171
rect 21925 6137 21959 6171
rect 22753 6137 22787 6171
rect 18981 6069 19015 6103
rect 20821 6069 20855 6103
rect 20913 6069 20947 6103
rect 21373 6069 21407 6103
rect 11069 5865 11103 5899
rect 12541 5865 12575 5899
rect 14013 5865 14047 5899
rect 14565 5865 14599 5899
rect 15301 5865 15335 5899
rect 17325 5865 17359 5899
rect 17693 5865 17727 5899
rect 18337 5865 18371 5899
rect 18613 5865 18647 5899
rect 19441 5865 19475 5899
rect 21557 5865 21591 5899
rect 9956 5797 9990 5831
rect 11428 5797 11462 5831
rect 12878 5797 12912 5831
rect 16190 5797 16224 5831
rect 21097 5797 21131 5831
rect 21281 5797 21315 5831
rect 22670 5797 22704 5831
rect 9689 5729 9723 5763
rect 11161 5729 11195 5763
rect 14381 5729 14415 5763
rect 14657 5729 14691 5763
rect 15393 5729 15427 5763
rect 15945 5729 15979 5763
rect 17785 5729 17819 5763
rect 18429 5729 18463 5763
rect 19073 5729 19107 5763
rect 19892 5729 19926 5763
rect 22937 5729 22971 5763
rect 12633 5661 12667 5695
rect 15209 5661 15243 5695
rect 17601 5661 17635 5695
rect 18889 5661 18923 5695
rect 18981 5661 19015 5695
rect 19625 5661 19659 5695
rect 14841 5593 14875 5627
rect 21005 5593 21039 5627
rect 15761 5525 15795 5559
rect 18153 5525 18187 5559
rect 21465 5525 21499 5559
rect 12265 5321 12299 5355
rect 18337 5321 18371 5355
rect 16037 5253 16071 5287
rect 13645 5185 13679 5219
rect 16129 5185 16163 5219
rect 16957 5185 16991 5219
rect 18889 5185 18923 5219
rect 18981 5185 19015 5219
rect 19441 5185 19475 5219
rect 19625 5185 19659 5219
rect 21005 5185 21039 5219
rect 21281 5185 21315 5219
rect 22661 5185 22695 5219
rect 22753 5185 22787 5219
rect 13389 5117 13423 5151
rect 15853 5117 15887 5151
rect 16589 5117 16623 5151
rect 17224 5117 17258 5151
rect 19809 5117 19843 5151
rect 21465 5117 21499 5151
rect 19901 5049 19935 5083
rect 21557 5049 21591 5083
rect 23029 5049 23063 5083
rect 16773 4981 16807 5015
rect 18429 4981 18463 5015
rect 18797 4981 18831 5015
rect 20269 4981 20303 5015
rect 20361 4981 20395 5015
rect 20729 4981 20763 5015
rect 20821 4981 20855 5015
rect 21925 4981 21959 5015
rect 22201 4981 22235 5015
rect 22569 4981 22603 5015
rect 16313 4777 16347 4811
rect 18613 4777 18647 4811
rect 17540 4709 17574 4743
rect 19892 4709 19926 4743
rect 21373 4709 21407 4743
rect 16129 4641 16163 4675
rect 18153 4641 18187 4675
rect 18245 4641 18279 4675
rect 19073 4641 19107 4675
rect 21189 4641 21223 4675
rect 22578 4641 22612 4675
rect 22845 4641 22879 4675
rect 23121 4641 23155 4675
rect 17785 4573 17819 4607
rect 18061 4573 18095 4607
rect 19165 4573 19199 4607
rect 19257 4573 19291 4607
rect 19625 4573 19659 4607
rect 16405 4505 16439 4539
rect 21465 4505 21499 4539
rect 18705 4437 18739 4471
rect 21005 4437 21039 4471
rect 22937 4437 22971 4471
rect 16037 4233 16071 4267
rect 22201 4233 22235 4267
rect 18337 4165 18371 4199
rect 22017 4165 22051 4199
rect 16589 4097 16623 4131
rect 16957 4097 16991 4131
rect 20177 4097 20211 4131
rect 20545 4097 20579 4131
rect 22753 4097 22787 4131
rect 16405 4029 16439 4063
rect 17224 4029 17258 4063
rect 18429 4029 18463 4063
rect 20361 4029 20395 4063
rect 20637 4029 20671 4063
rect 22569 4029 22603 4063
rect 15945 3961 15979 3995
rect 18696 3961 18730 3995
rect 19993 3961 20027 3995
rect 20904 3961 20938 3995
rect 22661 3961 22695 3995
rect 16497 3893 16531 3927
rect 19809 3893 19843 3927
rect 23121 3893 23155 3927
rect 23581 3893 23615 3927
rect 16405 3689 16439 3723
rect 19349 3689 19383 3723
rect 21373 3689 21407 3723
rect 22845 3689 22879 3723
rect 22937 3689 22971 3723
rect 3341 3621 3375 3655
rect 17632 3621 17666 3655
rect 19717 3621 19751 3655
rect 19901 3621 19935 3655
rect 20260 3621 20294 3655
rect 2697 3553 2731 3587
rect 17877 3553 17911 3587
rect 17969 3553 18003 3587
rect 18236 3553 18270 3587
rect 19993 3553 20027 3587
rect 21465 3553 21499 3587
rect 21732 3553 21766 3587
rect 23121 3553 23155 3587
rect 3709 3349 3743 3383
rect 16497 3349 16531 3383
rect 2421 3145 2455 3179
rect 18429 3145 18463 3179
rect 19349 3145 19383 3179
rect 19441 3145 19475 3179
rect 20913 3145 20947 3179
rect 1409 3077 1443 3111
rect 19073 3009 19107 3043
rect 21465 3009 21499 3043
rect 23581 3009 23615 3043
rect 1593 2941 1627 2975
rect 1961 2941 1995 2975
rect 2237 2941 2271 2975
rect 2697 2941 2731 2975
rect 6101 2941 6135 2975
rect 16957 2941 16991 2975
rect 17224 2941 17258 2975
rect 18889 2941 18923 2975
rect 20821 2941 20855 2975
rect 21281 2941 21315 2975
rect 21833 2941 21867 2975
rect 22661 2941 22695 2975
rect 22937 2941 22971 2975
rect 18797 2873 18831 2907
rect 20576 2873 20610 2907
rect 22385 2873 22419 2907
rect 2513 2805 2547 2839
rect 2881 2805 2915 2839
rect 18337 2805 18371 2839
rect 21373 2805 21407 2839
rect 21925 2805 21959 2839
rect 23029 2805 23063 2839
rect 10701 2601 10735 2635
rect 18613 2601 18647 2635
rect 19165 2601 19199 2635
rect 19717 2601 19751 2635
rect 22569 2601 22603 2635
rect 2237 2533 2271 2567
rect 6285 2533 6319 2567
rect 10425 2533 10459 2567
rect 17500 2533 17534 2567
rect 22937 2533 22971 2567
rect 14749 2465 14783 2499
rect 17233 2465 17267 2499
rect 18889 2465 18923 2499
rect 19533 2465 19567 2499
rect 19993 2465 20027 2499
rect 20361 2465 20395 2499
rect 20637 2465 20671 2499
rect 20904 2465 20938 2499
rect 22201 2465 22235 2499
rect 22753 2465 22787 2499
rect 20545 2397 20579 2431
rect 22385 2397 22419 2431
rect 2053 2329 2087 2363
rect 6101 2329 6135 2363
rect 10241 2329 10275 2363
rect 18981 2329 19015 2363
rect 23121 2329 23155 2363
rect 23581 2329 23615 2363
rect 14841 2261 14875 2295
rect 17049 2261 17083 2295
rect 19441 2261 19475 2295
rect 20177 2261 20211 2295
rect 22017 2261 22051 2295
rect 23581 1377 23615 1411
<< metal1 >>
rect 10134 22516 10140 22568
rect 10192 22556 10198 22568
rect 10594 22556 10600 22568
rect 10192 22528 10600 22556
rect 10192 22516 10198 22528
rect 10594 22516 10600 22528
rect 10652 22556 10658 22568
rect 11606 22556 11612 22568
rect 10652 22528 11612 22556
rect 10652 22516 10658 22528
rect 11606 22516 11612 22528
rect 11664 22516 11670 22568
rect 15102 22516 15108 22568
rect 15160 22556 15166 22568
rect 16206 22556 16212 22568
rect 15160 22528 16212 22556
rect 15160 22516 15166 22528
rect 16206 22516 16212 22528
rect 16264 22516 16270 22568
rect 9858 22448 9864 22500
rect 9916 22488 9922 22500
rect 17402 22488 17408 22500
rect 9916 22460 17408 22488
rect 9916 22448 9922 22460
rect 17402 22448 17408 22460
rect 17460 22488 17466 22500
rect 18414 22488 18420 22500
rect 17460 22460 18420 22488
rect 17460 22448 17466 22460
rect 18414 22448 18420 22460
rect 18472 22448 18478 22500
rect 5442 22380 5448 22432
rect 5500 22420 5506 22432
rect 5902 22420 5908 22432
rect 5500 22392 5908 22420
rect 5500 22380 5506 22392
rect 5902 22380 5908 22392
rect 5960 22420 5966 22432
rect 6638 22420 6644 22432
rect 5960 22392 6644 22420
rect 5960 22380 5966 22392
rect 6638 22380 6644 22392
rect 6696 22380 6702 22432
rect 9950 22380 9956 22432
rect 10008 22420 10014 22432
rect 12250 22420 12256 22432
rect 10008 22392 12256 22420
rect 10008 22380 10014 22392
rect 12250 22380 12256 22392
rect 12308 22380 12314 22432
rect 15010 22380 15016 22432
rect 15068 22420 15074 22432
rect 18874 22420 18880 22432
rect 15068 22392 18880 22420
rect 15068 22380 15074 22392
rect 18874 22380 18880 22392
rect 18932 22380 18938 22432
rect 1104 22330 23460 22352
rect 1104 22278 8446 22330
rect 8498 22278 8510 22330
rect 8562 22278 8574 22330
rect 8626 22278 8638 22330
rect 8690 22278 15910 22330
rect 15962 22278 15974 22330
rect 16026 22278 16038 22330
rect 16090 22278 16102 22330
rect 16154 22278 23460 22330
rect 1104 22256 23460 22278
rect 3697 22219 3755 22225
rect 3697 22185 3709 22219
rect 3743 22185 3755 22219
rect 3697 22179 3755 22185
rect 5169 22219 5227 22225
rect 5169 22185 5181 22219
rect 5215 22185 5227 22219
rect 5169 22179 5227 22185
rect 5644 22188 6224 22216
rect 3712 22148 3740 22179
rect 4065 22151 4123 22157
rect 4065 22148 4077 22151
rect 3712 22120 4077 22148
rect 4065 22117 4077 22120
rect 4111 22117 4123 22151
rect 4065 22111 4123 22117
rect 4433 22151 4491 22157
rect 4433 22117 4445 22151
rect 4479 22148 4491 22151
rect 5184 22148 5212 22179
rect 5644 22157 5672 22188
rect 4479 22120 5212 22148
rect 5629 22151 5687 22157
rect 4479 22117 4491 22120
rect 4433 22111 4491 22117
rect 5629 22117 5641 22151
rect 5675 22117 5687 22151
rect 5629 22111 5687 22117
rect 5902 22108 5908 22160
rect 5960 22148 5966 22160
rect 6196 22148 6224 22188
rect 7466 22176 7472 22228
rect 7524 22216 7530 22228
rect 7837 22219 7895 22225
rect 7837 22216 7849 22219
rect 7524 22188 7849 22216
rect 7524 22176 7530 22188
rect 7837 22185 7849 22188
rect 7883 22185 7895 22219
rect 7837 22179 7895 22185
rect 8205 22219 8263 22225
rect 8205 22185 8217 22219
rect 8251 22216 8263 22219
rect 8481 22219 8539 22225
rect 8481 22216 8493 22219
rect 8251 22188 8493 22216
rect 8251 22185 8263 22188
rect 8205 22179 8263 22185
rect 8481 22185 8493 22188
rect 8527 22185 8539 22219
rect 8481 22179 8539 22185
rect 11698 22176 11704 22228
rect 11756 22216 11762 22228
rect 12161 22219 12219 22225
rect 12161 22216 12173 22219
rect 11756 22188 12173 22216
rect 11756 22176 11762 22188
rect 12161 22185 12173 22188
rect 12207 22185 12219 22219
rect 12161 22179 12219 22185
rect 14458 22176 14464 22228
rect 14516 22216 14522 22228
rect 15010 22216 15016 22228
rect 14516 22188 15016 22216
rect 14516 22176 14522 22188
rect 15010 22176 15016 22188
rect 15068 22176 15074 22228
rect 15657 22219 15715 22225
rect 15657 22216 15669 22219
rect 15580 22188 15669 22216
rect 8294 22148 8300 22160
rect 5960 22120 6132 22148
rect 6196 22120 8300 22148
rect 5960 22108 5966 22120
rect 290 22040 296 22092
rect 348 22080 354 22092
rect 1397 22083 1455 22089
rect 1397 22080 1409 22083
rect 348 22052 1409 22080
rect 348 22040 354 22052
rect 1397 22049 1409 22052
rect 1443 22049 1455 22083
rect 1578 22080 1584 22092
rect 1539 22052 1584 22080
rect 1397 22043 1455 22049
rect 1578 22040 1584 22052
rect 1636 22040 1642 22092
rect 1946 22080 1952 22092
rect 1907 22052 1952 22080
rect 1946 22040 1952 22052
rect 2004 22040 2010 22092
rect 2314 22080 2320 22092
rect 2275 22052 2320 22080
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 2682 22080 2688 22092
rect 2643 22052 2688 22080
rect 2682 22040 2688 22052
rect 2740 22040 2746 22092
rect 2866 22080 2872 22092
rect 2827 22052 2872 22080
rect 2866 22040 2872 22052
rect 2924 22040 2930 22092
rect 3053 22083 3111 22089
rect 3053 22049 3065 22083
rect 3099 22080 3111 22083
rect 3326 22080 3332 22092
rect 3099 22052 3332 22080
rect 3099 22049 3111 22052
rect 3053 22043 3111 22049
rect 3326 22040 3332 22052
rect 3384 22040 3390 22092
rect 3513 22083 3571 22089
rect 3513 22049 3525 22083
rect 3559 22049 3571 22083
rect 3513 22043 3571 22049
rect 934 21972 940 22024
rect 992 22012 998 22024
rect 1765 22015 1823 22021
rect 1765 22012 1777 22015
rect 992 21984 1777 22012
rect 992 21972 998 21984
rect 1765 21981 1777 21984
rect 1811 21981 1823 22015
rect 1765 21975 1823 21981
rect 2222 21972 2228 22024
rect 2280 22012 2286 22024
rect 2501 22015 2559 22021
rect 2501 22012 2513 22015
rect 2280 21984 2513 22012
rect 2280 21972 2286 21984
rect 2501 21981 2513 21984
rect 2547 21981 2559 22015
rect 2501 21975 2559 21981
rect 2590 21972 2596 22024
rect 2648 22012 2654 22024
rect 3528 22012 3556 22043
rect 4154 22040 4160 22092
rect 4212 22080 4218 22092
rect 4249 22083 4307 22089
rect 4249 22080 4261 22083
rect 4212 22052 4261 22080
rect 4212 22040 4218 22052
rect 4249 22049 4261 22052
rect 4295 22049 4307 22083
rect 4798 22080 4804 22092
rect 4759 22052 4804 22080
rect 4249 22043 4307 22049
rect 4798 22040 4804 22052
rect 4856 22040 4862 22092
rect 4985 22083 5043 22089
rect 4985 22049 4997 22083
rect 5031 22049 5043 22083
rect 5350 22080 5356 22092
rect 5311 22052 5356 22080
rect 4985 22043 5043 22049
rect 4522 22012 4528 22024
rect 2648 21984 4528 22012
rect 2648 21972 2654 21984
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 5000 22012 5028 22043
rect 5350 22040 5356 22052
rect 5408 22040 5414 22092
rect 6104 22089 6132 22120
rect 8294 22108 8300 22120
rect 8352 22108 8358 22160
rect 9582 22108 9588 22160
rect 9640 22148 9646 22160
rect 10778 22148 10784 22160
rect 9640 22120 10088 22148
rect 10739 22120 10784 22148
rect 9640 22108 9646 22120
rect 5989 22083 6047 22089
rect 5989 22080 6001 22083
rect 5920 22052 6001 22080
rect 5000 21984 5856 22012
rect 1670 21904 1676 21956
rect 1728 21944 1734 21956
rect 2133 21947 2191 21953
rect 2133 21944 2145 21947
rect 1728 21916 2145 21944
rect 1728 21904 1734 21916
rect 2133 21913 2145 21916
rect 2179 21913 2191 21947
rect 2133 21907 2191 21913
rect 3510 21904 3516 21956
rect 3568 21944 3574 21956
rect 5828 21953 5856 21984
rect 3881 21947 3939 21953
rect 3881 21944 3893 21947
rect 3568 21916 3893 21944
rect 3568 21904 3574 21916
rect 3881 21913 3893 21916
rect 3927 21913 3939 21947
rect 3881 21907 3939 21913
rect 4709 21947 4767 21953
rect 4709 21913 4721 21947
rect 4755 21944 4767 21947
rect 5813 21947 5871 21953
rect 4755 21916 5764 21944
rect 4755 21913 4767 21916
rect 4709 21907 4767 21913
rect 2406 21836 2412 21888
rect 2464 21876 2470 21888
rect 3329 21879 3387 21885
rect 3329 21876 3341 21879
rect 2464 21848 3341 21876
rect 2464 21836 2470 21848
rect 3329 21845 3341 21848
rect 3375 21876 3387 21879
rect 5350 21876 5356 21888
rect 3375 21848 5356 21876
rect 3375 21845 3387 21848
rect 3329 21839 3387 21845
rect 5350 21836 5356 21848
rect 5408 21836 5414 21888
rect 5442 21836 5448 21888
rect 5500 21876 5506 21888
rect 5537 21879 5595 21885
rect 5537 21876 5549 21879
rect 5500 21848 5549 21876
rect 5500 21836 5506 21848
rect 5537 21845 5549 21848
rect 5583 21845 5595 21879
rect 5736 21876 5764 21916
rect 5813 21913 5825 21947
rect 5859 21913 5871 21947
rect 5920 21944 5948 22052
rect 5989 22049 6001 22052
rect 6035 22049 6047 22083
rect 5989 22043 6047 22049
rect 6081 22083 6139 22089
rect 6081 22049 6093 22083
rect 6127 22049 6139 22083
rect 6081 22043 6139 22049
rect 6270 22040 6276 22092
rect 6328 22080 6334 22092
rect 6733 22083 6791 22089
rect 6733 22080 6745 22083
rect 6328 22052 6745 22080
rect 6328 22040 6334 22052
rect 6733 22049 6745 22052
rect 6779 22049 6791 22083
rect 7006 22080 7012 22092
rect 6967 22052 7012 22080
rect 6733 22043 6791 22049
rect 7006 22040 7012 22052
rect 7064 22040 7070 22092
rect 7374 22080 7380 22092
rect 7287 22052 7380 22080
rect 7374 22040 7380 22052
rect 7432 22040 7438 22092
rect 7834 22040 7840 22092
rect 7892 22080 7898 22092
rect 8665 22083 8723 22089
rect 7892 22052 8524 22080
rect 7892 22040 7898 22052
rect 7392 21944 7420 22040
rect 7558 22012 7564 22024
rect 7519 21984 7564 22012
rect 7558 21972 7564 21984
rect 7616 21972 7622 22024
rect 7742 22012 7748 22024
rect 7703 21984 7748 22012
rect 7742 21972 7748 21984
rect 7800 21972 7806 22024
rect 7926 21972 7932 22024
rect 7984 22012 7990 22024
rect 8389 22015 8447 22021
rect 8389 22012 8401 22015
rect 7984 21984 8401 22012
rect 7984 21972 7990 21984
rect 8389 21981 8401 21984
rect 8435 21981 8447 22015
rect 8389 21975 8447 21981
rect 8110 21944 8116 21956
rect 5920 21916 7328 21944
rect 7392 21916 8116 21944
rect 5813 21907 5871 21913
rect 6086 21876 6092 21888
rect 5736 21848 6092 21876
rect 5537 21839 5595 21845
rect 6086 21836 6092 21848
rect 6144 21836 6150 21888
rect 6270 21876 6276 21888
rect 6231 21848 6276 21876
rect 6270 21836 6276 21848
rect 6328 21836 6334 21888
rect 6546 21876 6552 21888
rect 6507 21848 6552 21876
rect 6546 21836 6552 21848
rect 6604 21836 6610 21888
rect 6638 21836 6644 21888
rect 6696 21876 6702 21888
rect 6825 21879 6883 21885
rect 6825 21876 6837 21879
rect 6696 21848 6837 21876
rect 6696 21836 6702 21848
rect 6825 21845 6837 21848
rect 6871 21845 6883 21879
rect 6825 21839 6883 21845
rect 7098 21836 7104 21888
rect 7156 21876 7162 21888
rect 7193 21879 7251 21885
rect 7193 21876 7205 21879
rect 7156 21848 7205 21876
rect 7156 21836 7162 21848
rect 7193 21845 7205 21848
rect 7239 21845 7251 21879
rect 7300 21876 7328 21916
rect 8110 21904 8116 21916
rect 8168 21904 8174 21956
rect 8496 21944 8524 22052
rect 8665 22049 8677 22083
rect 8711 22080 8723 22083
rect 9217 22083 9275 22089
rect 9217 22080 9229 22083
rect 8711 22052 9229 22080
rect 8711 22049 8723 22052
rect 8665 22043 8723 22049
rect 9217 22049 9229 22052
rect 9263 22049 9275 22083
rect 9217 22043 9275 22049
rect 9674 22040 9680 22092
rect 9732 22080 9738 22092
rect 10060 22089 10088 22120
rect 10778 22108 10784 22120
rect 10836 22108 10842 22160
rect 13630 22108 13636 22160
rect 13688 22148 13694 22160
rect 13725 22151 13783 22157
rect 13725 22148 13737 22151
rect 13688 22120 13737 22148
rect 13688 22108 13694 22120
rect 13725 22117 13737 22120
rect 13771 22117 13783 22151
rect 13725 22111 13783 22117
rect 13814 22108 13820 22160
rect 13872 22148 13878 22160
rect 15580 22157 15608 22188
rect 15657 22185 15669 22188
rect 15703 22185 15715 22219
rect 18874 22216 18880 22228
rect 18835 22188 18880 22216
rect 15657 22179 15715 22185
rect 18874 22176 18880 22188
rect 18932 22176 18938 22228
rect 22278 22216 22284 22228
rect 22204 22188 22284 22216
rect 15565 22151 15623 22157
rect 13872 22120 14412 22148
rect 13872 22108 13878 22120
rect 14384 22092 14412 22120
rect 15565 22117 15577 22151
rect 15611 22117 15623 22151
rect 16206 22148 16212 22160
rect 15565 22111 15623 22117
rect 15856 22120 16212 22148
rect 9861 22083 9919 22089
rect 9861 22080 9873 22083
rect 9732 22052 9873 22080
rect 9732 22040 9738 22052
rect 9861 22049 9873 22052
rect 9907 22049 9919 22083
rect 9861 22043 9919 22049
rect 10045 22083 10103 22089
rect 10045 22049 10057 22083
rect 10091 22080 10103 22083
rect 11606 22080 11612 22092
rect 10091 22052 10125 22080
rect 11567 22052 11612 22080
rect 10091 22049 10103 22052
rect 10045 22043 10103 22049
rect 11606 22040 11612 22052
rect 11664 22040 11670 22092
rect 11882 22040 11888 22092
rect 11940 22080 11946 22092
rect 12069 22083 12127 22089
rect 12069 22080 12081 22083
rect 11940 22052 12081 22080
rect 11940 22040 11946 22052
rect 12069 22049 12081 22052
rect 12115 22049 12127 22083
rect 12069 22043 12127 22049
rect 12250 22040 12256 22092
rect 12308 22080 12314 22092
rect 12345 22083 12403 22089
rect 12345 22080 12357 22083
rect 12308 22052 12357 22080
rect 12308 22040 12314 22052
rect 12345 22049 12357 22052
rect 12391 22049 12403 22083
rect 12710 22080 12716 22092
rect 12671 22052 12716 22080
rect 12345 22043 12403 22049
rect 12710 22040 12716 22052
rect 12768 22040 12774 22092
rect 12802 22040 12808 22092
rect 12860 22080 12866 22092
rect 12860 22052 12905 22080
rect 12860 22040 12866 22052
rect 12986 22040 12992 22092
rect 13044 22080 13050 22092
rect 13081 22083 13139 22089
rect 13081 22080 13093 22083
rect 13044 22052 13093 22080
rect 13044 22040 13050 22052
rect 13081 22049 13093 22052
rect 13127 22080 13139 22083
rect 13170 22080 13176 22092
rect 13127 22052 13176 22080
rect 13127 22049 13139 22052
rect 13081 22043 13139 22049
rect 13170 22040 13176 22052
rect 13228 22040 13234 22092
rect 14366 22080 14372 22092
rect 14279 22052 14372 22080
rect 14366 22040 14372 22052
rect 14424 22040 14430 22092
rect 14553 22083 14611 22089
rect 14553 22049 14565 22083
rect 14599 22080 14611 22083
rect 15010 22080 15016 22092
rect 14599 22052 14872 22080
rect 14971 22052 15016 22080
rect 14599 22049 14611 22052
rect 14553 22043 14611 22049
rect 8754 21972 8760 22024
rect 8812 22012 8818 22024
rect 8959 22015 9017 22021
rect 8959 22012 8971 22015
rect 8812 21984 8971 22012
rect 8812 21972 8818 21984
rect 8959 21981 8971 21984
rect 9005 22012 9017 22015
rect 9122 22012 9128 22024
rect 9005 21984 9128 22012
rect 9005 21981 9017 21984
rect 8959 21975 9017 21981
rect 9122 21972 9128 21984
rect 9180 21972 9186 22024
rect 9766 22012 9772 22024
rect 9727 21984 9772 22012
rect 9766 21972 9772 21984
rect 9824 21972 9830 22024
rect 10502 22012 10508 22024
rect 10463 21984 10508 22012
rect 10502 21972 10508 21984
rect 10560 21972 10566 22024
rect 10594 21972 10600 22024
rect 10652 22012 10658 22024
rect 10689 22015 10747 22021
rect 10689 22012 10701 22015
rect 10652 21984 10701 22012
rect 10652 21972 10658 21984
rect 10689 21981 10701 21984
rect 10735 21981 10747 22015
rect 10689 21975 10747 21981
rect 10873 22015 10931 22021
rect 10873 21981 10885 22015
rect 10919 22012 10931 22015
rect 11054 22012 11060 22024
rect 10919 21984 11060 22012
rect 10919 21981 10931 21984
rect 10873 21975 10931 21981
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 13722 21972 13728 22024
rect 13780 22012 13786 22024
rect 13817 22015 13875 22021
rect 13817 22012 13829 22015
rect 13780 21984 13829 22012
rect 13780 21972 13786 21984
rect 13817 21981 13829 21984
rect 13863 21981 13875 22015
rect 13817 21975 13875 21981
rect 13906 21972 13912 22024
rect 13964 22012 13970 22024
rect 13964 21984 14009 22012
rect 13964 21972 13970 21984
rect 10042 21944 10048 21956
rect 8496 21916 10048 21944
rect 10042 21904 10048 21916
rect 10100 21904 10106 21956
rect 11422 21944 11428 21956
rect 11383 21916 11428 21944
rect 11422 21904 11428 21916
rect 11480 21904 11486 21956
rect 13170 21904 13176 21956
rect 13228 21944 13234 21956
rect 14844 21953 14872 22052
rect 15010 22040 15016 22052
rect 15068 22040 15074 22092
rect 15378 22080 15384 22092
rect 15339 22052 15384 22080
rect 15378 22040 15384 22052
rect 15436 22040 15442 22092
rect 15856 22089 15884 22120
rect 16206 22108 16212 22120
rect 16264 22108 16270 22160
rect 17402 22148 17408 22160
rect 17363 22120 17408 22148
rect 17402 22108 17408 22120
rect 17460 22108 17466 22160
rect 17954 22157 17960 22160
rect 17911 22151 17960 22157
rect 17911 22117 17923 22151
rect 17957 22117 17960 22151
rect 17911 22111 17960 22117
rect 17954 22108 17960 22111
rect 18012 22108 18018 22160
rect 18616 22120 19288 22148
rect 15841 22083 15899 22089
rect 15841 22049 15853 22083
rect 15887 22049 15899 22083
rect 15841 22043 15899 22049
rect 16022 22040 16028 22092
rect 16080 22080 16086 22092
rect 16117 22083 16175 22089
rect 16117 22080 16129 22083
rect 16080 22052 16129 22080
rect 16080 22040 16086 22052
rect 16117 22049 16129 22052
rect 16163 22049 16175 22083
rect 16482 22080 16488 22092
rect 16443 22052 16488 22080
rect 16117 22043 16175 22049
rect 16482 22040 16488 22052
rect 16540 22040 16546 22092
rect 16574 22040 16580 22092
rect 16632 22080 16638 22092
rect 17034 22080 17040 22092
rect 16632 22052 16677 22080
rect 16947 22052 17040 22080
rect 16632 22040 16638 22052
rect 17034 22040 17040 22052
rect 17092 22080 17098 22092
rect 17221 22083 17279 22089
rect 17221 22080 17233 22083
rect 17092 22052 17233 22080
rect 17092 22040 17098 22052
rect 17221 22049 17233 22052
rect 17267 22049 17279 22083
rect 17221 22043 17279 22049
rect 18049 22083 18107 22089
rect 18049 22049 18061 22083
rect 18095 22080 18107 22083
rect 18616 22080 18644 22120
rect 18095 22052 18644 22080
rect 18693 22083 18751 22089
rect 18095 22049 18107 22052
rect 18049 22043 18107 22049
rect 18693 22049 18705 22083
rect 18739 22080 18751 22083
rect 19058 22080 19064 22092
rect 18739 22052 19064 22080
rect 18739 22049 18751 22052
rect 18693 22043 18751 22049
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 19153 22083 19211 22089
rect 19153 22049 19165 22083
rect 19199 22049 19211 22083
rect 19260 22080 19288 22120
rect 20162 22108 20168 22160
rect 20220 22148 20226 22160
rect 22204 22157 22232 22188
rect 22278 22176 22284 22188
rect 22336 22176 22342 22228
rect 20441 22151 20499 22157
rect 20441 22148 20453 22151
rect 20220 22120 20453 22148
rect 20220 22108 20226 22120
rect 20441 22117 20453 22120
rect 20487 22117 20499 22151
rect 20441 22111 20499 22117
rect 22189 22151 22247 22157
rect 22189 22117 22201 22151
rect 22235 22117 22247 22151
rect 22925 22151 22983 22157
rect 22925 22148 22937 22151
rect 22189 22111 22247 22117
rect 22296 22120 22937 22148
rect 19334 22080 19340 22092
rect 19260 22052 19340 22080
rect 19153 22043 19211 22049
rect 18141 22015 18199 22021
rect 18141 21981 18153 22015
rect 18187 22012 18199 22015
rect 18782 22012 18788 22024
rect 18187 21984 18788 22012
rect 18187 21981 18199 21984
rect 18141 21975 18199 21981
rect 18782 21972 18788 21984
rect 18840 21972 18846 22024
rect 19168 22012 19196 22043
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 19426 22040 19432 22092
rect 19484 22080 19490 22092
rect 19521 22083 19579 22089
rect 19521 22080 19533 22083
rect 19484 22052 19533 22080
rect 19484 22040 19490 22052
rect 19521 22049 19533 22052
rect 19567 22049 19579 22083
rect 19521 22043 19579 22049
rect 19610 22040 19616 22092
rect 19668 22080 19674 22092
rect 19889 22083 19947 22089
rect 19889 22080 19901 22083
rect 19668 22052 19901 22080
rect 19668 22040 19674 22052
rect 19889 22049 19901 22052
rect 19935 22049 19947 22083
rect 20070 22080 20076 22092
rect 20031 22052 20076 22080
rect 19889 22043 19947 22049
rect 20070 22040 20076 22052
rect 20128 22040 20134 22092
rect 20254 22080 20260 22092
rect 20215 22052 20260 22080
rect 20254 22040 20260 22052
rect 20312 22040 20318 22092
rect 20806 22080 20812 22092
rect 20767 22052 20812 22080
rect 20806 22040 20812 22052
rect 20864 22040 20870 22092
rect 20898 22040 20904 22092
rect 20956 22080 20962 22092
rect 21082 22080 21088 22092
rect 20956 22052 21001 22080
rect 21043 22052 21088 22080
rect 20956 22040 20962 22052
rect 21082 22040 21088 22052
rect 21140 22040 21146 22092
rect 21450 22080 21456 22092
rect 21411 22052 21456 22080
rect 21450 22040 21456 22052
rect 21508 22040 21514 22092
rect 21634 22080 21640 22092
rect 21595 22052 21640 22080
rect 21634 22040 21640 22052
rect 21692 22040 21698 22092
rect 21818 22080 21824 22092
rect 21779 22052 21824 22080
rect 21818 22040 21824 22052
rect 21876 22040 21882 22092
rect 21910 22040 21916 22092
rect 21968 22080 21974 22092
rect 22296 22080 22324 22120
rect 22925 22117 22937 22120
rect 22971 22117 22983 22151
rect 22925 22111 22983 22117
rect 23106 22080 23112 22092
rect 21968 22052 22324 22080
rect 23067 22052 23112 22080
rect 21968 22040 21974 22052
rect 23106 22040 23112 22052
rect 23164 22040 23170 22092
rect 19242 22012 19248 22024
rect 19168 21984 19248 22012
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 19705 22015 19763 22021
rect 19705 21981 19717 22015
rect 19751 22012 19763 22015
rect 21542 22012 21548 22024
rect 19751 21984 21548 22012
rect 19751 21981 19763 21984
rect 19705 21975 19763 21981
rect 21542 21972 21548 21984
rect 21600 21972 21606 22024
rect 22002 21972 22008 22024
rect 22060 22012 22066 22024
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22060 21984 22385 22012
rect 22060 21972 22066 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 13357 21947 13415 21953
rect 13357 21944 13369 21947
rect 13228 21916 13369 21944
rect 13228 21904 13234 21916
rect 13357 21913 13369 21916
rect 13403 21913 13415 21947
rect 13357 21907 13415 21913
rect 14829 21947 14887 21953
rect 14829 21913 14841 21947
rect 14875 21913 14887 21947
rect 14829 21907 14887 21913
rect 17678 21904 17684 21956
rect 17736 21944 17742 21956
rect 18509 21947 18567 21953
rect 18509 21944 18521 21947
rect 17736 21916 18521 21944
rect 17736 21904 17742 21916
rect 18509 21913 18521 21916
rect 18555 21913 18567 21947
rect 18509 21907 18567 21913
rect 19337 21947 19395 21953
rect 19337 21913 19349 21947
rect 19383 21944 19395 21947
rect 22186 21944 22192 21956
rect 19383 21916 22192 21944
rect 19383 21913 19395 21916
rect 19337 21907 19395 21913
rect 22186 21904 22192 21916
rect 22244 21904 22250 21956
rect 9858 21876 9864 21888
rect 7300 21848 9864 21876
rect 7193 21839 7251 21845
rect 9858 21836 9864 21848
rect 9916 21836 9922 21888
rect 11238 21876 11244 21888
rect 11199 21848 11244 21876
rect 11238 21836 11244 21848
rect 11296 21836 11302 21888
rect 11606 21836 11612 21888
rect 11664 21876 11670 21888
rect 11885 21879 11943 21885
rect 11885 21876 11897 21879
rect 11664 21848 11897 21876
rect 11664 21836 11670 21848
rect 11885 21845 11897 21848
rect 11931 21845 11943 21879
rect 12526 21876 12532 21888
rect 12487 21848 12532 21876
rect 11885 21839 11943 21845
rect 12526 21836 12532 21848
rect 12584 21836 12590 21888
rect 12989 21879 13047 21885
rect 12989 21845 13001 21879
rect 13035 21876 13047 21879
rect 13078 21876 13084 21888
rect 13035 21848 13084 21876
rect 13035 21845 13047 21848
rect 12989 21839 13047 21845
rect 13078 21836 13084 21848
rect 13136 21836 13142 21888
rect 13262 21876 13268 21888
rect 13223 21848 13268 21876
rect 13262 21836 13268 21848
rect 13320 21836 13326 21888
rect 13998 21836 14004 21888
rect 14056 21876 14062 21888
rect 14185 21879 14243 21885
rect 14185 21876 14197 21879
rect 14056 21848 14197 21876
rect 14056 21836 14062 21848
rect 14185 21845 14197 21848
rect 14231 21845 14243 21879
rect 14734 21876 14740 21888
rect 14695 21848 14740 21876
rect 14185 21839 14243 21845
rect 14734 21836 14740 21848
rect 14792 21836 14798 21888
rect 15197 21879 15255 21885
rect 15197 21845 15209 21879
rect 15243 21876 15255 21879
rect 15286 21876 15292 21888
rect 15243 21848 15292 21876
rect 15243 21845 15255 21848
rect 15197 21839 15255 21845
rect 15286 21836 15292 21848
rect 15344 21836 15350 21888
rect 15470 21836 15476 21888
rect 15528 21876 15534 21888
rect 15933 21879 15991 21885
rect 15933 21876 15945 21879
rect 15528 21848 15945 21876
rect 15528 21836 15534 21848
rect 15933 21845 15945 21848
rect 15979 21845 15991 21879
rect 16758 21876 16764 21888
rect 16719 21848 16764 21876
rect 15933 21839 15991 21845
rect 16758 21836 16764 21848
rect 16816 21836 16822 21888
rect 16853 21879 16911 21885
rect 16853 21845 16865 21879
rect 16899 21876 16911 21879
rect 16942 21876 16948 21888
rect 16899 21848 16948 21876
rect 16899 21845 16911 21848
rect 16853 21839 16911 21845
rect 16942 21836 16948 21848
rect 17000 21836 17006 21888
rect 18966 21836 18972 21888
rect 19024 21876 19030 21888
rect 20625 21879 20683 21885
rect 20625 21876 20637 21879
rect 19024 21848 20637 21876
rect 19024 21836 19030 21848
rect 20625 21845 20637 21848
rect 20671 21845 20683 21879
rect 20625 21839 20683 21845
rect 21913 21879 21971 21885
rect 21913 21845 21925 21879
rect 21959 21876 21971 21879
rect 22094 21876 22100 21888
rect 21959 21848 22100 21876
rect 21959 21845 21971 21848
rect 21913 21839 21971 21845
rect 22094 21836 22100 21848
rect 22152 21836 22158 21888
rect 1104 21786 23460 21808
rect 1104 21734 4714 21786
rect 4766 21734 4778 21786
rect 4830 21734 4842 21786
rect 4894 21734 4906 21786
rect 4958 21734 12178 21786
rect 12230 21734 12242 21786
rect 12294 21734 12306 21786
rect 12358 21734 12370 21786
rect 12422 21734 19642 21786
rect 19694 21734 19706 21786
rect 19758 21734 19770 21786
rect 19822 21734 19834 21786
rect 19886 21734 23460 21786
rect 1104 21712 23460 21734
rect 1578 21632 1584 21684
rect 1636 21672 1642 21684
rect 1857 21675 1915 21681
rect 1857 21672 1869 21675
rect 1636 21644 1869 21672
rect 1636 21632 1642 21644
rect 1857 21641 1869 21644
rect 1903 21641 1915 21675
rect 1857 21635 1915 21641
rect 1946 21632 1952 21684
rect 2004 21672 2010 21684
rect 2133 21675 2191 21681
rect 2133 21672 2145 21675
rect 2004 21644 2145 21672
rect 2004 21632 2010 21644
rect 2133 21641 2145 21644
rect 2179 21641 2191 21675
rect 2133 21635 2191 21641
rect 3326 21632 3332 21684
rect 3384 21672 3390 21684
rect 4065 21675 4123 21681
rect 4065 21672 4077 21675
rect 3384 21644 4077 21672
rect 3384 21632 3390 21644
rect 4065 21641 4077 21644
rect 4111 21641 4123 21675
rect 4065 21635 4123 21641
rect 5994 21632 6000 21684
rect 6052 21672 6058 21684
rect 6457 21675 6515 21681
rect 6457 21672 6469 21675
rect 6052 21644 6469 21672
rect 6052 21632 6058 21644
rect 6457 21641 6469 21644
rect 6503 21641 6515 21675
rect 6730 21672 6736 21684
rect 6691 21644 6736 21672
rect 6457 21635 6515 21641
rect 6730 21632 6736 21644
rect 6788 21632 6794 21684
rect 6917 21675 6975 21681
rect 6917 21641 6929 21675
rect 6963 21672 6975 21675
rect 7926 21672 7932 21684
rect 6963 21644 7932 21672
rect 6963 21641 6975 21644
rect 6917 21635 6975 21641
rect 7926 21632 7932 21644
rect 7984 21632 7990 21684
rect 8110 21632 8116 21684
rect 8168 21672 8174 21684
rect 9217 21675 9275 21681
rect 9217 21672 9229 21675
rect 8168 21644 9229 21672
rect 8168 21632 8174 21644
rect 9217 21641 9229 21644
rect 9263 21641 9275 21675
rect 9217 21635 9275 21641
rect 9401 21675 9459 21681
rect 9401 21641 9413 21675
rect 9447 21672 9459 21675
rect 9858 21672 9864 21684
rect 9447 21644 9864 21672
rect 9447 21641 9459 21644
rect 9401 21635 9459 21641
rect 9858 21632 9864 21644
rect 9916 21672 9922 21684
rect 10594 21672 10600 21684
rect 9916 21644 10600 21672
rect 9916 21632 9922 21644
rect 10594 21632 10600 21644
rect 10652 21632 10658 21684
rect 10965 21675 11023 21681
rect 10965 21641 10977 21675
rect 11011 21672 11023 21675
rect 11790 21672 11796 21684
rect 11011 21644 11796 21672
rect 11011 21641 11023 21644
rect 10965 21635 11023 21641
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 12986 21632 12992 21684
rect 13044 21672 13050 21684
rect 13044 21644 14320 21672
rect 13044 21632 13050 21644
rect 2498 21604 2504 21616
rect 2056 21576 2504 21604
rect 1578 21468 1584 21480
rect 1539 21440 1584 21468
rect 1578 21428 1584 21440
rect 1636 21468 1642 21480
rect 2056 21477 2084 21576
rect 2498 21564 2504 21576
rect 2556 21564 2562 21616
rect 3973 21607 4031 21613
rect 3973 21573 3985 21607
rect 4019 21604 4031 21607
rect 4154 21604 4160 21616
rect 4019 21576 4160 21604
rect 4019 21573 4031 21576
rect 3973 21567 4031 21573
rect 4154 21564 4160 21576
rect 4212 21564 4218 21616
rect 9030 21604 9036 21616
rect 8312 21576 9036 21604
rect 2130 21496 2136 21548
rect 2188 21536 2194 21548
rect 5905 21539 5963 21545
rect 2188 21508 2636 21536
rect 2188 21496 2194 21508
rect 1673 21471 1731 21477
rect 1673 21468 1685 21471
rect 1636 21440 1685 21468
rect 1636 21428 1642 21440
rect 1673 21437 1685 21440
rect 1719 21437 1731 21471
rect 1673 21431 1731 21437
rect 2041 21471 2099 21477
rect 2041 21437 2053 21471
rect 2087 21437 2099 21471
rect 2041 21431 2099 21437
rect 2317 21471 2375 21477
rect 2317 21437 2329 21471
rect 2363 21468 2375 21471
rect 2406 21468 2412 21480
rect 2363 21440 2412 21468
rect 2363 21437 2375 21440
rect 2317 21431 2375 21437
rect 2406 21428 2412 21440
rect 2464 21428 2470 21480
rect 2608 21477 2636 21508
rect 5905 21505 5917 21539
rect 5951 21536 5963 21539
rect 6914 21536 6920 21548
rect 5951 21508 6920 21536
rect 5951 21505 5963 21508
rect 5905 21499 5963 21505
rect 6914 21496 6920 21508
rect 6972 21496 6978 21548
rect 8312 21545 8340 21576
rect 9030 21564 9036 21576
rect 9088 21564 9094 21616
rect 10870 21564 10876 21616
rect 10928 21604 10934 21616
rect 11333 21607 11391 21613
rect 11333 21604 11345 21607
rect 10928 21576 11345 21604
rect 10928 21564 10934 21576
rect 11333 21573 11345 21576
rect 11379 21573 11391 21607
rect 11333 21567 11391 21573
rect 8297 21539 8355 21545
rect 8297 21505 8309 21539
rect 8343 21505 8355 21539
rect 8297 21499 8355 21505
rect 8570 21496 8576 21548
rect 8628 21536 8634 21548
rect 10781 21539 10839 21545
rect 8628 21508 9674 21536
rect 8628 21496 8634 21508
rect 2593 21471 2651 21477
rect 2593 21437 2605 21471
rect 2639 21468 2651 21471
rect 4246 21468 4252 21480
rect 2639 21440 3556 21468
rect 4207 21440 4252 21468
rect 2639 21437 2651 21440
rect 2593 21431 2651 21437
rect 2860 21403 2918 21409
rect 2860 21369 2872 21403
rect 2906 21400 2918 21403
rect 3418 21400 3424 21412
rect 2906 21372 3424 21400
rect 2906 21369 2918 21372
rect 2860 21363 2918 21369
rect 3418 21360 3424 21372
rect 3476 21360 3482 21412
rect 3528 21400 3556 21440
rect 4246 21428 4252 21440
rect 4304 21428 4310 21480
rect 4430 21468 4436 21480
rect 4391 21440 4436 21468
rect 4430 21428 4436 21440
rect 4488 21428 4494 21480
rect 4522 21428 4528 21480
rect 4580 21468 4586 21480
rect 6638 21468 6644 21480
rect 4580 21440 6224 21468
rect 6599 21440 6644 21468
rect 4580 21428 4586 21440
rect 4448 21400 4476 21428
rect 3528 21372 4476 21400
rect 4700 21403 4758 21409
rect 4700 21369 4712 21403
rect 4746 21400 4758 21403
rect 5258 21400 5264 21412
rect 4746 21372 5264 21400
rect 4746 21369 4758 21372
rect 4700 21363 4758 21369
rect 5258 21360 5264 21372
rect 5316 21400 5322 21412
rect 6089 21403 6147 21409
rect 6089 21400 6101 21403
rect 5316 21372 6101 21400
rect 5316 21360 5322 21372
rect 6089 21369 6101 21372
rect 6135 21369 6147 21403
rect 6089 21363 6147 21369
rect 5810 21332 5816 21344
rect 5771 21304 5816 21332
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 6196 21332 6224 21440
rect 6638 21428 6644 21440
rect 6696 21428 6702 21480
rect 8041 21471 8099 21477
rect 8041 21437 8053 21471
rect 8087 21468 8099 21471
rect 8386 21468 8392 21480
rect 8087 21440 8392 21468
rect 8087 21437 8099 21440
rect 8041 21431 8099 21437
rect 8386 21428 8392 21440
rect 8444 21428 8450 21480
rect 8481 21471 8539 21477
rect 8481 21437 8493 21471
rect 8527 21468 8539 21471
rect 8754 21468 8760 21480
rect 8527 21440 8760 21468
rect 8527 21437 8539 21440
rect 8481 21431 8539 21437
rect 8754 21428 8760 21440
rect 8812 21428 8818 21480
rect 9646 21468 9674 21508
rect 10781 21505 10793 21539
rect 10827 21536 10839 21539
rect 10962 21536 10968 21548
rect 10827 21508 10968 21536
rect 10827 21505 10839 21508
rect 10781 21499 10839 21505
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 11606 21536 11612 21548
rect 11072 21508 11612 21536
rect 10686 21468 10692 21480
rect 9646 21440 10692 21468
rect 10686 21428 10692 21440
rect 10744 21428 10750 21480
rect 11072 21477 11100 21508
rect 11606 21496 11612 21508
rect 11664 21496 11670 21548
rect 11698 21496 11704 21548
rect 11756 21536 11762 21548
rect 11793 21539 11851 21545
rect 11793 21536 11805 21539
rect 11756 21508 11805 21536
rect 11756 21496 11762 21508
rect 11793 21505 11805 21508
rect 11839 21505 11851 21539
rect 14292 21536 14320 21644
rect 15378 21632 15384 21684
rect 15436 21672 15442 21684
rect 16117 21675 16175 21681
rect 16117 21672 16129 21675
rect 15436 21644 15884 21672
rect 15436 21632 15442 21644
rect 14642 21604 14648 21616
rect 14603 21576 14648 21604
rect 14642 21564 14648 21576
rect 14700 21564 14706 21616
rect 15856 21604 15884 21644
rect 16040 21644 16129 21672
rect 16040 21604 16068 21644
rect 16117 21641 16129 21644
rect 16163 21672 16175 21675
rect 16390 21672 16396 21684
rect 16163 21644 16396 21672
rect 16163 21641 16175 21644
rect 16117 21635 16175 21641
rect 16390 21632 16396 21644
rect 16448 21632 16454 21684
rect 16574 21632 16580 21684
rect 16632 21672 16638 21684
rect 16761 21675 16819 21681
rect 16761 21672 16773 21675
rect 16632 21644 16773 21672
rect 16632 21632 16638 21644
rect 16761 21641 16773 21644
rect 16807 21672 16819 21675
rect 18322 21672 18328 21684
rect 16807 21644 18328 21672
rect 16807 21641 16819 21644
rect 16761 21635 16819 21641
rect 18322 21632 18328 21644
rect 18380 21632 18386 21684
rect 19429 21675 19487 21681
rect 19429 21641 19441 21675
rect 19475 21672 19487 21675
rect 22830 21672 22836 21684
rect 19475 21644 22836 21672
rect 19475 21641 19487 21644
rect 19429 21635 19487 21641
rect 22830 21632 22836 21644
rect 22888 21632 22894 21684
rect 16206 21604 16212 21616
rect 15856 21576 16068 21604
rect 16167 21576 16212 21604
rect 16206 21564 16212 21576
rect 16264 21564 16270 21616
rect 18046 21564 18052 21616
rect 18104 21604 18110 21616
rect 19705 21607 19763 21613
rect 19705 21604 19717 21607
rect 18104 21576 19717 21604
rect 18104 21564 18110 21576
rect 19705 21573 19717 21576
rect 19751 21604 19763 21607
rect 20070 21604 20076 21616
rect 19751 21576 20076 21604
rect 19751 21573 19763 21576
rect 19705 21567 19763 21573
rect 20070 21564 20076 21576
rect 20128 21564 20134 21616
rect 22741 21607 22799 21613
rect 22741 21573 22753 21607
rect 22787 21604 22799 21607
rect 23474 21604 23480 21616
rect 22787 21576 23480 21604
rect 22787 21573 22799 21576
rect 22741 21567 22799 21573
rect 23474 21564 23480 21576
rect 23532 21564 23538 21616
rect 14292 21508 14872 21536
rect 11793 21499 11851 21505
rect 11049 21471 11107 21477
rect 11049 21437 11061 21471
rect 11095 21437 11107 21471
rect 11049 21431 11107 21437
rect 11330 21428 11336 21480
rect 11388 21468 11394 21480
rect 11517 21471 11575 21477
rect 11517 21468 11529 21471
rect 11388 21440 11529 21468
rect 11388 21428 11394 21440
rect 11517 21437 11529 21440
rect 11563 21437 11575 21471
rect 12342 21468 12348 21480
rect 11517 21431 11575 21437
rect 11624 21440 12348 21468
rect 6273 21403 6331 21409
rect 6273 21369 6285 21403
rect 6319 21400 6331 21403
rect 7834 21400 7840 21412
rect 6319 21372 7840 21400
rect 6319 21369 6331 21372
rect 6273 21363 6331 21369
rect 7834 21360 7840 21372
rect 7892 21360 7898 21412
rect 8938 21360 8944 21412
rect 8996 21400 9002 21412
rect 8996 21372 9041 21400
rect 8996 21360 9002 21372
rect 9122 21360 9128 21412
rect 9180 21400 9186 21412
rect 10410 21400 10416 21412
rect 9180 21372 10416 21400
rect 9180 21360 9186 21372
rect 10410 21360 10416 21372
rect 10468 21360 10474 21412
rect 10536 21403 10594 21409
rect 10536 21369 10548 21403
rect 10582 21400 10594 21403
rect 10962 21400 10968 21412
rect 10582 21372 10968 21400
rect 10582 21369 10594 21372
rect 10536 21363 10594 21369
rect 10962 21360 10968 21372
rect 11020 21360 11026 21412
rect 11624 21400 11652 21440
rect 12342 21428 12348 21440
rect 12400 21428 12406 21480
rect 12894 21428 12900 21480
rect 12952 21468 12958 21480
rect 13265 21471 13323 21477
rect 13265 21468 13277 21471
rect 12952 21440 13277 21468
rect 12952 21428 12958 21440
rect 13265 21437 13277 21440
rect 13311 21437 13323 21471
rect 13265 21431 13323 21437
rect 14090 21428 14096 21480
rect 14148 21468 14154 21480
rect 14737 21471 14795 21477
rect 14737 21468 14749 21471
rect 14148 21440 14749 21468
rect 14148 21428 14154 21440
rect 14737 21437 14749 21440
rect 14783 21437 14795 21471
rect 14844 21468 14872 21508
rect 16022 21496 16028 21548
rect 16080 21536 16086 21548
rect 16080 21508 16528 21536
rect 16080 21496 16086 21508
rect 14844 21440 15240 21468
rect 14737 21431 14795 21437
rect 12066 21409 12072 21412
rect 12060 21400 12072 21409
rect 11072 21372 11652 21400
rect 12027 21372 12072 21400
rect 11072 21332 11100 21372
rect 12060 21363 12072 21372
rect 12066 21360 12072 21363
rect 12124 21360 12130 21412
rect 13354 21400 13360 21412
rect 13188 21372 13360 21400
rect 6196 21304 11100 21332
rect 11241 21335 11299 21341
rect 11241 21301 11253 21335
rect 11287 21332 11299 21335
rect 11606 21332 11612 21344
rect 11287 21304 11612 21332
rect 11287 21301 11299 21304
rect 11241 21295 11299 21301
rect 11606 21292 11612 21304
rect 11664 21292 11670 21344
rect 11701 21335 11759 21341
rect 11701 21301 11713 21335
rect 11747 21332 11759 21335
rect 12894 21332 12900 21344
rect 11747 21304 12900 21332
rect 11747 21301 11759 21304
rect 11701 21295 11759 21301
rect 12894 21292 12900 21304
rect 12952 21292 12958 21344
rect 13188 21341 13216 21372
rect 13354 21360 13360 21372
rect 13412 21400 13418 21412
rect 13510 21403 13568 21409
rect 13510 21400 13522 21403
rect 13412 21372 13522 21400
rect 13412 21360 13418 21372
rect 13510 21369 13522 21372
rect 13556 21369 13568 21403
rect 13510 21363 13568 21369
rect 14274 21360 14280 21412
rect 14332 21400 14338 21412
rect 14982 21403 15040 21409
rect 14982 21400 14994 21403
rect 14332 21372 14994 21400
rect 14332 21360 14338 21372
rect 14982 21369 14994 21372
rect 15028 21400 15040 21403
rect 15102 21400 15108 21412
rect 15028 21372 15108 21400
rect 15028 21369 15040 21372
rect 14982 21363 15040 21369
rect 15102 21360 15108 21372
rect 15160 21360 15166 21412
rect 15212 21400 15240 21440
rect 15286 21428 15292 21480
rect 15344 21468 15350 21480
rect 16393 21471 16451 21477
rect 16393 21468 16405 21471
rect 15344 21440 16405 21468
rect 15344 21428 15350 21440
rect 16393 21437 16405 21440
rect 16439 21437 16451 21471
rect 16500 21468 16528 21508
rect 16758 21496 16764 21548
rect 16816 21536 16822 21548
rect 16816 21508 17080 21536
rect 16816 21496 16822 21508
rect 16942 21468 16948 21480
rect 16500 21440 16948 21468
rect 16393 21431 16451 21437
rect 16942 21428 16948 21440
rect 17000 21428 17006 21480
rect 17052 21468 17080 21508
rect 18690 21496 18696 21548
rect 18748 21536 18754 21548
rect 18785 21539 18843 21545
rect 18785 21536 18797 21539
rect 18748 21508 18797 21536
rect 18748 21496 18754 21508
rect 18785 21505 18797 21508
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 19242 21496 19248 21548
rect 19300 21536 19306 21548
rect 19889 21539 19947 21545
rect 19889 21536 19901 21539
rect 19300 21508 19901 21536
rect 19300 21496 19306 21508
rect 19889 21505 19901 21508
rect 19935 21505 19947 21539
rect 23106 21536 23112 21548
rect 23067 21508 23112 21536
rect 19889 21499 19947 21505
rect 23106 21496 23112 21508
rect 23164 21496 23170 21548
rect 18509 21471 18567 21477
rect 18509 21468 18521 21471
rect 17052 21440 18521 21468
rect 18509 21437 18521 21440
rect 18555 21437 18567 21471
rect 18509 21431 18567 21437
rect 18598 21428 18604 21480
rect 18656 21468 18662 21480
rect 20073 21471 20131 21477
rect 20073 21468 20085 21471
rect 18656 21440 20085 21468
rect 18656 21428 18662 21440
rect 20073 21437 20085 21440
rect 20119 21468 20131 21471
rect 20162 21468 20168 21480
rect 20119 21440 20168 21468
rect 20119 21437 20131 21440
rect 20073 21431 20131 21437
rect 20162 21428 20168 21440
rect 20220 21428 20226 21480
rect 21634 21428 21640 21480
rect 21692 21468 21698 21480
rect 22925 21471 22983 21477
rect 22925 21468 22937 21471
rect 21692 21440 22937 21468
rect 21692 21428 21698 21440
rect 22925 21437 22937 21440
rect 22971 21437 22983 21471
rect 22925 21431 22983 21437
rect 17218 21409 17224 21412
rect 16485 21403 16543 21409
rect 16485 21400 16497 21403
rect 15212 21372 16497 21400
rect 16485 21369 16497 21372
rect 16531 21369 16543 21403
rect 17212 21400 17224 21409
rect 17179 21372 17224 21400
rect 16485 21363 16543 21369
rect 17212 21363 17224 21372
rect 17218 21360 17224 21363
rect 17276 21360 17282 21412
rect 17310 21360 17316 21412
rect 17368 21400 17374 21412
rect 17368 21372 19012 21400
rect 17368 21360 17374 21372
rect 13173 21335 13231 21341
rect 13173 21301 13185 21335
rect 13219 21301 13231 21335
rect 13173 21295 13231 21301
rect 18325 21335 18383 21341
rect 18325 21301 18337 21335
rect 18371 21332 18383 21335
rect 18874 21332 18880 21344
rect 18371 21304 18880 21332
rect 18371 21301 18383 21304
rect 18325 21295 18383 21301
rect 18874 21292 18880 21304
rect 18932 21292 18938 21344
rect 18984 21332 19012 21372
rect 19150 21360 19156 21412
rect 19208 21400 19214 21412
rect 19337 21403 19395 21409
rect 19337 21400 19349 21403
rect 19208 21372 19349 21400
rect 19208 21360 19214 21372
rect 19337 21369 19349 21372
rect 19383 21369 19395 21403
rect 22557 21403 22615 21409
rect 22557 21400 22569 21403
rect 19337 21363 19395 21369
rect 22066 21372 22569 21400
rect 20717 21335 20775 21341
rect 20717 21332 20729 21335
rect 18984 21304 20729 21332
rect 20717 21301 20729 21304
rect 20763 21332 20775 21335
rect 21082 21332 21088 21344
rect 20763 21304 21088 21332
rect 20763 21301 20775 21304
rect 20717 21295 20775 21301
rect 21082 21292 21088 21304
rect 21140 21292 21146 21344
rect 21358 21332 21364 21344
rect 21319 21304 21364 21332
rect 21358 21292 21364 21304
rect 21416 21292 21422 21344
rect 21542 21292 21548 21344
rect 21600 21332 21606 21344
rect 21913 21335 21971 21341
rect 21913 21332 21925 21335
rect 21600 21304 21925 21332
rect 21600 21292 21606 21304
rect 21913 21301 21925 21304
rect 21959 21332 21971 21335
rect 22066 21332 22094 21372
rect 22557 21369 22569 21372
rect 22603 21369 22615 21403
rect 22557 21363 22615 21369
rect 22186 21332 22192 21344
rect 21959 21304 22094 21332
rect 22147 21304 22192 21332
rect 21959 21301 21971 21304
rect 21913 21295 21971 21301
rect 22186 21292 22192 21304
rect 22244 21292 22250 21344
rect 1104 21242 23460 21264
rect 1104 21190 8446 21242
rect 8498 21190 8510 21242
rect 8562 21190 8574 21242
rect 8626 21190 8638 21242
rect 8690 21190 15910 21242
rect 15962 21190 15974 21242
rect 16026 21190 16038 21242
rect 16090 21190 16102 21242
rect 16154 21190 23460 21242
rect 1104 21168 23460 21190
rect 1949 21131 2007 21137
rect 1949 21097 1961 21131
rect 1995 21128 2007 21131
rect 2314 21128 2320 21140
rect 1995 21100 2320 21128
rect 1995 21097 2007 21100
rect 1949 21091 2007 21097
rect 2314 21088 2320 21100
rect 2372 21088 2378 21140
rect 2682 21088 2688 21140
rect 2740 21128 2746 21140
rect 3513 21131 3571 21137
rect 3513 21128 3525 21131
rect 2740 21100 3525 21128
rect 2740 21088 2746 21100
rect 3513 21097 3525 21100
rect 3559 21097 3571 21131
rect 5258 21128 5264 21140
rect 5219 21100 5264 21128
rect 3513 21091 3571 21097
rect 5258 21088 5264 21100
rect 5316 21088 5322 21140
rect 5350 21088 5356 21140
rect 5408 21128 5414 21140
rect 8297 21131 8355 21137
rect 5408 21100 8064 21128
rect 5408 21088 5414 21100
rect 1489 21063 1547 21069
rect 1489 21029 1501 21063
rect 1535 21060 1547 21063
rect 2590 21060 2596 21072
rect 1535 21032 2596 21060
rect 1535 21029 1547 21032
rect 1489 21023 1547 21029
rect 2590 21020 2596 21032
rect 2648 21020 2654 21072
rect 4154 21069 4160 21072
rect 4148 21060 4160 21069
rect 4115 21032 4160 21060
rect 4148 21023 4160 21032
rect 4154 21020 4160 21023
rect 4212 21020 4218 21072
rect 5620 21063 5678 21069
rect 5620 21029 5632 21063
rect 5666 21060 5678 21063
rect 5810 21060 5816 21072
rect 5666 21032 5816 21060
rect 5666 21029 5678 21032
rect 5620 21023 5678 21029
rect 5810 21020 5816 21032
rect 5868 21020 5874 21072
rect 8036 21060 8064 21100
rect 8297 21097 8309 21131
rect 8343 21128 8355 21131
rect 8573 21131 8631 21137
rect 8343 21100 8432 21128
rect 8343 21097 8355 21100
rect 8297 21091 8355 21097
rect 8404 21072 8432 21100
rect 8573 21097 8585 21131
rect 8619 21128 8631 21131
rect 8754 21128 8760 21140
rect 8619 21100 8760 21128
rect 8619 21097 8631 21100
rect 8573 21091 8631 21097
rect 8754 21088 8760 21100
rect 8812 21088 8818 21140
rect 8846 21088 8852 21140
rect 8904 21128 8910 21140
rect 9125 21131 9183 21137
rect 9125 21128 9137 21131
rect 8904 21100 9137 21128
rect 8904 21088 8910 21100
rect 9125 21097 9137 21100
rect 9171 21097 9183 21131
rect 9125 21091 9183 21097
rect 9306 21088 9312 21140
rect 9364 21128 9370 21140
rect 9364 21100 9720 21128
rect 9364 21088 9370 21100
rect 8036 21032 8340 21060
rect 1765 20995 1823 21001
rect 1765 20992 1777 20995
rect 1688 20964 1777 20992
rect 1688 20868 1716 20964
rect 1765 20961 1777 20964
rect 1811 20961 1823 20995
rect 1765 20955 1823 20961
rect 2041 20995 2099 21001
rect 2041 20961 2053 20995
rect 2087 20992 2099 20995
rect 2130 20992 2136 21004
rect 2087 20964 2136 20992
rect 2087 20961 2099 20964
rect 2041 20955 2099 20961
rect 2130 20952 2136 20964
rect 2188 20952 2194 21004
rect 2308 20995 2366 21001
rect 2308 20961 2320 20995
rect 2354 20992 2366 20995
rect 2866 20992 2872 21004
rect 2354 20964 2872 20992
rect 2354 20961 2366 20964
rect 2308 20955 2366 20961
rect 2866 20952 2872 20964
rect 2924 20952 2930 21004
rect 3694 20992 3700 21004
rect 3655 20964 3700 20992
rect 3694 20952 3700 20964
rect 3752 20952 3758 21004
rect 3881 20995 3939 21001
rect 3881 20961 3893 20995
rect 3927 20992 3939 20995
rect 4430 20992 4436 21004
rect 3927 20964 4436 20992
rect 3927 20961 3939 20964
rect 3881 20955 3939 20961
rect 4430 20952 4436 20964
rect 4488 20952 4494 21004
rect 5353 20995 5411 21001
rect 5353 20961 5365 20995
rect 5399 20992 5411 20995
rect 5399 20964 6684 20992
rect 5399 20961 5411 20964
rect 5353 20955 5411 20961
rect 6656 20936 6684 20964
rect 6730 20952 6736 21004
rect 6788 20992 6794 21004
rect 7081 20995 7139 21001
rect 7081 20992 7093 20995
rect 6788 20964 7093 20992
rect 6788 20952 6794 20964
rect 7081 20961 7093 20964
rect 7127 20961 7139 20995
rect 7081 20955 7139 20961
rect 6638 20884 6644 20936
rect 6696 20924 6702 20936
rect 6825 20927 6883 20933
rect 6825 20924 6837 20927
rect 6696 20896 6837 20924
rect 6696 20884 6702 20896
rect 6825 20893 6837 20896
rect 6871 20893 6883 20927
rect 6825 20887 6883 20893
rect 1670 20856 1676 20868
rect 1631 20828 1676 20856
rect 1670 20816 1676 20828
rect 1728 20816 1734 20868
rect 3418 20856 3424 20868
rect 3379 20828 3424 20856
rect 3418 20816 3424 20828
rect 3476 20816 3482 20868
rect 8312 20856 8340 21032
rect 8386 21020 8392 21072
rect 8444 21020 8450 21072
rect 8864 21060 8892 21088
rect 9582 21069 9588 21072
rect 9576 21060 9588 21069
rect 8496 21032 8892 21060
rect 9543 21032 9588 21060
rect 8496 21001 8524 21032
rect 9576 21023 9588 21032
rect 9582 21020 9588 21023
rect 9640 21020 9646 21072
rect 9692 21060 9720 21100
rect 9766 21088 9772 21140
rect 9824 21128 9830 21140
rect 10781 21131 10839 21137
rect 10781 21128 10793 21131
rect 9824 21100 10793 21128
rect 9824 21088 9830 21100
rect 10781 21097 10793 21100
rect 10827 21097 10839 21131
rect 11054 21128 11060 21140
rect 11015 21100 11060 21128
rect 10781 21091 10839 21097
rect 11054 21088 11060 21100
rect 11112 21088 11118 21140
rect 11517 21131 11575 21137
rect 11517 21097 11529 21131
rect 11563 21097 11575 21131
rect 11517 21091 11575 21097
rect 11330 21060 11336 21072
rect 9692 21032 11336 21060
rect 11330 21020 11336 21032
rect 11388 21020 11394 21072
rect 11532 21060 11560 21091
rect 13354 21088 13360 21140
rect 13412 21128 13418 21140
rect 13722 21128 13728 21140
rect 13412 21100 13457 21128
rect 13683 21100 13728 21128
rect 13412 21088 13418 21100
rect 13722 21088 13728 21100
rect 13780 21088 13786 21140
rect 13906 21128 13912 21140
rect 13867 21100 13912 21128
rect 13906 21088 13912 21100
rect 13964 21088 13970 21140
rect 14090 21088 14096 21140
rect 14148 21128 14154 21140
rect 14148 21100 15056 21128
rect 14148 21088 14154 21100
rect 12066 21060 12072 21072
rect 11532 21032 12072 21060
rect 12066 21020 12072 21032
rect 12124 21060 12130 21072
rect 13265 21063 13323 21069
rect 12124 21032 13032 21060
rect 12124 21020 12130 21032
rect 8481 20995 8539 21001
rect 8481 20961 8493 20995
rect 8527 20961 8539 20995
rect 8481 20955 8539 20961
rect 8757 20995 8815 21001
rect 8757 20961 8769 20995
rect 8803 20992 8815 20995
rect 10502 20992 10508 21004
rect 8803 20964 8837 20992
rect 8956 20964 10508 20992
rect 8803 20961 8815 20964
rect 8757 20955 8815 20961
rect 8386 20884 8392 20936
rect 8444 20924 8450 20936
rect 8772 20924 8800 20955
rect 8849 20927 8907 20933
rect 8849 20924 8861 20927
rect 8444 20896 8861 20924
rect 8444 20884 8450 20896
rect 8849 20893 8861 20896
rect 8895 20893 8907 20927
rect 8849 20887 8907 20893
rect 8956 20856 8984 20964
rect 10502 20952 10508 20964
rect 10560 20992 10566 21004
rect 12342 20992 12348 21004
rect 10560 20964 12348 20992
rect 10560 20952 10566 20964
rect 12342 20952 12348 20964
rect 12400 20952 12406 21004
rect 12618 20952 12624 21004
rect 12676 21001 12682 21004
rect 12676 20992 12688 21001
rect 12894 20992 12900 21004
rect 12676 20964 12721 20992
rect 12855 20964 12900 20992
rect 12676 20955 12688 20964
rect 12676 20952 12682 20955
rect 12894 20952 12900 20964
rect 12952 20952 12958 21004
rect 13004 20992 13032 21032
rect 13265 21029 13277 21063
rect 13311 21029 13323 21063
rect 13998 21060 14004 21072
rect 13959 21032 14004 21060
rect 13265 21023 13323 21029
rect 13280 20992 13308 21023
rect 13998 21020 14004 21032
rect 14056 21020 14062 21072
rect 14642 21069 14648 21072
rect 14636 21060 14648 21069
rect 14603 21032 14648 21060
rect 14636 21023 14648 21032
rect 14642 21020 14648 21023
rect 14700 21020 14706 21072
rect 15028 21060 15056 21100
rect 15102 21088 15108 21140
rect 15160 21128 15166 21140
rect 15749 21131 15807 21137
rect 15749 21128 15761 21131
rect 15160 21100 15761 21128
rect 15160 21088 15166 21100
rect 15749 21097 15761 21100
rect 15795 21097 15807 21131
rect 18598 21128 18604 21140
rect 15749 21091 15807 21097
rect 15856 21100 18604 21128
rect 15856 21072 15884 21100
rect 18598 21088 18604 21100
rect 18656 21088 18662 21140
rect 18782 21128 18788 21140
rect 18743 21100 18788 21128
rect 18782 21088 18788 21100
rect 18840 21088 18846 21140
rect 19058 21128 19064 21140
rect 19019 21100 19064 21128
rect 19058 21088 19064 21100
rect 19116 21088 19122 21140
rect 19150 21088 19156 21140
rect 19208 21128 19214 21140
rect 19613 21131 19671 21137
rect 19613 21128 19625 21131
rect 19208 21100 19625 21128
rect 19208 21088 19214 21100
rect 19613 21097 19625 21100
rect 19659 21097 19671 21131
rect 19613 21091 19671 21097
rect 21177 21131 21235 21137
rect 21177 21097 21189 21131
rect 21223 21128 21235 21131
rect 21450 21128 21456 21140
rect 21223 21100 21456 21128
rect 21223 21097 21235 21100
rect 21177 21091 21235 21097
rect 21450 21088 21456 21100
rect 21508 21088 21514 21140
rect 21729 21131 21787 21137
rect 21729 21097 21741 21131
rect 21775 21128 21787 21131
rect 22094 21128 22100 21140
rect 21775 21100 22100 21128
rect 21775 21097 21787 21100
rect 21729 21091 21787 21097
rect 22094 21088 22100 21100
rect 22152 21088 22158 21140
rect 22281 21131 22339 21137
rect 22281 21097 22293 21131
rect 22327 21128 22339 21131
rect 24118 21128 24124 21140
rect 22327 21100 24124 21128
rect 22327 21097 22339 21100
rect 22281 21091 22339 21097
rect 24118 21088 24124 21100
rect 24176 21088 24182 21140
rect 15286 21060 15292 21072
rect 15028 21032 15292 21060
rect 15286 21020 15292 21032
rect 15344 21060 15350 21072
rect 15654 21060 15660 21072
rect 15344 21032 15660 21060
rect 15344 21020 15350 21032
rect 15654 21020 15660 21032
rect 15712 21020 15718 21072
rect 15838 21020 15844 21072
rect 15896 21020 15902 21072
rect 16108 21063 16166 21069
rect 16108 21029 16120 21063
rect 16154 21060 16166 21063
rect 16390 21060 16396 21072
rect 16154 21032 16396 21060
rect 16154 21029 16166 21032
rect 16108 21023 16166 21029
rect 16390 21020 16396 21032
rect 16448 21020 16454 21072
rect 19426 21060 19432 21072
rect 16500 21032 19432 21060
rect 13004 20964 13308 20992
rect 14458 20952 14464 21004
rect 14516 20992 14522 21004
rect 16500 20992 16528 21032
rect 19426 21020 19432 21032
rect 19484 21020 19490 21072
rect 21008 21032 21772 21060
rect 14516 20964 16528 20992
rect 17580 20995 17638 21001
rect 14516 20952 14522 20964
rect 17580 20961 17592 20995
rect 17626 20992 17638 20995
rect 18874 20992 18880 21004
rect 17626 20964 18880 20992
rect 17626 20961 17638 20964
rect 17580 20955 17638 20961
rect 18874 20952 18880 20964
rect 18932 20952 18938 21004
rect 19245 20995 19303 21001
rect 19245 20961 19257 20995
rect 19291 20992 19303 20995
rect 19337 20995 19395 21001
rect 19337 20992 19349 20995
rect 19291 20964 19349 20992
rect 19291 20961 19303 20964
rect 19245 20955 19303 20961
rect 19337 20961 19349 20964
rect 19383 20992 19395 20995
rect 20438 20992 20444 21004
rect 19383 20964 20444 20992
rect 19383 20961 19395 20964
rect 19337 20955 19395 20961
rect 20438 20952 20444 20964
rect 20496 20952 20502 21004
rect 21008 21001 21036 21032
rect 21744 21004 21772 21032
rect 22002 21020 22008 21072
rect 22060 21060 22066 21072
rect 22557 21063 22615 21069
rect 22557 21060 22569 21063
rect 22060 21032 22569 21060
rect 22060 21020 22066 21032
rect 22557 21029 22569 21032
rect 22603 21029 22615 21063
rect 22557 21023 22615 21029
rect 20717 20995 20775 21001
rect 20717 20961 20729 20995
rect 20763 20992 20775 20995
rect 20993 20995 21051 21001
rect 20993 20992 21005 20995
rect 20763 20964 21005 20992
rect 20763 20961 20775 20964
rect 20717 20955 20775 20961
rect 20993 20961 21005 20964
rect 21039 20961 21051 20995
rect 20993 20955 21051 20961
rect 21174 20952 21180 21004
rect 21232 20992 21238 21004
rect 21269 20995 21327 21001
rect 21269 20992 21281 20995
rect 21232 20964 21281 20992
rect 21232 20952 21238 20964
rect 21269 20961 21281 20964
rect 21315 20961 21327 20995
rect 21269 20955 21327 20961
rect 21358 20952 21364 21004
rect 21416 20992 21422 21004
rect 21545 20995 21603 21001
rect 21545 20992 21557 20995
rect 21416 20964 21557 20992
rect 21416 20952 21422 20964
rect 21545 20961 21557 20964
rect 21591 20961 21603 20995
rect 21545 20955 21603 20961
rect 21726 20952 21732 21004
rect 21784 20952 21790 21004
rect 21821 20995 21879 21001
rect 21821 20961 21833 20995
rect 21867 20992 21879 20995
rect 22094 20992 22100 21004
rect 21867 20964 22100 20992
rect 21867 20961 21879 20964
rect 21821 20955 21879 20961
rect 22094 20952 22100 20964
rect 22152 20952 22158 21004
rect 22189 20995 22247 21001
rect 22189 20961 22201 20995
rect 22235 20961 22247 20995
rect 22189 20955 22247 20961
rect 9030 20884 9036 20936
rect 9088 20924 9094 20936
rect 9309 20927 9367 20933
rect 9309 20924 9321 20927
rect 9088 20896 9321 20924
rect 9088 20884 9094 20896
rect 9309 20893 9321 20896
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 13173 20927 13231 20933
rect 13173 20893 13185 20927
rect 13219 20924 13231 20927
rect 13446 20924 13452 20936
rect 13219 20896 13452 20924
rect 13219 20893 13231 20896
rect 13173 20887 13231 20893
rect 13446 20884 13452 20896
rect 13504 20884 13510 20936
rect 14090 20884 14096 20936
rect 14148 20924 14154 20936
rect 14369 20927 14427 20933
rect 14369 20924 14381 20927
rect 14148 20896 14381 20924
rect 14148 20884 14154 20896
rect 14369 20893 14381 20896
rect 14415 20893 14427 20927
rect 14369 20887 14427 20893
rect 15654 20884 15660 20936
rect 15712 20924 15718 20936
rect 15841 20927 15899 20933
rect 15841 20924 15853 20927
rect 15712 20896 15853 20924
rect 15712 20884 15718 20896
rect 15841 20893 15853 20896
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 16942 20884 16948 20936
rect 17000 20924 17006 20936
rect 17313 20927 17371 20933
rect 17313 20924 17325 20927
rect 17000 20896 17325 20924
rect 17000 20884 17006 20896
rect 17313 20893 17325 20896
rect 17359 20893 17371 20927
rect 17313 20887 17371 20893
rect 18414 20884 18420 20936
rect 18472 20924 18478 20936
rect 22204 20924 22232 20955
rect 22278 20952 22284 21004
rect 22336 20992 22342 21004
rect 22925 20995 22983 21001
rect 22925 20992 22937 20995
rect 22336 20964 22937 20992
rect 22336 20952 22342 20964
rect 22925 20961 22937 20964
rect 22971 20961 22983 20995
rect 22925 20955 22983 20961
rect 23474 20924 23480 20936
rect 18472 20896 22232 20924
rect 22296 20896 23480 20924
rect 18472 20884 18478 20896
rect 11330 20856 11336 20868
rect 8312 20828 8984 20856
rect 10612 20828 11336 20856
rect 3436 20788 3464 20816
rect 4246 20788 4252 20800
rect 3436 20760 4252 20788
rect 4246 20748 4252 20760
rect 4304 20748 4310 20800
rect 6454 20748 6460 20800
rect 6512 20788 6518 20800
rect 6730 20788 6736 20800
rect 6512 20760 6736 20788
rect 6512 20748 6518 20760
rect 6730 20748 6736 20760
rect 6788 20748 6794 20800
rect 7558 20748 7564 20800
rect 7616 20788 7622 20800
rect 8205 20791 8263 20797
rect 8205 20788 8217 20791
rect 7616 20760 8217 20788
rect 7616 20748 7622 20760
rect 8205 20757 8217 20760
rect 8251 20757 8263 20791
rect 8205 20751 8263 20757
rect 8478 20748 8484 20800
rect 8536 20788 8542 20800
rect 10612 20788 10640 20828
rect 11330 20816 11336 20828
rect 11388 20816 11394 20868
rect 14182 20856 14188 20868
rect 13280 20828 14188 20856
rect 8536 20760 10640 20788
rect 10689 20791 10747 20797
rect 8536 20748 8542 20760
rect 10689 20757 10701 20791
rect 10735 20788 10747 20791
rect 11054 20788 11060 20800
rect 10735 20760 11060 20788
rect 10735 20757 10747 20760
rect 10689 20751 10747 20757
rect 11054 20748 11060 20760
rect 11112 20748 11118 20800
rect 11348 20788 11376 20816
rect 13280 20788 13308 20828
rect 14182 20816 14188 20828
rect 14240 20816 14246 20868
rect 18506 20816 18512 20868
rect 18564 20856 18570 20868
rect 20809 20859 20867 20865
rect 20809 20856 20821 20859
rect 18564 20828 20821 20856
rect 18564 20816 18570 20828
rect 20809 20825 20821 20828
rect 20855 20856 20867 20859
rect 21174 20856 21180 20868
rect 20855 20828 21180 20856
rect 20855 20825 20867 20828
rect 20809 20819 20867 20825
rect 21174 20816 21180 20828
rect 21232 20816 21238 20868
rect 21453 20859 21511 20865
rect 21453 20825 21465 20859
rect 21499 20856 21511 20859
rect 21818 20856 21824 20868
rect 21499 20828 21824 20856
rect 21499 20825 21511 20828
rect 21453 20819 21511 20825
rect 21818 20816 21824 20828
rect 21876 20816 21882 20868
rect 21910 20816 21916 20868
rect 21968 20856 21974 20868
rect 22005 20859 22063 20865
rect 22005 20856 22017 20859
rect 21968 20828 22017 20856
rect 21968 20816 21974 20828
rect 22005 20825 22017 20828
rect 22051 20825 22063 20859
rect 22005 20819 22063 20825
rect 22094 20816 22100 20868
rect 22152 20856 22158 20868
rect 22296 20856 22324 20896
rect 23474 20884 23480 20896
rect 23532 20884 23538 20936
rect 22738 20856 22744 20868
rect 22152 20828 22324 20856
rect 22699 20828 22744 20856
rect 22152 20816 22158 20828
rect 22738 20816 22744 20828
rect 22796 20816 22802 20868
rect 11348 20760 13308 20788
rect 13354 20748 13360 20800
rect 13412 20788 13418 20800
rect 15838 20788 15844 20800
rect 13412 20760 15844 20788
rect 13412 20748 13418 20760
rect 15838 20748 15844 20760
rect 15896 20748 15902 20800
rect 16574 20748 16580 20800
rect 16632 20788 16638 20800
rect 17218 20788 17224 20800
rect 16632 20760 17224 20788
rect 16632 20748 16638 20760
rect 17218 20748 17224 20760
rect 17276 20748 17282 20800
rect 18693 20791 18751 20797
rect 18693 20757 18705 20791
rect 18739 20788 18751 20791
rect 18966 20788 18972 20800
rect 18739 20760 18972 20788
rect 18739 20757 18751 20760
rect 18693 20751 18751 20757
rect 18966 20748 18972 20760
rect 19024 20748 19030 20800
rect 23014 20788 23020 20800
rect 22975 20760 23020 20788
rect 23014 20748 23020 20760
rect 23072 20748 23078 20800
rect 1104 20698 23460 20720
rect 1104 20646 4714 20698
rect 4766 20646 4778 20698
rect 4830 20646 4842 20698
rect 4894 20646 4906 20698
rect 4958 20646 12178 20698
rect 12230 20646 12242 20698
rect 12294 20646 12306 20698
rect 12358 20646 12370 20698
rect 12422 20646 19642 20698
rect 19694 20646 19706 20698
rect 19758 20646 19770 20698
rect 19822 20646 19834 20698
rect 19886 20646 23460 20698
rect 1104 20624 23460 20646
rect 2866 20544 2872 20596
rect 2924 20584 2930 20596
rect 2961 20587 3019 20593
rect 2961 20584 2973 20587
rect 2924 20556 2973 20584
rect 2924 20544 2930 20556
rect 2961 20553 2973 20556
rect 3007 20553 3019 20587
rect 2961 20547 3019 20553
rect 1581 20383 1639 20389
rect 1581 20349 1593 20383
rect 1627 20380 1639 20383
rect 2130 20380 2136 20392
rect 1627 20352 2136 20380
rect 1627 20349 1639 20352
rect 1581 20343 1639 20349
rect 2130 20340 2136 20352
rect 2188 20380 2194 20392
rect 2866 20380 2872 20392
rect 2188 20352 2872 20380
rect 2188 20340 2194 20352
rect 2866 20340 2872 20352
rect 2924 20340 2930 20392
rect 2976 20380 3004 20547
rect 6822 20544 6828 20596
rect 6880 20584 6886 20596
rect 7009 20587 7067 20593
rect 7009 20584 7021 20587
rect 6880 20556 7021 20584
rect 6880 20544 6886 20556
rect 7009 20553 7021 20556
rect 7055 20553 7067 20587
rect 8665 20587 8723 20593
rect 8665 20584 8677 20587
rect 7009 20547 7067 20553
rect 7116 20556 8677 20584
rect 7116 20516 7144 20556
rect 8665 20553 8677 20556
rect 8711 20553 8723 20587
rect 8665 20547 8723 20553
rect 9217 20587 9275 20593
rect 9217 20553 9229 20587
rect 9263 20584 9275 20587
rect 9582 20584 9588 20596
rect 9263 20556 9588 20584
rect 9263 20553 9275 20556
rect 9217 20547 9275 20553
rect 9582 20544 9588 20556
rect 9640 20544 9646 20596
rect 10870 20584 10876 20596
rect 9692 20556 10876 20584
rect 9692 20516 9720 20556
rect 10870 20544 10876 20556
rect 10928 20544 10934 20596
rect 11330 20584 11336 20596
rect 11291 20556 11336 20584
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 12710 20544 12716 20596
rect 12768 20584 12774 20596
rect 13173 20587 13231 20593
rect 13173 20584 13185 20587
rect 12768 20556 13185 20584
rect 12768 20544 12774 20556
rect 13173 20553 13185 20556
rect 13219 20553 13231 20587
rect 13173 20547 13231 20553
rect 13630 20544 13636 20596
rect 13688 20584 13694 20596
rect 13909 20587 13967 20593
rect 13909 20584 13921 20587
rect 13688 20556 13921 20584
rect 13688 20544 13694 20556
rect 13909 20553 13921 20556
rect 13955 20553 13967 20587
rect 13909 20547 13967 20553
rect 16298 20544 16304 20596
rect 16356 20584 16362 20596
rect 16669 20587 16727 20593
rect 16669 20584 16681 20587
rect 16356 20556 16681 20584
rect 16356 20544 16362 20556
rect 16669 20553 16681 20556
rect 16715 20553 16727 20587
rect 16669 20547 16727 20553
rect 17313 20587 17371 20593
rect 17313 20553 17325 20587
rect 17359 20584 17371 20587
rect 17954 20584 17960 20596
rect 17359 20556 17960 20584
rect 17359 20553 17371 20556
rect 17313 20547 17371 20553
rect 17954 20544 17960 20556
rect 18012 20544 18018 20596
rect 18322 20544 18328 20596
rect 18380 20584 18386 20596
rect 19242 20584 19248 20596
rect 18380 20556 19248 20584
rect 18380 20544 18386 20556
rect 19242 20544 19248 20556
rect 19300 20544 19306 20596
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 19613 20587 19671 20593
rect 19613 20584 19625 20587
rect 19392 20556 19625 20584
rect 19392 20544 19398 20556
rect 19613 20553 19625 20556
rect 19659 20553 19671 20587
rect 19613 20547 19671 20553
rect 21634 20544 21640 20596
rect 21692 20584 21698 20596
rect 21729 20587 21787 20593
rect 21729 20584 21741 20587
rect 21692 20556 21741 20584
rect 21692 20544 21698 20556
rect 21729 20553 21741 20556
rect 21775 20553 21787 20587
rect 22002 20584 22008 20596
rect 21963 20556 22008 20584
rect 21729 20547 21787 20553
rect 22002 20544 22008 20556
rect 22060 20544 22066 20596
rect 4908 20488 7144 20516
rect 8864 20488 9720 20516
rect 4908 20460 4936 20488
rect 3237 20451 3295 20457
rect 3237 20417 3249 20451
rect 3283 20448 3295 20451
rect 4065 20451 4123 20457
rect 4065 20448 4077 20451
rect 3283 20420 4077 20448
rect 3283 20417 3295 20420
rect 3237 20411 3295 20417
rect 4065 20417 4077 20420
rect 4111 20448 4123 20451
rect 4430 20448 4436 20460
rect 4111 20420 4436 20448
rect 4111 20417 4123 20420
rect 4065 20411 4123 20417
rect 4430 20408 4436 20420
rect 4488 20408 4494 20460
rect 4890 20448 4896 20460
rect 4803 20420 4896 20448
rect 4890 20408 4896 20420
rect 4948 20408 4954 20460
rect 5721 20451 5779 20457
rect 5721 20417 5733 20451
rect 5767 20448 5779 20451
rect 5810 20448 5816 20460
rect 5767 20420 5816 20448
rect 5767 20417 5779 20420
rect 5721 20411 5779 20417
rect 5810 20408 5816 20420
rect 5868 20408 5874 20460
rect 6086 20408 6092 20460
rect 6144 20448 6150 20460
rect 6638 20448 6644 20460
rect 6144 20420 6644 20448
rect 6144 20408 6150 20420
rect 6638 20408 6644 20420
rect 6696 20448 6702 20460
rect 7193 20451 7251 20457
rect 7193 20448 7205 20451
rect 6696 20420 7205 20448
rect 6696 20408 6702 20420
rect 7193 20417 7205 20420
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 2976 20352 3433 20380
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3421 20343 3479 20349
rect 4154 20340 4160 20392
rect 4212 20380 4218 20392
rect 4249 20383 4307 20389
rect 4249 20380 4261 20383
rect 4212 20352 4261 20380
rect 4212 20340 4218 20352
rect 4249 20349 4261 20352
rect 4295 20349 4307 20383
rect 6914 20380 6920 20392
rect 6875 20352 6920 20380
rect 4249 20343 4307 20349
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 7460 20383 7518 20389
rect 7460 20349 7472 20383
rect 7506 20380 7518 20383
rect 7926 20380 7932 20392
rect 7506 20352 7932 20380
rect 7506 20349 7518 20352
rect 7460 20343 7518 20349
rect 7926 20340 7932 20352
rect 7984 20340 7990 20392
rect 8864 20389 8892 20488
rect 14918 20476 14924 20528
rect 14976 20516 14982 20528
rect 20717 20519 20775 20525
rect 14976 20488 16988 20516
rect 14976 20476 14982 20488
rect 10873 20451 10931 20457
rect 10873 20448 10885 20451
rect 10520 20420 10885 20448
rect 8849 20383 8907 20389
rect 8849 20349 8861 20383
rect 8895 20349 8907 20383
rect 10520 20380 10548 20420
rect 10873 20417 10885 20420
rect 10919 20417 10931 20451
rect 14461 20451 14519 20457
rect 14461 20448 14473 20451
rect 10873 20411 10931 20417
rect 13648 20420 14473 20448
rect 8849 20343 8907 20349
rect 8956 20352 10548 20380
rect 1670 20272 1676 20324
rect 1728 20312 1734 20324
rect 1848 20315 1906 20321
rect 1848 20312 1860 20315
rect 1728 20284 1860 20312
rect 1728 20272 1734 20284
rect 1848 20281 1860 20284
rect 1894 20312 1906 20315
rect 3329 20315 3387 20321
rect 3329 20312 3341 20315
rect 1894 20284 3341 20312
rect 1894 20281 1906 20284
rect 1848 20275 1906 20281
rect 3329 20281 3341 20284
rect 3375 20281 3387 20315
rect 3329 20275 3387 20281
rect 3694 20272 3700 20324
rect 3752 20312 3758 20324
rect 4985 20315 5043 20321
rect 4985 20312 4997 20315
rect 3752 20284 4997 20312
rect 3752 20272 3758 20284
rect 4985 20281 4997 20284
rect 5031 20281 5043 20315
rect 4985 20275 5043 20281
rect 5813 20315 5871 20321
rect 5813 20281 5825 20315
rect 5859 20312 5871 20315
rect 6362 20312 6368 20324
rect 5859 20284 6368 20312
rect 5859 20281 5871 20284
rect 5813 20275 5871 20281
rect 6362 20272 6368 20284
rect 6420 20272 6426 20324
rect 6472 20284 6960 20312
rect 3789 20247 3847 20253
rect 3789 20213 3801 20247
rect 3835 20244 3847 20247
rect 4062 20244 4068 20256
rect 3835 20216 4068 20244
rect 3835 20213 3847 20216
rect 3789 20207 3847 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 4157 20247 4215 20253
rect 4157 20213 4169 20247
rect 4203 20244 4215 20247
rect 4246 20244 4252 20256
rect 4203 20216 4252 20244
rect 4203 20213 4215 20216
rect 4157 20207 4215 20213
rect 4246 20204 4252 20216
rect 4304 20204 4310 20256
rect 4614 20244 4620 20256
rect 4575 20216 4620 20244
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 4706 20204 4712 20256
rect 4764 20244 4770 20256
rect 5077 20247 5135 20253
rect 5077 20244 5089 20247
rect 4764 20216 5089 20244
rect 4764 20204 4770 20216
rect 5077 20213 5089 20216
rect 5123 20213 5135 20247
rect 5077 20207 5135 20213
rect 5445 20247 5503 20253
rect 5445 20213 5457 20247
rect 5491 20244 5503 20247
rect 5718 20244 5724 20256
rect 5491 20216 5724 20244
rect 5491 20213 5503 20216
rect 5445 20207 5503 20213
rect 5718 20204 5724 20216
rect 5776 20204 5782 20256
rect 5902 20204 5908 20256
rect 5960 20244 5966 20256
rect 6273 20247 6331 20253
rect 5960 20216 6005 20244
rect 5960 20204 5966 20216
rect 6273 20213 6285 20247
rect 6319 20244 6331 20247
rect 6472 20244 6500 20284
rect 6932 20256 6960 20284
rect 8754 20272 8760 20324
rect 8812 20312 8818 20324
rect 8956 20312 8984 20352
rect 10594 20340 10600 20392
rect 10652 20380 10658 20392
rect 11514 20380 11520 20392
rect 10652 20352 11520 20380
rect 10652 20340 10658 20352
rect 11514 20340 11520 20352
rect 11572 20380 11578 20392
rect 12986 20380 12992 20392
rect 11572 20352 12992 20380
rect 11572 20340 11578 20352
rect 12986 20340 12992 20352
rect 13044 20380 13050 20392
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 13044 20352 13093 20380
rect 13044 20340 13050 20352
rect 13081 20349 13093 20352
rect 13127 20349 13139 20383
rect 13081 20343 13139 20349
rect 13262 20340 13268 20392
rect 13320 20380 13326 20392
rect 13357 20383 13415 20389
rect 13357 20380 13369 20383
rect 13320 20352 13369 20380
rect 13320 20340 13326 20352
rect 13357 20349 13369 20352
rect 13403 20349 13415 20383
rect 13357 20343 13415 20349
rect 8812 20284 8984 20312
rect 9125 20315 9183 20321
rect 8812 20272 8818 20284
rect 9125 20281 9137 20315
rect 9171 20312 9183 20315
rect 10134 20312 10140 20324
rect 9171 20284 10140 20312
rect 9171 20281 9183 20284
rect 9125 20275 9183 20281
rect 10134 20272 10140 20284
rect 10192 20272 10198 20324
rect 10226 20272 10232 20324
rect 10284 20312 10290 20324
rect 10330 20315 10388 20321
rect 10330 20312 10342 20315
rect 10284 20284 10342 20312
rect 10284 20272 10290 20284
rect 10330 20281 10342 20284
rect 10376 20281 10388 20315
rect 10330 20275 10388 20281
rect 10502 20272 10508 20324
rect 10560 20312 10566 20324
rect 10781 20315 10839 20321
rect 10781 20312 10793 20315
rect 10560 20284 10793 20312
rect 10560 20272 10566 20284
rect 10781 20281 10793 20284
rect 10827 20281 10839 20315
rect 10781 20275 10839 20281
rect 12802 20272 12808 20324
rect 12860 20321 12866 20324
rect 12860 20312 12872 20321
rect 12860 20284 12905 20312
rect 12860 20275 12872 20284
rect 12860 20272 12866 20275
rect 13446 20272 13452 20324
rect 13504 20312 13510 20324
rect 13648 20321 13676 20420
rect 14461 20417 14473 20420
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 14734 20408 14740 20460
rect 14792 20448 14798 20460
rect 14829 20451 14887 20457
rect 14829 20448 14841 20451
rect 14792 20420 14841 20448
rect 14792 20408 14798 20420
rect 14829 20417 14841 20420
rect 14875 20417 14887 20451
rect 14829 20411 14887 20417
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20448 15807 20451
rect 16206 20448 16212 20460
rect 15795 20420 16212 20448
rect 15795 20417 15807 20420
rect 15749 20411 15807 20417
rect 16206 20408 16212 20420
rect 16264 20408 16270 20460
rect 14274 20380 14280 20392
rect 14235 20352 14280 20380
rect 14274 20340 14280 20352
rect 14332 20340 14338 20392
rect 14369 20383 14427 20389
rect 14369 20349 14381 20383
rect 14415 20380 14427 20383
rect 14642 20380 14648 20392
rect 14415 20352 14648 20380
rect 14415 20349 14427 20352
rect 14369 20343 14427 20349
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 15841 20383 15899 20389
rect 15841 20380 15853 20383
rect 15252 20352 15853 20380
rect 15252 20340 15258 20352
rect 15841 20349 15853 20352
rect 15887 20380 15899 20383
rect 16577 20383 16635 20389
rect 16577 20380 16589 20383
rect 15887 20352 16589 20380
rect 15887 20349 15899 20352
rect 15841 20343 15899 20349
rect 16577 20349 16589 20352
rect 16623 20349 16635 20383
rect 16577 20343 16635 20349
rect 13633 20315 13691 20321
rect 13633 20312 13645 20315
rect 13504 20284 13645 20312
rect 13504 20272 13510 20284
rect 13633 20281 13645 20284
rect 13679 20281 13691 20315
rect 13633 20275 13691 20281
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 15105 20315 15163 20321
rect 15105 20312 15117 20315
rect 13872 20284 15117 20312
rect 13872 20272 13878 20284
rect 15105 20281 15117 20284
rect 15151 20281 15163 20315
rect 15933 20315 15991 20321
rect 15933 20312 15945 20315
rect 15105 20275 15163 20281
rect 15488 20284 15945 20312
rect 6638 20244 6644 20256
rect 6319 20216 6500 20244
rect 6599 20216 6644 20244
rect 6319 20213 6331 20216
rect 6273 20207 6331 20213
rect 6638 20204 6644 20216
rect 6696 20204 6702 20256
rect 6730 20204 6736 20256
rect 6788 20244 6794 20256
rect 6788 20216 6833 20244
rect 6788 20204 6794 20216
rect 6914 20204 6920 20256
rect 6972 20204 6978 20256
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 8573 20247 8631 20253
rect 8573 20244 8585 20247
rect 8352 20216 8585 20244
rect 8352 20204 8358 20216
rect 8573 20213 8585 20216
rect 8619 20213 8631 20247
rect 8573 20207 8631 20213
rect 9766 20204 9772 20256
rect 9824 20244 9830 20256
rect 10873 20247 10931 20253
rect 10873 20244 10885 20247
rect 9824 20216 10885 20244
rect 9824 20204 9830 20216
rect 10873 20213 10885 20216
rect 10919 20213 10931 20247
rect 10873 20207 10931 20213
rect 11701 20247 11759 20253
rect 11701 20213 11713 20247
rect 11747 20244 11759 20247
rect 12618 20244 12624 20256
rect 11747 20216 12624 20244
rect 11747 20213 11759 20216
rect 11701 20207 11759 20213
rect 12618 20204 12624 20216
rect 12676 20244 12682 20256
rect 12894 20244 12900 20256
rect 12676 20216 12900 20244
rect 12676 20204 12682 20216
rect 12894 20204 12900 20216
rect 12952 20204 12958 20256
rect 15010 20244 15016 20256
rect 14971 20216 15016 20244
rect 15010 20204 15016 20216
rect 15068 20204 15074 20256
rect 15488 20253 15516 20284
rect 15933 20281 15945 20284
rect 15979 20312 15991 20315
rect 16850 20312 16856 20324
rect 15979 20284 16856 20312
rect 15979 20281 15991 20284
rect 15933 20275 15991 20281
rect 16850 20272 16856 20284
rect 16908 20272 16914 20324
rect 16960 20312 16988 20488
rect 20717 20485 20729 20519
rect 20763 20516 20775 20519
rect 21542 20516 21548 20528
rect 20763 20488 21548 20516
rect 20763 20485 20775 20488
rect 20717 20479 20775 20485
rect 21542 20476 21548 20488
rect 21600 20476 21606 20528
rect 18874 20448 18880 20460
rect 18835 20420 18880 20448
rect 18874 20408 18880 20420
rect 18932 20408 18938 20460
rect 18966 20408 18972 20460
rect 19024 20448 19030 20460
rect 20165 20451 20223 20457
rect 20165 20448 20177 20451
rect 19024 20420 20177 20448
rect 19024 20408 19030 20420
rect 20165 20417 20177 20420
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 21284 20420 22094 20448
rect 17129 20383 17187 20389
rect 17129 20349 17141 20383
rect 17175 20380 17187 20383
rect 18693 20383 18751 20389
rect 17175 20352 18552 20380
rect 17175 20349 17187 20352
rect 17129 20343 17187 20349
rect 18322 20312 18328 20324
rect 16960 20284 18328 20312
rect 18322 20272 18328 20284
rect 18380 20272 18386 20324
rect 18426 20315 18484 20321
rect 18426 20281 18438 20315
rect 18472 20281 18484 20315
rect 18524 20312 18552 20352
rect 18693 20349 18705 20383
rect 18739 20380 18751 20383
rect 18782 20380 18788 20392
rect 18739 20352 18788 20380
rect 18739 20349 18751 20352
rect 18693 20343 18751 20349
rect 18782 20340 18788 20352
rect 18840 20340 18846 20392
rect 20898 20340 20904 20392
rect 20956 20380 20962 20392
rect 21284 20389 21312 20420
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20956 20352 21005 20380
rect 20956 20340 20962 20352
rect 20993 20349 21005 20352
rect 21039 20349 21051 20383
rect 20993 20343 21051 20349
rect 21269 20383 21327 20389
rect 21269 20349 21281 20383
rect 21315 20349 21327 20383
rect 21545 20383 21603 20389
rect 21545 20380 21557 20383
rect 21269 20343 21327 20349
rect 21376 20352 21557 20380
rect 19153 20315 19211 20321
rect 19153 20312 19165 20315
rect 18524 20284 19165 20312
rect 18426 20275 18484 20281
rect 19153 20281 19165 20284
rect 19199 20281 19211 20315
rect 19981 20315 20039 20321
rect 19981 20312 19993 20315
rect 19153 20275 19211 20281
rect 19536 20284 19993 20312
rect 15473 20247 15531 20253
rect 15473 20213 15485 20247
rect 15519 20213 15531 20247
rect 15473 20207 15531 20213
rect 16206 20204 16212 20256
rect 16264 20244 16270 20256
rect 16301 20247 16359 20253
rect 16301 20244 16313 20247
rect 16264 20216 16313 20244
rect 16264 20204 16270 20216
rect 16301 20213 16313 20216
rect 16347 20213 16359 20247
rect 16301 20207 16359 20213
rect 16390 20204 16396 20256
rect 16448 20244 16454 20256
rect 18432 20244 18460 20275
rect 19536 20256 19564 20284
rect 19981 20281 19993 20284
rect 20027 20281 20039 20315
rect 21376 20312 21404 20352
rect 21545 20349 21557 20352
rect 21591 20349 21603 20383
rect 21545 20343 21603 20349
rect 21634 20340 21640 20392
rect 21692 20380 21698 20392
rect 21821 20383 21879 20389
rect 21821 20380 21833 20383
rect 21692 20352 21833 20380
rect 21692 20340 21698 20352
rect 21821 20349 21833 20352
rect 21867 20349 21879 20383
rect 21821 20343 21879 20349
rect 22066 20312 22094 20420
rect 22186 20340 22192 20392
rect 22244 20380 22250 20392
rect 22465 20383 22523 20389
rect 22465 20380 22477 20383
rect 22244 20352 22477 20380
rect 22244 20340 22250 20352
rect 22465 20349 22477 20352
rect 22511 20349 22523 20383
rect 22465 20343 22523 20349
rect 22830 20312 22836 20324
rect 19981 20275 20039 20281
rect 20456 20284 21404 20312
rect 21468 20284 21956 20312
rect 22066 20284 22324 20312
rect 22791 20284 22836 20312
rect 18966 20244 18972 20256
rect 16448 20216 16493 20244
rect 18432 20216 18972 20244
rect 16448 20204 16454 20216
rect 18966 20204 18972 20216
rect 19024 20204 19030 20256
rect 19058 20204 19064 20256
rect 19116 20244 19122 20256
rect 19518 20244 19524 20256
rect 19116 20216 19161 20244
rect 19479 20216 19524 20244
rect 19116 20204 19122 20216
rect 19518 20204 19524 20216
rect 19576 20204 19582 20256
rect 20070 20244 20076 20256
rect 20031 20216 20076 20244
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 20254 20204 20260 20256
rect 20312 20244 20318 20256
rect 20456 20253 20484 20284
rect 20441 20247 20499 20253
rect 20441 20244 20453 20247
rect 20312 20216 20453 20244
rect 20312 20204 20318 20216
rect 20441 20213 20453 20216
rect 20487 20213 20499 20247
rect 20898 20244 20904 20256
rect 20859 20216 20904 20244
rect 20441 20207 20499 20213
rect 20898 20204 20904 20216
rect 20956 20204 20962 20256
rect 21174 20244 21180 20256
rect 21135 20216 21180 20244
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 21468 20253 21496 20284
rect 21453 20247 21511 20253
rect 21453 20213 21465 20247
rect 21499 20213 21511 20247
rect 21928 20244 21956 20284
rect 22094 20244 22100 20256
rect 21928 20216 22100 20244
rect 21453 20207 21511 20213
rect 22094 20204 22100 20216
rect 22152 20204 22158 20256
rect 22296 20253 22324 20284
rect 22830 20272 22836 20284
rect 22888 20272 22894 20324
rect 22281 20247 22339 20253
rect 22281 20213 22293 20247
rect 22327 20244 22339 20247
rect 23569 20247 23627 20253
rect 23569 20244 23581 20247
rect 22327 20216 23581 20244
rect 22327 20213 22339 20216
rect 22281 20207 22339 20213
rect 23569 20213 23581 20216
rect 23615 20213 23627 20247
rect 23569 20207 23627 20213
rect 1104 20154 23460 20176
rect 1104 20102 8446 20154
rect 8498 20102 8510 20154
rect 8562 20102 8574 20154
rect 8626 20102 8638 20154
rect 8690 20102 15910 20154
rect 15962 20102 15974 20154
rect 16026 20102 16038 20154
rect 16090 20102 16102 20154
rect 16154 20102 23460 20154
rect 1104 20080 23460 20102
rect 1581 20043 1639 20049
rect 1581 20009 1593 20043
rect 1627 20040 1639 20043
rect 1670 20040 1676 20052
rect 1627 20012 1676 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 1670 20000 1676 20012
rect 1728 20000 1734 20052
rect 3694 20040 3700 20052
rect 3655 20012 3700 20040
rect 3694 20000 3700 20012
rect 3752 20000 3758 20052
rect 3881 20043 3939 20049
rect 3881 20009 3893 20043
rect 3927 20009 3939 20043
rect 3881 20003 3939 20009
rect 4249 20043 4307 20049
rect 4249 20009 4261 20043
rect 4295 20040 4307 20043
rect 4614 20040 4620 20052
rect 4295 20012 4620 20040
rect 4295 20009 4307 20012
rect 4249 20003 4307 20009
rect 3896 19972 3924 20003
rect 4614 20000 4620 20012
rect 4672 20000 4678 20052
rect 5445 20043 5503 20049
rect 5445 20009 5457 20043
rect 5491 20040 5503 20043
rect 5626 20040 5632 20052
rect 5491 20012 5632 20040
rect 5491 20009 5503 20012
rect 5445 20003 5503 20009
rect 5626 20000 5632 20012
rect 5684 20040 5690 20052
rect 5813 20043 5871 20049
rect 5813 20040 5825 20043
rect 5684 20012 5825 20040
rect 5684 20000 5690 20012
rect 5813 20009 5825 20012
rect 5859 20009 5871 20043
rect 6362 20040 6368 20052
rect 6323 20012 6368 20040
rect 5813 20003 5871 20009
rect 6362 20000 6368 20012
rect 6420 20000 6426 20052
rect 7101 20043 7159 20049
rect 7101 20009 7113 20043
rect 7147 20040 7159 20043
rect 7834 20040 7840 20052
rect 7147 20012 7840 20040
rect 7147 20009 7159 20012
rect 7101 20003 7159 20009
rect 7834 20000 7840 20012
rect 7892 20040 7898 20052
rect 8754 20040 8760 20052
rect 7892 20012 8616 20040
rect 8715 20012 8760 20040
rect 7892 20000 7898 20012
rect 3252 19944 3924 19972
rect 2705 19907 2763 19913
rect 2705 19873 2717 19907
rect 2751 19904 2763 19907
rect 3050 19904 3056 19916
rect 2751 19876 3056 19904
rect 2751 19873 2763 19876
rect 2705 19867 2763 19873
rect 3050 19864 3056 19876
rect 3108 19864 3114 19916
rect 3252 19913 3280 19944
rect 4062 19932 4068 19984
rect 4120 19972 4126 19984
rect 4341 19975 4399 19981
rect 4341 19972 4353 19975
rect 4120 19944 4353 19972
rect 4120 19932 4126 19944
rect 4341 19941 4353 19944
rect 4387 19941 4399 19975
rect 4341 19935 4399 19941
rect 5718 19932 5724 19984
rect 5776 19972 5782 19984
rect 5905 19975 5963 19981
rect 5905 19972 5917 19975
rect 5776 19944 5917 19972
rect 5776 19932 5782 19944
rect 5905 19941 5917 19944
rect 5951 19941 5963 19975
rect 6730 19972 6736 19984
rect 5905 19935 5963 19941
rect 6196 19944 6736 19972
rect 3237 19907 3295 19913
rect 3237 19873 3249 19907
rect 3283 19873 3295 19907
rect 3510 19904 3516 19916
rect 3471 19876 3516 19904
rect 3237 19867 3295 19873
rect 3510 19864 3516 19876
rect 3568 19864 3574 19916
rect 5077 19907 5135 19913
rect 5077 19873 5089 19907
rect 5123 19904 5135 19907
rect 5166 19904 5172 19916
rect 5123 19876 5172 19904
rect 5123 19873 5135 19876
rect 5077 19867 5135 19873
rect 5166 19864 5172 19876
rect 5224 19864 5230 19916
rect 2958 19836 2964 19848
rect 2919 19808 2964 19836
rect 2958 19796 2964 19808
rect 3016 19796 3022 19848
rect 4522 19836 4528 19848
rect 4483 19808 4528 19836
rect 4522 19796 4528 19808
rect 4580 19796 4586 19848
rect 4890 19836 4896 19848
rect 4851 19808 4896 19836
rect 4890 19796 4896 19808
rect 4948 19796 4954 19848
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19805 5043 19839
rect 4985 19799 5043 19805
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19836 5779 19839
rect 6196 19836 6224 19944
rect 6730 19932 6736 19944
rect 6788 19932 6794 19984
rect 8294 19981 8300 19984
rect 8236 19975 8300 19981
rect 8236 19941 8248 19975
rect 8282 19941 8300 19975
rect 8236 19935 8300 19941
rect 8294 19932 8300 19935
rect 8352 19932 8358 19984
rect 8588 19972 8616 20012
rect 8754 20000 8760 20012
rect 8812 20000 8818 20052
rect 10502 20040 10508 20052
rect 9048 20012 10508 20040
rect 9048 19972 9076 20012
rect 10502 20000 10508 20012
rect 10560 20000 10566 20052
rect 10778 20000 10784 20052
rect 10836 20040 10842 20052
rect 11149 20043 11207 20049
rect 11149 20040 11161 20043
rect 10836 20012 11161 20040
rect 10836 20000 10842 20012
rect 11149 20009 11161 20012
rect 11195 20009 11207 20043
rect 11974 20040 11980 20052
rect 11935 20012 11980 20040
rect 11149 20003 11207 20009
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 12437 20043 12495 20049
rect 12437 20009 12449 20043
rect 12483 20040 12495 20043
rect 12894 20040 12900 20052
rect 12483 20012 12756 20040
rect 12855 20012 12900 20040
rect 12483 20009 12495 20012
rect 12437 20003 12495 20009
rect 8588 19944 9076 19972
rect 9858 19932 9864 19984
rect 9916 19981 9922 19984
rect 9916 19975 9980 19981
rect 9916 19941 9934 19975
rect 9968 19941 9980 19975
rect 9916 19935 9980 19941
rect 9916 19932 9922 19935
rect 11054 19932 11060 19984
rect 11112 19972 11118 19984
rect 12728 19972 12756 20012
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 13265 20043 13323 20049
rect 13265 20009 13277 20043
rect 13311 20040 13323 20043
rect 13725 20043 13783 20049
rect 13725 20040 13737 20043
rect 13311 20012 13737 20040
rect 13311 20009 13323 20012
rect 13265 20003 13323 20009
rect 13725 20009 13737 20012
rect 13771 20009 13783 20043
rect 13725 20003 13783 20009
rect 14366 20000 14372 20052
rect 14424 20040 14430 20052
rect 14424 20012 14872 20040
rect 14424 20000 14430 20012
rect 13814 19972 13820 19984
rect 11112 19944 11744 19972
rect 12728 19944 13820 19972
rect 11112 19932 11118 19944
rect 6549 19907 6607 19913
rect 6549 19904 6561 19907
rect 5767 19808 6224 19836
rect 6288 19876 6561 19904
rect 5767 19805 5779 19808
rect 5721 19799 5779 19805
rect 3421 19771 3479 19777
rect 3421 19737 3433 19771
rect 3467 19768 3479 19771
rect 4706 19768 4712 19780
rect 3467 19740 4712 19768
rect 3467 19737 3479 19740
rect 3421 19731 3479 19737
rect 4706 19728 4712 19740
rect 4764 19728 4770 19780
rect 5000 19768 5028 19799
rect 5074 19768 5080 19780
rect 5000 19740 5080 19768
rect 5074 19728 5080 19740
rect 5132 19728 5138 19780
rect 6288 19777 6316 19876
rect 6549 19873 6561 19876
rect 6595 19873 6607 19907
rect 6549 19867 6607 19873
rect 6822 19864 6828 19916
rect 6880 19904 6886 19916
rect 8938 19904 8944 19916
rect 6880 19876 8944 19904
rect 6880 19864 6886 19876
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 9306 19864 9312 19916
rect 9364 19904 9370 19916
rect 11517 19907 11575 19913
rect 11517 19904 11529 19907
rect 9364 19876 11529 19904
rect 9364 19864 9370 19876
rect 11517 19873 11529 19876
rect 11563 19873 11575 19907
rect 11517 19867 11575 19873
rect 8481 19839 8539 19845
rect 8481 19805 8493 19839
rect 8527 19836 8539 19839
rect 8754 19836 8760 19848
rect 8527 19808 8760 19836
rect 8527 19805 8539 19808
rect 8481 19799 8539 19805
rect 8754 19796 8760 19808
rect 8812 19836 8818 19848
rect 9030 19836 9036 19848
rect 8812 19808 9036 19836
rect 8812 19796 8818 19808
rect 9030 19796 9036 19808
rect 9088 19836 9094 19848
rect 9677 19839 9735 19845
rect 9677 19836 9689 19839
rect 9088 19808 9689 19836
rect 9088 19796 9094 19808
rect 9677 19805 9689 19808
rect 9723 19805 9735 19839
rect 9677 19799 9735 19805
rect 6273 19771 6331 19777
rect 6273 19737 6285 19771
rect 6319 19737 6331 19771
rect 6273 19731 6331 19737
rect 3142 19700 3148 19712
rect 3103 19672 3148 19700
rect 3142 19660 3148 19672
rect 3200 19660 3206 19712
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 6733 19703 6791 19709
rect 6733 19700 6745 19703
rect 5592 19672 6745 19700
rect 5592 19660 5598 19672
rect 6733 19669 6745 19672
rect 6779 19700 6791 19703
rect 8570 19700 8576 19712
rect 6779 19672 8576 19700
rect 6779 19669 6791 19672
rect 6733 19663 6791 19669
rect 8570 19660 8576 19672
rect 8628 19660 8634 19712
rect 9217 19703 9275 19709
rect 9217 19669 9229 19703
rect 9263 19700 9275 19703
rect 9398 19700 9404 19712
rect 9263 19672 9404 19700
rect 9263 19669 9275 19672
rect 9217 19663 9275 19669
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 9692 19700 9720 19799
rect 10962 19796 10968 19848
rect 11020 19836 11026 19848
rect 11716 19845 11744 19944
rect 13814 19932 13820 19944
rect 13872 19932 13878 19984
rect 13906 19932 13912 19984
rect 13964 19932 13970 19984
rect 14550 19932 14556 19984
rect 14608 19972 14614 19984
rect 14737 19975 14795 19981
rect 14737 19972 14749 19975
rect 14608 19944 14749 19972
rect 14608 19932 14614 19944
rect 14737 19941 14749 19944
rect 14783 19941 14795 19975
rect 14844 19972 14872 20012
rect 15010 20000 15016 20052
rect 15068 20040 15074 20052
rect 15289 20043 15347 20049
rect 15289 20040 15301 20043
rect 15068 20012 15301 20040
rect 15068 20000 15074 20012
rect 15289 20009 15301 20012
rect 15335 20009 15347 20043
rect 15289 20003 15347 20009
rect 15933 20043 15991 20049
rect 15933 20009 15945 20043
rect 15979 20009 15991 20043
rect 16390 20040 16396 20052
rect 16351 20012 16396 20040
rect 15933 20003 15991 20009
rect 15565 19975 15623 19981
rect 15565 19972 15577 19975
rect 14844 19944 15577 19972
rect 14737 19935 14795 19941
rect 15565 19941 15577 19944
rect 15611 19941 15623 19975
rect 15948 19972 15976 20003
rect 16390 20000 16396 20012
rect 16448 20000 16454 20052
rect 16761 20043 16819 20049
rect 16761 20009 16773 20043
rect 16807 20040 16819 20043
rect 19058 20040 19064 20052
rect 16807 20012 19064 20040
rect 16807 20009 16819 20012
rect 16761 20003 16819 20009
rect 19058 20000 19064 20012
rect 19116 20000 19122 20052
rect 19242 20000 19248 20052
rect 19300 20040 19306 20052
rect 21450 20040 21456 20052
rect 19300 20012 21456 20040
rect 19300 20000 19306 20012
rect 21450 20000 21456 20012
rect 21508 20000 21514 20052
rect 22649 20043 22707 20049
rect 22649 20009 22661 20043
rect 22695 20009 22707 20043
rect 22649 20003 22707 20009
rect 16301 19975 16359 19981
rect 16301 19972 16313 19975
rect 15948 19944 16313 19972
rect 15565 19935 15623 19941
rect 16301 19941 16313 19944
rect 16347 19941 16359 19975
rect 16301 19935 16359 19941
rect 16482 19932 16488 19984
rect 16540 19972 16546 19984
rect 17313 19975 17371 19981
rect 17313 19972 17325 19975
rect 16540 19944 17325 19972
rect 16540 19932 16546 19944
rect 17313 19941 17325 19944
rect 17359 19941 17371 19975
rect 17313 19935 17371 19941
rect 17954 19932 17960 19984
rect 18012 19972 18018 19984
rect 18702 19975 18760 19981
rect 18702 19972 18714 19975
rect 18012 19944 18714 19972
rect 18012 19932 18018 19944
rect 18702 19941 18714 19944
rect 18748 19941 18760 19975
rect 20070 19972 20076 19984
rect 18702 19935 18760 19941
rect 18800 19944 20076 19972
rect 12253 19907 12311 19913
rect 12253 19873 12265 19907
rect 12299 19904 12311 19907
rect 13170 19904 13176 19916
rect 12299 19876 13176 19904
rect 12299 19873 12311 19876
rect 12253 19867 12311 19873
rect 13170 19864 13176 19876
rect 13228 19864 13234 19916
rect 13924 19904 13952 19932
rect 14826 19904 14832 19916
rect 13556 19876 13952 19904
rect 14787 19876 14832 19904
rect 11609 19839 11667 19845
rect 11609 19836 11621 19839
rect 11020 19808 11621 19836
rect 11020 19796 11026 19808
rect 11609 19805 11621 19808
rect 11655 19805 11667 19839
rect 11609 19799 11667 19805
rect 11701 19839 11759 19845
rect 11701 19805 11713 19839
rect 11747 19805 11759 19839
rect 11701 19799 11759 19805
rect 12713 19839 12771 19845
rect 12713 19805 12725 19839
rect 12759 19805 12771 19839
rect 12713 19799 12771 19805
rect 12728 19768 12756 19799
rect 12802 19796 12808 19848
rect 12860 19836 12866 19848
rect 13078 19836 13084 19848
rect 12860 19808 13084 19836
rect 12860 19796 12866 19808
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 13556 19845 13584 19876
rect 14826 19864 14832 19876
rect 14884 19864 14890 19916
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 15749 19907 15807 19913
rect 15749 19873 15761 19907
rect 15795 19904 15807 19907
rect 16206 19904 16212 19916
rect 15795 19876 16212 19904
rect 15795 19873 15807 19876
rect 15749 19867 15807 19873
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 13633 19839 13691 19845
rect 13633 19805 13645 19839
rect 13679 19836 13691 19839
rect 13906 19836 13912 19848
rect 13679 19808 13912 19836
rect 13679 19805 13691 19808
rect 13633 19799 13691 19805
rect 13906 19796 13912 19808
rect 13964 19796 13970 19848
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19836 14703 19839
rect 14734 19836 14740 19848
rect 14691 19808 14740 19836
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 12894 19768 12900 19780
rect 12728 19740 12900 19768
rect 12894 19728 12900 19740
rect 12952 19768 12958 19780
rect 13446 19768 13452 19780
rect 12952 19740 13452 19768
rect 12952 19728 12958 19740
rect 13446 19728 13452 19740
rect 13504 19728 13510 19780
rect 14093 19771 14151 19777
rect 14093 19737 14105 19771
rect 14139 19768 14151 19771
rect 15488 19768 15516 19867
rect 16206 19864 16212 19876
rect 16264 19864 16270 19916
rect 16574 19904 16580 19916
rect 16316 19876 16580 19904
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19836 16175 19839
rect 16316 19836 16344 19876
rect 16574 19864 16580 19876
rect 16632 19864 16638 19916
rect 16850 19904 16856 19916
rect 16811 19876 16856 19904
rect 16850 19864 16856 19876
rect 16908 19864 16914 19916
rect 17402 19864 17408 19916
rect 17460 19904 17466 19916
rect 18800 19904 18828 19944
rect 20070 19932 20076 19944
rect 20128 19932 20134 19984
rect 22664 19972 22692 20003
rect 22925 19975 22983 19981
rect 22925 19972 22937 19975
rect 22664 19944 22937 19972
rect 22925 19941 22937 19944
rect 22971 19941 22983 19975
rect 22925 19935 22983 19941
rect 19978 19904 19984 19916
rect 17460 19876 18828 19904
rect 19939 19876 19984 19904
rect 17460 19864 17466 19876
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 20622 19864 20628 19916
rect 20680 19904 20686 19916
rect 20717 19907 20775 19913
rect 20717 19904 20729 19907
rect 20680 19876 20729 19904
rect 20680 19864 20686 19876
rect 20717 19873 20729 19876
rect 20763 19873 20775 19907
rect 21082 19904 21088 19916
rect 20717 19867 20775 19873
rect 20824 19876 21088 19904
rect 18966 19836 18972 19848
rect 16163 19808 16344 19836
rect 18927 19808 18972 19836
rect 16163 19805 16175 19808
rect 16117 19799 16175 19805
rect 18966 19796 18972 19808
rect 19024 19796 19030 19848
rect 19797 19839 19855 19845
rect 19797 19805 19809 19839
rect 19843 19805 19855 19839
rect 19797 19799 19855 19805
rect 19889 19839 19947 19845
rect 19889 19805 19901 19839
rect 19935 19836 19947 19839
rect 20070 19836 20076 19848
rect 19935 19808 20076 19836
rect 19935 19805 19947 19808
rect 19889 19799 19947 19805
rect 14139 19740 15516 19768
rect 14139 19737 14151 19740
rect 14093 19731 14151 19737
rect 15562 19728 15568 19780
rect 15620 19768 15626 19780
rect 17129 19771 17187 19777
rect 17129 19768 17141 19771
rect 15620 19740 17141 19768
rect 15620 19728 15626 19740
rect 17129 19737 17141 19740
rect 17175 19737 17187 19771
rect 19812 19768 19840 19799
rect 20070 19796 20076 19808
rect 20128 19796 20134 19848
rect 20714 19768 20720 19780
rect 19812 19740 20720 19768
rect 17129 19731 17187 19737
rect 20714 19728 20720 19740
rect 20772 19728 20778 19780
rect 20824 19768 20852 19876
rect 21082 19864 21088 19876
rect 21140 19864 21146 19916
rect 21260 19907 21318 19913
rect 21260 19873 21272 19907
rect 21306 19904 21318 19907
rect 22370 19904 22376 19916
rect 21306 19876 22376 19904
rect 21306 19873 21318 19876
rect 21260 19867 21318 19873
rect 22370 19864 22376 19876
rect 22428 19864 22434 19916
rect 22465 19907 22523 19913
rect 22465 19873 22477 19907
rect 22511 19904 22523 19907
rect 23198 19904 23204 19916
rect 22511 19876 23204 19904
rect 22511 19873 22523 19876
rect 22465 19867 22523 19873
rect 23198 19864 23204 19876
rect 23256 19864 23262 19916
rect 20990 19836 20996 19848
rect 20951 19808 20996 19836
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 20901 19771 20959 19777
rect 20901 19768 20913 19771
rect 20824 19740 20913 19768
rect 20901 19737 20913 19740
rect 20947 19737 20959 19771
rect 23106 19768 23112 19780
rect 23067 19740 23112 19768
rect 20901 19731 20959 19737
rect 23106 19728 23112 19740
rect 23164 19728 23170 19780
rect 10594 19700 10600 19712
rect 9692 19672 10600 19700
rect 10594 19660 10600 19672
rect 10652 19660 10658 19712
rect 11054 19700 11060 19712
rect 11015 19672 11060 19700
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 11146 19660 11152 19712
rect 11204 19700 11210 19712
rect 14458 19700 14464 19712
rect 11204 19672 14464 19700
rect 11204 19660 11210 19672
rect 14458 19660 14464 19672
rect 14516 19700 14522 19712
rect 14918 19700 14924 19712
rect 14516 19672 14924 19700
rect 14516 19660 14522 19672
rect 14918 19660 14924 19672
rect 14976 19660 14982 19712
rect 15194 19700 15200 19712
rect 15155 19672 15200 19700
rect 15194 19660 15200 19672
rect 15252 19660 15258 19712
rect 17034 19700 17040 19712
rect 16995 19672 17040 19700
rect 17034 19660 17040 19672
rect 17092 19660 17098 19712
rect 17586 19700 17592 19712
rect 17547 19672 17592 19700
rect 17586 19660 17592 19672
rect 17644 19660 17650 19712
rect 20162 19660 20168 19712
rect 20220 19700 20226 19712
rect 20349 19703 20407 19709
rect 20349 19700 20361 19703
rect 20220 19672 20361 19700
rect 20220 19660 20226 19672
rect 20349 19669 20361 19672
rect 20395 19669 20407 19703
rect 20622 19700 20628 19712
rect 20583 19672 20628 19700
rect 20349 19663 20407 19669
rect 20622 19660 20628 19672
rect 20680 19660 20686 19712
rect 22373 19703 22431 19709
rect 22373 19669 22385 19703
rect 22419 19700 22431 19703
rect 22554 19700 22560 19712
rect 22419 19672 22560 19700
rect 22419 19669 22431 19672
rect 22373 19663 22431 19669
rect 22554 19660 22560 19672
rect 22612 19660 22618 19712
rect 1104 19610 23460 19632
rect 1104 19558 4714 19610
rect 4766 19558 4778 19610
rect 4830 19558 4842 19610
rect 4894 19558 4906 19610
rect 4958 19558 12178 19610
rect 12230 19558 12242 19610
rect 12294 19558 12306 19610
rect 12358 19558 12370 19610
rect 12422 19558 19642 19610
rect 19694 19558 19706 19610
rect 19758 19558 19770 19610
rect 19822 19558 19834 19610
rect 19886 19558 23460 19610
rect 1104 19536 23460 19558
rect 3510 19456 3516 19508
rect 3568 19496 3574 19508
rect 3973 19499 4031 19505
rect 3973 19496 3985 19499
rect 3568 19468 3985 19496
rect 3568 19456 3574 19468
rect 3973 19465 3985 19468
rect 4019 19465 4031 19499
rect 3973 19459 4031 19465
rect 5813 19499 5871 19505
rect 5813 19465 5825 19499
rect 5859 19496 5871 19499
rect 5902 19496 5908 19508
rect 5859 19468 5908 19496
rect 5859 19465 5871 19468
rect 5813 19459 5871 19465
rect 5902 19456 5908 19468
rect 5960 19456 5966 19508
rect 6012 19468 8892 19496
rect 3142 19388 3148 19440
rect 3200 19428 3206 19440
rect 4338 19428 4344 19440
rect 3200 19400 4344 19428
rect 3200 19388 3206 19400
rect 4338 19388 4344 19400
rect 4396 19428 4402 19440
rect 6012 19428 6040 19468
rect 4396 19400 6040 19428
rect 8864 19428 8892 19468
rect 9122 19456 9128 19508
rect 9180 19496 9186 19508
rect 9309 19499 9367 19505
rect 9309 19496 9321 19499
rect 9180 19468 9321 19496
rect 9180 19456 9186 19468
rect 9309 19465 9321 19468
rect 9355 19465 9367 19499
rect 11514 19496 11520 19508
rect 11475 19468 11520 19496
rect 9309 19459 9367 19465
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 13078 19496 13084 19508
rect 13039 19468 13084 19496
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 19797 19499 19855 19505
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 20070 19496 20076 19508
rect 19843 19468 20076 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 20070 19456 20076 19468
rect 20128 19456 20134 19508
rect 21545 19499 21603 19505
rect 21545 19465 21557 19499
rect 21591 19496 21603 19499
rect 22278 19496 22284 19508
rect 21591 19468 22284 19496
rect 21591 19465 21603 19468
rect 21545 19459 21603 19465
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 11146 19428 11152 19440
rect 8864 19400 11152 19428
rect 4396 19388 4402 19400
rect 11146 19388 11152 19400
rect 11204 19388 11210 19440
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 4430 19360 4436 19372
rect 3375 19332 4436 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 4522 19320 4528 19372
rect 4580 19360 4586 19372
rect 4617 19363 4675 19369
rect 4617 19360 4629 19363
rect 4580 19332 4629 19360
rect 4580 19320 4586 19332
rect 4617 19329 4629 19332
rect 4663 19360 4675 19363
rect 5442 19360 5448 19372
rect 4663 19332 5448 19360
rect 4663 19329 4675 19332
rect 4617 19323 4675 19329
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 6454 19320 6460 19372
rect 6512 19360 6518 19372
rect 6549 19363 6607 19369
rect 6549 19360 6561 19363
rect 6512 19332 6561 19360
rect 6512 19320 6518 19332
rect 6549 19329 6561 19332
rect 6595 19329 6607 19363
rect 6549 19323 6607 19329
rect 6733 19363 6791 19369
rect 6733 19329 6745 19363
rect 6779 19360 6791 19363
rect 6914 19360 6920 19372
rect 6779 19332 6920 19360
rect 6779 19329 6791 19332
rect 6733 19323 6791 19329
rect 6914 19320 6920 19332
rect 6972 19320 6978 19372
rect 7932 19363 7990 19369
rect 7932 19360 7944 19363
rect 7576 19332 7944 19360
rect 1673 19295 1731 19301
rect 1673 19261 1685 19295
rect 1719 19292 1731 19295
rect 5626 19292 5632 19304
rect 1719 19264 2176 19292
rect 5587 19264 5632 19292
rect 1719 19261 1731 19264
rect 1673 19255 1731 19261
rect 2148 19236 2176 19264
rect 5626 19252 5632 19264
rect 5684 19252 5690 19304
rect 5718 19252 5724 19304
rect 5776 19292 5782 19304
rect 5905 19295 5963 19301
rect 5905 19292 5917 19295
rect 5776 19264 5917 19292
rect 5776 19252 5782 19264
rect 5905 19261 5917 19264
rect 5951 19261 5963 19295
rect 5905 19255 5963 19261
rect 6638 19252 6644 19304
rect 6696 19292 6702 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6696 19264 6837 19292
rect 6696 19252 6702 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 6825 19255 6883 19261
rect 7374 19252 7380 19304
rect 7432 19292 7438 19304
rect 7469 19295 7527 19301
rect 7469 19292 7481 19295
rect 7432 19264 7481 19292
rect 7432 19252 7438 19264
rect 7469 19261 7481 19264
rect 7515 19261 7527 19295
rect 7469 19255 7527 19261
rect 1946 19233 1952 19236
rect 1940 19224 1952 19233
rect 1907 19196 1952 19224
rect 1940 19187 1952 19196
rect 1946 19184 1952 19187
rect 2004 19184 2010 19236
rect 2130 19184 2136 19236
rect 2188 19184 2194 19236
rect 2222 19184 2228 19236
rect 2280 19224 2286 19236
rect 3513 19227 3571 19233
rect 3513 19224 3525 19227
rect 2280 19196 3525 19224
rect 2280 19184 2286 19196
rect 3513 19193 3525 19196
rect 3559 19193 3571 19227
rect 4433 19227 4491 19233
rect 4433 19224 4445 19227
rect 3513 19187 3571 19193
rect 3896 19196 4445 19224
rect 3050 19156 3056 19168
rect 3011 19128 3056 19156
rect 3050 19116 3056 19128
rect 3108 19116 3114 19168
rect 3326 19116 3332 19168
rect 3384 19156 3390 19168
rect 3896 19165 3924 19196
rect 4433 19193 4445 19196
rect 4479 19193 4491 19227
rect 4433 19187 4491 19193
rect 5169 19227 5227 19233
rect 5169 19193 5181 19227
rect 5215 19224 5227 19227
rect 5810 19224 5816 19236
rect 5215 19196 5816 19224
rect 5215 19193 5227 19196
rect 5169 19187 5227 19193
rect 5810 19184 5816 19196
rect 5868 19184 5874 19236
rect 7576 19224 7604 19332
rect 7932 19329 7944 19332
rect 7978 19360 7990 19363
rect 8110 19360 8116 19372
rect 7978 19332 8116 19360
rect 7978 19329 7990 19332
rect 7932 19323 7990 19329
rect 8110 19320 8116 19332
rect 8168 19320 8174 19372
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 8628 19332 9812 19360
rect 8628 19320 8634 19332
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 8205 19295 8263 19301
rect 8205 19292 8217 19295
rect 7800 19264 8217 19292
rect 7800 19252 7806 19264
rect 8205 19261 8217 19264
rect 8251 19261 8263 19295
rect 9784 19292 9812 19332
rect 9858 19320 9864 19372
rect 9916 19360 9922 19372
rect 10226 19360 10232 19372
rect 9916 19332 10232 19360
rect 9916 19320 9922 19332
rect 10226 19320 10232 19332
rect 10284 19320 10290 19372
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 10597 19363 10655 19369
rect 10597 19360 10609 19363
rect 10468 19332 10609 19360
rect 10468 19320 10474 19332
rect 10597 19329 10609 19332
rect 10643 19329 10655 19363
rect 10597 19323 10655 19329
rect 10686 19320 10692 19372
rect 10744 19320 10750 19372
rect 10704 19292 10732 19320
rect 11330 19292 11336 19304
rect 9784 19264 10732 19292
rect 11291 19264 11336 19292
rect 8205 19255 8263 19261
rect 11330 19252 11336 19264
rect 11388 19252 11394 19304
rect 11532 19292 11560 19456
rect 13740 19400 15424 19428
rect 13740 19372 13768 19400
rect 12894 19320 12900 19372
rect 12952 19360 12958 19372
rect 13265 19363 13323 19369
rect 13265 19360 13277 19363
rect 12952 19332 13277 19360
rect 12952 19320 12958 19332
rect 13265 19329 13277 19332
rect 13311 19360 13323 19363
rect 13722 19360 13728 19372
rect 13311 19332 13728 19360
rect 13311 19329 13323 19332
rect 13265 19323 13323 19329
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 13998 19320 14004 19372
rect 14056 19360 14062 19372
rect 15396 19369 15424 19400
rect 20916 19400 22876 19428
rect 14093 19363 14151 19369
rect 14093 19360 14105 19363
rect 14056 19332 14105 19360
rect 14056 19320 14062 19332
rect 14093 19329 14105 19332
rect 14139 19329 14151 19363
rect 14093 19323 14151 19329
rect 15381 19363 15439 19369
rect 15381 19329 15393 19363
rect 15427 19360 15439 19363
rect 16209 19363 16267 19369
rect 16209 19360 16221 19363
rect 15427 19332 16221 19360
rect 15427 19329 15439 19332
rect 15381 19323 15439 19329
rect 16209 19329 16221 19332
rect 16255 19329 16267 19363
rect 16209 19323 16267 19329
rect 19245 19363 19303 19369
rect 19245 19329 19257 19363
rect 19291 19360 19303 19363
rect 19291 19332 20024 19360
rect 19291 19329 19303 19332
rect 19245 19323 19303 19329
rect 11701 19295 11759 19301
rect 11701 19292 11713 19295
rect 11532 19264 11713 19292
rect 11701 19261 11713 19264
rect 11747 19292 11759 19295
rect 11790 19292 11796 19304
rect 11747 19264 11796 19292
rect 11747 19261 11759 19264
rect 11701 19255 11759 19261
rect 11790 19252 11796 19264
rect 11848 19252 11854 19304
rect 14369 19295 14427 19301
rect 14369 19261 14381 19295
rect 14415 19292 14427 19295
rect 14415 19264 15700 19292
rect 14415 19261 14427 19264
rect 14369 19255 14427 19261
rect 6104 19196 7604 19224
rect 3421 19159 3479 19165
rect 3421 19156 3433 19159
rect 3384 19128 3433 19156
rect 3384 19116 3390 19128
rect 3421 19125 3433 19128
rect 3467 19125 3479 19159
rect 3421 19119 3479 19125
rect 3881 19159 3939 19165
rect 3881 19125 3893 19159
rect 3927 19125 3939 19159
rect 4338 19156 4344 19168
rect 4299 19128 4344 19156
rect 3881 19119 3939 19125
rect 4338 19116 4344 19128
rect 4396 19116 4402 19168
rect 4798 19156 4804 19168
rect 4759 19128 4804 19156
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 6104 19165 6132 19196
rect 9582 19184 9588 19236
rect 9640 19224 9646 19236
rect 10045 19227 10103 19233
rect 10045 19224 10057 19227
rect 9640 19196 10057 19224
rect 9640 19184 9646 19196
rect 10045 19193 10057 19196
rect 10091 19224 10103 19227
rect 11146 19224 11152 19236
rect 10091 19196 11152 19224
rect 10091 19193 10103 19196
rect 10045 19187 10103 19193
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 11968 19227 12026 19233
rect 11968 19193 11980 19227
rect 12014 19224 12026 19227
rect 13262 19224 13268 19236
rect 12014 19196 13268 19224
rect 12014 19193 12026 19196
rect 11968 19187 12026 19193
rect 13262 19184 13268 19196
rect 13320 19224 13326 19236
rect 13541 19227 13599 19233
rect 13541 19224 13553 19227
rect 13320 19196 13553 19224
rect 13320 19184 13326 19196
rect 13541 19193 13553 19196
rect 13587 19193 13599 19227
rect 13541 19187 13599 19193
rect 14277 19227 14335 19233
rect 14277 19193 14289 19227
rect 14323 19224 14335 19227
rect 14323 19196 14872 19224
rect 14323 19193 14335 19196
rect 14277 19187 14335 19193
rect 6089 19159 6147 19165
rect 5316 19128 5361 19156
rect 5316 19116 5322 19128
rect 6089 19125 6101 19159
rect 6135 19125 6147 19159
rect 7190 19156 7196 19168
rect 7151 19128 7196 19156
rect 6089 19119 6147 19125
rect 7190 19116 7196 19128
rect 7248 19156 7254 19168
rect 7466 19156 7472 19168
rect 7248 19128 7472 19156
rect 7248 19116 7254 19128
rect 7466 19116 7472 19128
rect 7524 19116 7530 19168
rect 7935 19159 7993 19165
rect 7935 19125 7947 19159
rect 7981 19156 7993 19159
rect 9306 19156 9312 19168
rect 7981 19128 9312 19156
rect 7981 19125 7993 19128
rect 7935 19119 7993 19125
rect 9306 19116 9312 19128
rect 9364 19156 9370 19168
rect 9493 19159 9551 19165
rect 9493 19156 9505 19159
rect 9364 19128 9505 19156
rect 9364 19116 9370 19128
rect 9493 19125 9505 19128
rect 9539 19125 9551 19159
rect 9674 19156 9680 19168
rect 9635 19128 9680 19156
rect 9493 19119 9551 19125
rect 9674 19116 9680 19128
rect 9732 19116 9738 19168
rect 10134 19156 10140 19168
rect 10095 19128 10140 19156
rect 10134 19116 10140 19128
rect 10192 19116 10198 19168
rect 10778 19156 10784 19168
rect 10739 19128 10784 19156
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 11238 19156 11244 19168
rect 10928 19128 10973 19156
rect 11199 19128 11244 19156
rect 10928 19116 10934 19128
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 12158 19116 12164 19168
rect 12216 19156 12222 19168
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 12216 19128 13461 19156
rect 12216 19116 12222 19128
rect 13449 19125 13461 19128
rect 13495 19125 13507 19159
rect 13906 19156 13912 19168
rect 13867 19128 13912 19156
rect 13449 19119 13507 19125
rect 13906 19116 13912 19128
rect 13964 19116 13970 19168
rect 14642 19116 14648 19168
rect 14700 19156 14706 19168
rect 14844 19165 14872 19196
rect 14737 19159 14795 19165
rect 14737 19156 14749 19159
rect 14700 19128 14749 19156
rect 14700 19116 14706 19128
rect 14737 19125 14749 19128
rect 14783 19125 14795 19159
rect 14737 19119 14795 19125
rect 14829 19159 14887 19165
rect 14829 19125 14841 19159
rect 14875 19125 14887 19159
rect 15194 19156 15200 19168
rect 15155 19128 15200 19156
rect 14829 19119 14887 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 15286 19116 15292 19168
rect 15344 19156 15350 19168
rect 15672 19165 15700 19264
rect 17586 19252 17592 19304
rect 17644 19292 17650 19304
rect 18058 19295 18116 19301
rect 18058 19292 18070 19295
rect 17644 19264 18070 19292
rect 17644 19252 17650 19264
rect 18058 19261 18070 19264
rect 18104 19261 18116 19295
rect 18058 19255 18116 19261
rect 18325 19295 18383 19301
rect 18325 19261 18337 19295
rect 18371 19292 18383 19295
rect 18966 19292 18972 19304
rect 18371 19264 18972 19292
rect 18371 19261 18383 19264
rect 18325 19255 18383 19261
rect 18966 19252 18972 19264
rect 19024 19292 19030 19304
rect 19150 19292 19156 19304
rect 19024 19264 19156 19292
rect 19024 19252 19030 19264
rect 19150 19252 19156 19264
rect 19208 19292 19214 19304
rect 19889 19295 19947 19301
rect 19889 19292 19901 19295
rect 19208 19264 19901 19292
rect 19208 19252 19214 19264
rect 19889 19261 19901 19264
rect 19935 19261 19947 19295
rect 19996 19292 20024 19332
rect 20530 19292 20536 19304
rect 19996 19264 20536 19292
rect 19889 19255 19947 19261
rect 20530 19252 20536 19264
rect 20588 19292 20594 19304
rect 20916 19292 20944 19400
rect 22848 19372 22876 19400
rect 21634 19320 21640 19372
rect 21692 19360 21698 19372
rect 22005 19363 22063 19369
rect 22005 19360 22017 19363
rect 21692 19332 22017 19360
rect 21692 19320 21698 19332
rect 22005 19329 22017 19332
rect 22051 19329 22063 19363
rect 22830 19360 22836 19372
rect 22791 19332 22836 19360
rect 22005 19323 22063 19329
rect 22830 19320 22836 19332
rect 22888 19320 22894 19372
rect 23566 19360 23572 19372
rect 23527 19332 23572 19360
rect 23566 19320 23572 19332
rect 23624 19320 23630 19372
rect 20588 19264 20944 19292
rect 21361 19295 21419 19301
rect 20588 19252 20594 19264
rect 21361 19261 21373 19295
rect 21407 19292 21419 19295
rect 21726 19292 21732 19304
rect 21407 19264 21732 19292
rect 21407 19261 21419 19264
rect 21361 19255 21419 19261
rect 21726 19252 21732 19264
rect 21784 19252 21790 19304
rect 21821 19295 21879 19301
rect 21821 19261 21833 19295
rect 21867 19292 21879 19295
rect 21910 19292 21916 19304
rect 21867 19264 21916 19292
rect 21867 19261 21879 19264
rect 21821 19255 21879 19261
rect 21910 19252 21916 19264
rect 21968 19252 21974 19304
rect 22370 19252 22376 19304
rect 22428 19292 22434 19304
rect 22557 19295 22615 19301
rect 22557 19292 22569 19295
rect 22428 19264 22569 19292
rect 22428 19252 22434 19264
rect 22557 19261 22569 19264
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 20156 19227 20214 19233
rect 20156 19193 20168 19227
rect 20202 19224 20214 19227
rect 20346 19224 20352 19236
rect 20202 19196 20352 19224
rect 20202 19193 20214 19196
rect 20156 19187 20214 19193
rect 20346 19184 20352 19196
rect 20404 19184 20410 19236
rect 21174 19184 21180 19236
rect 21232 19224 21238 19236
rect 21637 19227 21695 19233
rect 21637 19224 21649 19227
rect 21232 19196 21649 19224
rect 21232 19184 21238 19196
rect 21637 19193 21649 19196
rect 21683 19193 21695 19227
rect 22649 19227 22707 19233
rect 22649 19224 22661 19227
rect 21637 19187 21695 19193
rect 21744 19196 22661 19224
rect 15657 19159 15715 19165
rect 15344 19128 15389 19156
rect 15344 19116 15350 19128
rect 15657 19125 15669 19159
rect 15703 19125 15715 19159
rect 15657 19119 15715 19125
rect 15746 19116 15752 19168
rect 15804 19156 15810 19168
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 15804 19128 16037 19156
rect 15804 19116 15810 19128
rect 16025 19125 16037 19128
rect 16071 19125 16083 19159
rect 16025 19119 16083 19125
rect 16117 19159 16175 19165
rect 16117 19125 16129 19159
rect 16163 19156 16175 19159
rect 16574 19156 16580 19168
rect 16163 19128 16580 19156
rect 16163 19125 16175 19128
rect 16117 19119 16175 19125
rect 16574 19116 16580 19128
rect 16632 19116 16638 19168
rect 16758 19156 16764 19168
rect 16719 19128 16764 19156
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 16942 19156 16948 19168
rect 16903 19128 16948 19156
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 19334 19156 19340 19168
rect 19295 19128 19340 19156
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 19426 19116 19432 19168
rect 19484 19156 19490 19168
rect 21269 19159 21327 19165
rect 19484 19128 19529 19156
rect 19484 19116 19490 19128
rect 21269 19125 21281 19159
rect 21315 19156 21327 19159
rect 21358 19156 21364 19168
rect 21315 19128 21364 19156
rect 21315 19125 21327 19128
rect 21269 19119 21327 19125
rect 21358 19116 21364 19128
rect 21416 19156 21422 19168
rect 21744 19156 21772 19196
rect 22649 19193 22661 19196
rect 22695 19193 22707 19227
rect 22649 19187 22707 19193
rect 21416 19128 21772 19156
rect 21416 19116 21422 19128
rect 21910 19116 21916 19168
rect 21968 19156 21974 19168
rect 22189 19159 22247 19165
rect 22189 19156 22201 19159
rect 21968 19128 22201 19156
rect 21968 19116 21974 19128
rect 22189 19125 22201 19128
rect 22235 19125 22247 19159
rect 23014 19156 23020 19168
rect 22975 19128 23020 19156
rect 22189 19119 22247 19125
rect 23014 19116 23020 19128
rect 23072 19116 23078 19168
rect 1104 19066 23460 19088
rect 1104 19014 8446 19066
rect 8498 19014 8510 19066
rect 8562 19014 8574 19066
rect 8626 19014 8638 19066
rect 8690 19014 15910 19066
rect 15962 19014 15974 19066
rect 16026 19014 16038 19066
rect 16090 19014 16102 19066
rect 16154 19014 23460 19066
rect 1104 18992 23460 19014
rect 1765 18955 1823 18961
rect 1765 18921 1777 18955
rect 1811 18952 1823 18955
rect 1946 18952 1952 18964
rect 1811 18924 1952 18952
rect 1811 18921 1823 18924
rect 1765 18915 1823 18921
rect 1946 18912 1952 18924
rect 2004 18952 2010 18964
rect 4157 18955 4215 18961
rect 4157 18952 4169 18955
rect 2004 18924 4169 18952
rect 2004 18912 2010 18924
rect 4157 18921 4169 18924
rect 4203 18921 4215 18955
rect 4157 18915 4215 18921
rect 4338 18912 4344 18964
rect 4396 18952 4402 18964
rect 4617 18955 4675 18961
rect 4617 18952 4629 18955
rect 4396 18924 4629 18952
rect 4396 18912 4402 18924
rect 4617 18921 4629 18924
rect 4663 18921 4675 18955
rect 4617 18915 4675 18921
rect 4985 18955 5043 18961
rect 4985 18921 4997 18955
rect 5031 18952 5043 18955
rect 5074 18952 5080 18964
rect 5031 18924 5080 18952
rect 5031 18921 5043 18924
rect 4985 18915 5043 18921
rect 5074 18912 5080 18924
rect 5132 18912 5138 18964
rect 5258 18952 5264 18964
rect 5219 18924 5264 18952
rect 5258 18912 5264 18924
rect 5316 18912 5322 18964
rect 8110 18912 8116 18964
rect 8168 18952 8174 18964
rect 8573 18955 8631 18961
rect 8573 18952 8585 18955
rect 8168 18924 8585 18952
rect 8168 18912 8174 18924
rect 8573 18921 8585 18924
rect 8619 18921 8631 18955
rect 8573 18915 8631 18921
rect 8941 18955 8999 18961
rect 8941 18921 8953 18955
rect 8987 18952 8999 18955
rect 9766 18952 9772 18964
rect 8987 18924 9772 18952
rect 8987 18921 8999 18924
rect 8941 18915 8999 18921
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 10778 18912 10784 18964
rect 10836 18952 10842 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 10836 18924 11069 18952
rect 10836 18912 10842 18924
rect 11057 18921 11069 18924
rect 11103 18921 11115 18955
rect 11057 18915 11115 18921
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11517 18955 11575 18961
rect 11517 18952 11529 18955
rect 11204 18924 11529 18952
rect 11204 18912 11210 18924
rect 11517 18921 11529 18924
rect 11563 18921 11575 18955
rect 13262 18952 13268 18964
rect 13223 18924 13268 18952
rect 11517 18915 11575 18921
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 14185 18955 14243 18961
rect 14185 18921 14197 18955
rect 14231 18921 14243 18955
rect 14550 18952 14556 18964
rect 14511 18924 14556 18952
rect 14185 18915 14243 18921
rect 2130 18844 2136 18896
rect 2188 18884 2194 18896
rect 2188 18856 3004 18884
rect 2188 18844 2194 18856
rect 2314 18776 2320 18828
rect 2372 18816 2378 18828
rect 2878 18819 2936 18825
rect 2878 18816 2890 18819
rect 2372 18788 2890 18816
rect 2372 18776 2378 18788
rect 2878 18785 2890 18788
rect 2924 18785 2936 18819
rect 2976 18816 3004 18856
rect 3050 18844 3056 18896
rect 3108 18884 3114 18896
rect 4249 18887 4307 18893
rect 4249 18884 4261 18887
rect 3108 18856 4261 18884
rect 3108 18844 3114 18856
rect 4249 18853 4261 18856
rect 4295 18853 4307 18887
rect 4249 18847 4307 18853
rect 5629 18887 5687 18893
rect 5629 18853 5641 18887
rect 5675 18884 5687 18887
rect 6178 18884 6184 18896
rect 5675 18856 6184 18884
rect 5675 18853 5687 18856
rect 5629 18847 5687 18853
rect 6178 18844 6184 18856
rect 6236 18844 6242 18896
rect 7834 18844 7840 18896
rect 7892 18893 7898 18896
rect 7892 18884 7904 18893
rect 8481 18887 8539 18893
rect 7892 18856 7937 18884
rect 7892 18847 7904 18856
rect 8481 18853 8493 18887
rect 8527 18884 8539 18887
rect 9122 18884 9128 18896
rect 8527 18856 9128 18884
rect 8527 18853 8539 18856
rect 8481 18847 8539 18853
rect 7892 18844 7898 18847
rect 9122 18844 9128 18856
rect 9180 18844 9186 18896
rect 11425 18887 11483 18893
rect 11425 18853 11437 18887
rect 11471 18884 11483 18887
rect 11698 18884 11704 18896
rect 11471 18856 11704 18884
rect 11471 18853 11483 18856
rect 11425 18847 11483 18853
rect 11698 18844 11704 18856
rect 11756 18844 11762 18896
rect 13998 18884 14004 18896
rect 13648 18856 14004 18884
rect 3145 18819 3203 18825
rect 3145 18816 3157 18819
rect 2976 18788 3157 18816
rect 2878 18779 2936 18785
rect 3145 18785 3157 18788
rect 3191 18816 3203 18819
rect 3602 18816 3608 18828
rect 3191 18788 3608 18816
rect 3191 18785 3203 18788
rect 3145 18779 3203 18785
rect 3602 18776 3608 18788
rect 3660 18776 3666 18828
rect 4798 18816 4804 18828
rect 4759 18788 4804 18816
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 6089 18819 6147 18825
rect 6089 18785 6101 18819
rect 6135 18816 6147 18819
rect 6362 18816 6368 18828
rect 6135 18788 6368 18816
rect 6135 18785 6147 18788
rect 6089 18779 6147 18785
rect 6362 18776 6368 18788
rect 6420 18776 6426 18828
rect 7374 18776 7380 18828
rect 7432 18816 7438 18828
rect 9140 18816 9168 18844
rect 9861 18819 9919 18825
rect 7432 18788 9076 18816
rect 9140 18788 9812 18816
rect 7432 18776 7438 18788
rect 9048 18760 9076 18788
rect 4065 18751 4123 18757
rect 4065 18717 4077 18751
rect 4111 18748 4123 18751
rect 4430 18748 4436 18760
rect 4111 18720 4436 18748
rect 4111 18717 4123 18720
rect 4065 18711 4123 18717
rect 4430 18708 4436 18720
rect 4488 18708 4494 18760
rect 5074 18708 5080 18760
rect 5132 18748 5138 18760
rect 5721 18751 5779 18757
rect 5721 18748 5733 18751
rect 5132 18720 5733 18748
rect 5132 18708 5138 18720
rect 5721 18717 5733 18720
rect 5767 18717 5779 18751
rect 5721 18711 5779 18717
rect 5905 18751 5963 18757
rect 5905 18717 5917 18751
rect 5951 18748 5963 18751
rect 6822 18748 6828 18760
rect 5951 18720 6828 18748
rect 5951 18717 5963 18720
rect 5905 18711 5963 18717
rect 6822 18708 6828 18720
rect 6880 18708 6886 18760
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18717 8171 18751
rect 8294 18748 8300 18760
rect 8255 18720 8300 18748
rect 8113 18711 8171 18717
rect 8128 18680 8156 18711
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 9030 18748 9036 18760
rect 8943 18720 9036 18748
rect 9030 18708 9036 18720
rect 9088 18748 9094 18760
rect 9125 18751 9183 18757
rect 9125 18748 9137 18751
rect 9088 18720 9137 18748
rect 9088 18708 9094 18720
rect 9125 18717 9137 18720
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 9306 18708 9312 18760
rect 9364 18748 9370 18760
rect 9674 18757 9680 18760
rect 9448 18751 9506 18757
rect 9448 18748 9460 18751
rect 9364 18720 9460 18748
rect 9364 18708 9370 18720
rect 9448 18717 9460 18720
rect 9494 18717 9506 18751
rect 9448 18711 9506 18717
rect 9631 18751 9680 18757
rect 9631 18717 9643 18751
rect 9677 18717 9680 18751
rect 9631 18711 9680 18717
rect 9674 18708 9680 18711
rect 9732 18708 9738 18760
rect 9784 18748 9812 18788
rect 9861 18785 9873 18819
rect 9907 18816 9919 18819
rect 10134 18816 10140 18828
rect 9907 18788 10140 18816
rect 9907 18785 9919 18788
rect 9861 18779 9919 18785
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 12158 18825 12164 18828
rect 12152 18816 12164 18825
rect 11112 18788 11652 18816
rect 12119 18788 12164 18816
rect 11112 18776 11118 18788
rect 10318 18748 10324 18760
rect 9784 18720 10324 18748
rect 10318 18708 10324 18720
rect 10376 18708 10382 18760
rect 11624 18757 11652 18788
rect 12152 18779 12164 18788
rect 12158 18776 12164 18779
rect 12216 18776 12222 18828
rect 11609 18751 11667 18757
rect 11609 18717 11621 18751
rect 11655 18717 11667 18751
rect 11609 18711 11667 18717
rect 11790 18708 11796 18760
rect 11848 18748 11854 18760
rect 13648 18757 13676 18856
rect 13998 18844 14004 18856
rect 14056 18844 14062 18896
rect 13817 18819 13875 18825
rect 13817 18785 13829 18819
rect 13863 18816 13875 18819
rect 13906 18816 13912 18828
rect 13863 18788 13912 18816
rect 13863 18785 13875 18788
rect 13817 18779 13875 18785
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 14200 18816 14228 18915
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 14826 18952 14832 18964
rect 14787 18924 14832 18952
rect 14826 18912 14832 18924
rect 14884 18912 14890 18964
rect 16758 18912 16764 18964
rect 16816 18952 16822 18964
rect 16816 18924 19012 18952
rect 16816 18912 16822 18924
rect 15378 18844 15384 18896
rect 15436 18884 15442 18896
rect 16485 18887 16543 18893
rect 16485 18884 16497 18887
rect 15436 18856 16497 18884
rect 15436 18844 15442 18856
rect 16485 18853 16497 18856
rect 16531 18853 16543 18887
rect 16485 18847 16543 18853
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 14200 18788 14381 18816
rect 14369 18785 14381 18788
rect 14415 18785 14427 18819
rect 14642 18816 14648 18828
rect 14603 18788 14648 18816
rect 14369 18779 14427 18785
rect 14642 18776 14648 18788
rect 14700 18776 14706 18828
rect 14734 18776 14740 18828
rect 14792 18816 14798 18828
rect 15194 18825 15200 18828
rect 15177 18819 15200 18825
rect 15177 18816 15189 18819
rect 14792 18788 15189 18816
rect 14792 18776 14798 18788
rect 15177 18785 15189 18788
rect 15252 18816 15258 18828
rect 16500 18816 16528 18847
rect 18230 18844 18236 18896
rect 18288 18884 18294 18896
rect 18984 18893 19012 18924
rect 20070 18912 20076 18964
rect 20128 18952 20134 18964
rect 20438 18952 20444 18964
rect 20128 18924 20444 18952
rect 20128 18912 20134 18924
rect 20438 18912 20444 18924
rect 20496 18912 20502 18964
rect 22370 18912 22376 18964
rect 22428 18952 22434 18964
rect 22465 18955 22523 18961
rect 22465 18952 22477 18955
rect 22428 18924 22477 18952
rect 22428 18912 22434 18924
rect 22465 18921 22477 18924
rect 22511 18921 22523 18955
rect 22465 18915 22523 18921
rect 21358 18893 21364 18896
rect 18785 18887 18843 18893
rect 18785 18884 18797 18887
rect 18288 18856 18797 18884
rect 18288 18844 18294 18856
rect 18785 18853 18797 18856
rect 18831 18853 18843 18887
rect 18785 18847 18843 18853
rect 18969 18887 19027 18893
rect 18969 18853 18981 18887
rect 19015 18853 19027 18887
rect 21352 18884 21364 18893
rect 21319 18856 21364 18884
rect 18969 18847 19027 18853
rect 21352 18847 21364 18856
rect 21358 18844 21364 18847
rect 21416 18844 21422 18896
rect 21726 18844 21732 18896
rect 21784 18884 21790 18896
rect 23014 18884 23020 18896
rect 21784 18856 23020 18884
rect 21784 18844 21790 18856
rect 23014 18844 23020 18856
rect 23072 18844 23078 18896
rect 16992 18819 17050 18825
rect 16992 18816 17004 18819
rect 15252 18788 15325 18816
rect 16500 18788 17004 18816
rect 15177 18779 15200 18785
rect 15194 18776 15200 18779
rect 15252 18776 15258 18788
rect 16992 18785 17004 18788
rect 17038 18785 17050 18819
rect 17402 18816 17408 18828
rect 17363 18788 17408 18816
rect 16992 18779 17050 18785
rect 17402 18776 17408 18788
rect 17460 18776 17466 18828
rect 19880 18819 19938 18825
rect 19880 18785 19892 18819
rect 19926 18816 19938 18819
rect 20438 18816 20444 18828
rect 19926 18788 20444 18816
rect 19926 18785 19938 18788
rect 19880 18779 19938 18785
rect 20438 18776 20444 18788
rect 20496 18776 20502 18828
rect 11885 18751 11943 18757
rect 11885 18748 11897 18751
rect 11848 18720 11897 18748
rect 11848 18708 11854 18720
rect 11885 18717 11897 18720
rect 11931 18717 11943 18751
rect 11885 18711 11943 18717
rect 13633 18751 13691 18757
rect 13633 18717 13645 18751
rect 13679 18717 13691 18751
rect 13633 18711 13691 18717
rect 13725 18751 13783 18757
rect 13725 18717 13737 18751
rect 13771 18748 13783 18751
rect 14918 18748 14924 18760
rect 13771 18720 13860 18748
rect 14879 18720 14924 18748
rect 13771 18717 13783 18720
rect 13725 18711 13783 18717
rect 8754 18680 8760 18692
rect 8128 18652 8760 18680
rect 8312 18624 8340 18652
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 10962 18680 10968 18692
rect 10923 18652 10968 18680
rect 10962 18640 10968 18652
rect 11020 18640 11026 18692
rect 1578 18572 1584 18624
rect 1636 18612 1642 18624
rect 4522 18612 4528 18624
rect 1636 18584 4528 18612
rect 1636 18572 1642 18584
rect 4522 18572 4528 18584
rect 4580 18572 4586 18624
rect 6086 18572 6092 18624
rect 6144 18612 6150 18624
rect 6273 18615 6331 18621
rect 6273 18612 6285 18615
rect 6144 18584 6285 18612
rect 6144 18572 6150 18584
rect 6273 18581 6285 18584
rect 6319 18581 6331 18615
rect 6273 18575 6331 18581
rect 6733 18615 6791 18621
rect 6733 18581 6745 18615
rect 6779 18612 6791 18615
rect 7926 18612 7932 18624
rect 6779 18584 7932 18612
rect 6779 18581 6791 18584
rect 6733 18575 6791 18581
rect 7926 18572 7932 18584
rect 7984 18572 7990 18624
rect 8294 18572 8300 18624
rect 8352 18572 8358 18624
rect 8386 18572 8392 18624
rect 8444 18612 8450 18624
rect 9490 18612 9496 18624
rect 8444 18584 9496 18612
rect 8444 18572 8450 18584
rect 9490 18572 9496 18584
rect 9548 18612 9554 18624
rect 10980 18612 11008 18640
rect 9548 18584 11008 18612
rect 11900 18612 11928 18711
rect 13832 18692 13860 18720
rect 14918 18708 14924 18720
rect 14976 18708 14982 18760
rect 16206 18708 16212 18760
rect 16264 18748 16270 18760
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 16264 18720 16681 18748
rect 16264 18708 16270 18720
rect 16669 18717 16681 18720
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 17126 18708 17132 18760
rect 17184 18748 17190 18760
rect 18693 18751 18751 18757
rect 18693 18748 18705 18751
rect 17184 18720 17229 18748
rect 18064 18720 18705 18748
rect 17184 18708 17190 18720
rect 13814 18640 13820 18692
rect 13872 18640 13878 18692
rect 13078 18612 13084 18624
rect 11900 18584 13084 18612
rect 9548 18572 9554 18584
rect 13078 18572 13084 18584
rect 13136 18572 13142 18624
rect 14366 18572 14372 18624
rect 14424 18612 14430 18624
rect 14936 18612 14964 18708
rect 16301 18683 16359 18689
rect 16301 18649 16313 18683
rect 16347 18680 16359 18683
rect 16574 18680 16580 18692
rect 16347 18652 16580 18680
rect 16347 18649 16359 18652
rect 16301 18643 16359 18649
rect 16574 18640 16580 18652
rect 16632 18640 16638 18692
rect 16114 18612 16120 18624
rect 14424 18584 16120 18612
rect 14424 18572 14430 18584
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16942 18572 16948 18624
rect 17000 18612 17006 18624
rect 18064 18612 18092 18720
rect 18693 18717 18705 18720
rect 18739 18717 18751 18751
rect 18693 18711 18751 18717
rect 19150 18708 19156 18760
rect 19208 18748 19214 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19208 18720 19625 18748
rect 19208 18708 19214 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 20990 18708 20996 18760
rect 21048 18748 21054 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 21048 18720 21097 18748
rect 21048 18708 21054 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 19242 18680 19248 18692
rect 19203 18652 19248 18680
rect 19242 18640 19248 18652
rect 19300 18640 19306 18692
rect 17000 18584 18092 18612
rect 17000 18572 17006 18584
rect 18322 18572 18328 18624
rect 18380 18612 18386 18624
rect 18509 18615 18567 18621
rect 18509 18612 18521 18615
rect 18380 18584 18521 18612
rect 18380 18572 18386 18584
rect 18509 18581 18521 18584
rect 18555 18581 18567 18615
rect 18509 18575 18567 18581
rect 20346 18572 20352 18624
rect 20404 18612 20410 18624
rect 20993 18615 21051 18621
rect 20993 18612 21005 18615
rect 20404 18584 21005 18612
rect 20404 18572 20410 18584
rect 20993 18581 21005 18584
rect 21039 18581 21051 18615
rect 20993 18575 21051 18581
rect 1104 18522 23460 18544
rect 1104 18470 4714 18522
rect 4766 18470 4778 18522
rect 4830 18470 4842 18522
rect 4894 18470 4906 18522
rect 4958 18470 12178 18522
rect 12230 18470 12242 18522
rect 12294 18470 12306 18522
rect 12358 18470 12370 18522
rect 12422 18470 19642 18522
rect 19694 18470 19706 18522
rect 19758 18470 19770 18522
rect 19822 18470 19834 18522
rect 19886 18470 23460 18522
rect 1104 18448 23460 18470
rect 2222 18408 2228 18420
rect 2183 18380 2228 18408
rect 2222 18368 2228 18380
rect 2280 18368 2286 18420
rect 3602 18368 3608 18420
rect 3660 18408 3666 18420
rect 4709 18411 4767 18417
rect 3660 18380 4568 18408
rect 3660 18368 3666 18380
rect 3697 18343 3755 18349
rect 3697 18340 3709 18343
rect 3620 18312 3709 18340
rect 1578 18272 1584 18284
rect 1539 18244 1584 18272
rect 1578 18232 1584 18244
rect 1636 18232 1642 18284
rect 3620 18272 3648 18312
rect 3697 18309 3709 18312
rect 3743 18309 3755 18343
rect 3697 18303 3755 18309
rect 3528 18244 3648 18272
rect 4341 18275 4399 18281
rect 1673 18207 1731 18213
rect 1673 18173 1685 18207
rect 1719 18204 1731 18207
rect 3050 18204 3056 18216
rect 1719 18176 3056 18204
rect 1719 18173 1731 18176
rect 1673 18167 1731 18173
rect 3050 18164 3056 18176
rect 3108 18164 3114 18216
rect 3326 18164 3332 18216
rect 3384 18213 3390 18216
rect 3384 18204 3396 18213
rect 3384 18176 3429 18204
rect 3384 18167 3396 18176
rect 3384 18164 3390 18167
rect 1765 18139 1823 18145
rect 1765 18105 1777 18139
rect 1811 18136 1823 18139
rect 3528 18136 3556 18244
rect 4341 18241 4353 18275
rect 4387 18272 4399 18275
rect 4430 18272 4436 18284
rect 4387 18244 4436 18272
rect 4387 18241 4399 18244
rect 4341 18235 4399 18241
rect 4430 18232 4436 18244
rect 4488 18232 4494 18284
rect 4540 18272 4568 18380
rect 4709 18377 4721 18411
rect 4755 18408 4767 18411
rect 5166 18408 5172 18420
rect 4755 18380 5172 18408
rect 4755 18377 4767 18380
rect 4709 18371 4767 18377
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 7193 18411 7251 18417
rect 7193 18377 7205 18411
rect 7239 18408 7251 18411
rect 7650 18408 7656 18420
rect 7239 18380 7656 18408
rect 7239 18377 7251 18380
rect 7193 18371 7251 18377
rect 7650 18368 7656 18380
rect 7708 18368 7714 18420
rect 9677 18411 9735 18417
rect 9677 18377 9689 18411
rect 9723 18408 9735 18411
rect 10042 18408 10048 18420
rect 9723 18380 10048 18408
rect 9723 18377 9735 18380
rect 9677 18371 9735 18377
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 13906 18408 13912 18420
rect 10152 18380 11560 18408
rect 9030 18300 9036 18352
rect 9088 18340 9094 18352
rect 10152 18340 10180 18380
rect 9088 18312 10180 18340
rect 9088 18300 9094 18312
rect 4614 18272 4620 18284
rect 4527 18244 4620 18272
rect 4614 18232 4620 18244
rect 4672 18272 4678 18284
rect 4801 18275 4859 18281
rect 4801 18272 4813 18275
rect 4672 18244 4813 18272
rect 4672 18232 4678 18244
rect 4801 18241 4813 18244
rect 4847 18241 4859 18275
rect 4801 18235 4859 18241
rect 8297 18275 8355 18281
rect 8297 18241 8309 18275
rect 8343 18272 8355 18275
rect 8386 18272 8392 18284
rect 8343 18244 8392 18272
rect 8343 18241 8355 18244
rect 8297 18235 8355 18241
rect 3602 18213 3608 18216
rect 3598 18167 3608 18213
rect 3660 18204 3666 18216
rect 3660 18176 3698 18204
rect 3602 18164 3608 18167
rect 3660 18164 3666 18176
rect 3786 18164 3792 18216
rect 3844 18204 3850 18216
rect 4157 18207 4215 18213
rect 4157 18204 4169 18207
rect 3844 18176 4169 18204
rect 3844 18164 3850 18176
rect 4157 18173 4169 18176
rect 4203 18173 4215 18207
rect 4157 18167 4215 18173
rect 4525 18207 4583 18213
rect 4525 18173 4537 18207
rect 4571 18173 4583 18207
rect 4525 18167 4583 18173
rect 4540 18136 4568 18167
rect 1811 18108 3556 18136
rect 3804 18108 4568 18136
rect 4816 18136 4844 18235
rect 8386 18232 8392 18244
rect 8444 18232 8450 18284
rect 8570 18275 8628 18281
rect 8570 18241 8582 18275
rect 8616 18272 8628 18275
rect 8754 18272 8760 18284
rect 8616 18244 8760 18272
rect 8616 18241 8628 18244
rect 8570 18235 8628 18241
rect 8754 18232 8760 18244
rect 8812 18232 8818 18284
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18272 9643 18275
rect 10870 18272 10876 18284
rect 9631 18244 10876 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 11054 18275 11112 18281
rect 11054 18241 11066 18275
rect 11100 18272 11112 18275
rect 11238 18272 11244 18284
rect 11100 18244 11244 18272
rect 11100 18241 11112 18244
rect 11054 18235 11112 18241
rect 11238 18232 11244 18244
rect 11296 18232 11302 18284
rect 5074 18213 5080 18216
rect 5068 18204 5080 18213
rect 5035 18176 5080 18204
rect 5068 18167 5080 18176
rect 5074 18164 5080 18167
rect 5132 18164 5138 18216
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 9088 18176 9133 18204
rect 9088 18164 9094 18176
rect 9214 18164 9220 18216
rect 9272 18204 9278 18216
rect 9674 18204 9680 18216
rect 9272 18176 9680 18204
rect 9272 18164 9278 18176
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 11532 18213 11560 18380
rect 11624 18380 13768 18408
rect 13867 18380 13912 18408
rect 10781 18207 10839 18213
rect 10781 18173 10793 18207
rect 10827 18204 10839 18207
rect 11517 18207 11575 18213
rect 10827 18176 11468 18204
rect 10827 18173 10839 18176
rect 10781 18167 10839 18173
rect 6086 18136 6092 18148
rect 4816 18108 6092 18136
rect 1811 18105 1823 18108
rect 1765 18099 1823 18105
rect 2133 18071 2191 18077
rect 2133 18037 2145 18071
rect 2179 18068 2191 18071
rect 3804 18068 3832 18108
rect 6086 18096 6092 18108
rect 6144 18096 6150 18148
rect 11440 18136 11468 18176
rect 11517 18173 11529 18207
rect 11563 18173 11575 18207
rect 11517 18167 11575 18173
rect 11624 18136 11652 18380
rect 11701 18343 11759 18349
rect 11701 18309 11713 18343
rect 11747 18340 11759 18343
rect 12066 18340 12072 18352
rect 11747 18312 12072 18340
rect 11747 18309 11759 18312
rect 11701 18303 11759 18309
rect 12066 18300 12072 18312
rect 12124 18300 12130 18352
rect 13740 18340 13768 18380
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 14734 18408 14740 18420
rect 14695 18380 14740 18408
rect 14734 18368 14740 18380
rect 14792 18368 14798 18420
rect 16666 18408 16672 18420
rect 14844 18380 16672 18408
rect 14844 18340 14872 18380
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 18230 18408 18236 18420
rect 18191 18380 18236 18408
rect 18230 18368 18236 18380
rect 18288 18368 18294 18420
rect 20349 18411 20407 18417
rect 20349 18377 20361 18411
rect 20395 18408 20407 18411
rect 22462 18408 22468 18420
rect 20395 18380 22468 18408
rect 20395 18377 20407 18380
rect 20349 18371 20407 18377
rect 22462 18368 22468 18380
rect 22520 18368 22526 18420
rect 13740 18312 14872 18340
rect 16393 18343 16451 18349
rect 16393 18309 16405 18343
rect 16439 18309 16451 18343
rect 16393 18303 16451 18309
rect 13078 18272 13084 18284
rect 13039 18244 13084 18272
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 13722 18232 13728 18284
rect 13780 18272 13786 18284
rect 14461 18275 14519 18281
rect 14461 18272 14473 18275
rect 13780 18244 14473 18272
rect 13780 18232 13786 18244
rect 14461 18241 14473 18244
rect 14507 18241 14519 18275
rect 16114 18272 16120 18284
rect 16075 18244 16120 18272
rect 14461 18235 14519 18241
rect 16114 18232 16120 18244
rect 16172 18272 16178 18284
rect 16298 18272 16304 18284
rect 16172 18244 16304 18272
rect 16172 18232 16178 18244
rect 16298 18232 16304 18244
rect 16356 18272 16362 18284
rect 16408 18272 16436 18303
rect 16850 18300 16856 18352
rect 16908 18340 16914 18352
rect 18417 18343 18475 18349
rect 18417 18340 18429 18343
rect 16908 18312 18429 18340
rect 16908 18300 16914 18312
rect 18417 18309 18429 18312
rect 18463 18309 18475 18343
rect 18417 18303 18475 18309
rect 17586 18272 17592 18284
rect 16356 18244 16436 18272
rect 17547 18244 17592 18272
rect 16356 18232 16362 18244
rect 17586 18232 17592 18244
rect 17644 18232 17650 18284
rect 17678 18232 17684 18284
rect 17736 18272 17742 18284
rect 18693 18275 18751 18281
rect 18693 18272 18705 18275
rect 17736 18244 18705 18272
rect 17736 18232 17742 18244
rect 18693 18241 18705 18244
rect 18739 18241 18751 18275
rect 22830 18272 22836 18284
rect 22791 18244 22836 18272
rect 18693 18235 18751 18241
rect 15286 18164 15292 18216
rect 15344 18204 15350 18216
rect 15850 18207 15908 18213
rect 15850 18204 15862 18207
rect 15344 18176 15862 18204
rect 15344 18164 15350 18176
rect 15850 18173 15862 18176
rect 15896 18173 15908 18207
rect 15850 18167 15908 18173
rect 16209 18207 16267 18213
rect 16209 18173 16221 18207
rect 16255 18173 16267 18207
rect 16209 18167 16267 18173
rect 11440 18108 11652 18136
rect 12836 18139 12894 18145
rect 12836 18105 12848 18139
rect 12882 18136 12894 18139
rect 15470 18136 15476 18148
rect 12882 18108 15476 18136
rect 12882 18105 12894 18108
rect 12836 18099 12894 18105
rect 15470 18096 15476 18108
rect 15528 18096 15534 18148
rect 15562 18096 15568 18148
rect 15620 18136 15626 18148
rect 16224 18136 16252 18167
rect 17126 18164 17132 18216
rect 17184 18204 17190 18216
rect 17865 18207 17923 18213
rect 17865 18204 17877 18207
rect 17184 18176 17877 18204
rect 17184 18164 17190 18176
rect 17865 18173 17877 18176
rect 17911 18173 17923 18207
rect 17865 18167 17923 18173
rect 17954 18164 17960 18216
rect 18012 18204 18018 18216
rect 18601 18207 18659 18213
rect 18601 18204 18613 18207
rect 18012 18176 18613 18204
rect 18012 18164 18018 18176
rect 18601 18173 18613 18176
rect 18647 18173 18659 18207
rect 18601 18167 18659 18173
rect 15620 18108 16252 18136
rect 18708 18136 18736 18235
rect 22830 18232 22836 18244
rect 22888 18232 22894 18284
rect 18960 18207 19018 18213
rect 18960 18173 18972 18207
rect 19006 18204 19018 18207
rect 19426 18204 19432 18216
rect 19006 18176 19432 18204
rect 19006 18173 19018 18176
rect 18960 18167 19018 18173
rect 19426 18164 19432 18176
rect 19484 18204 19490 18216
rect 19702 18204 19708 18216
rect 19484 18176 19708 18204
rect 19484 18164 19490 18176
rect 19702 18164 19708 18176
rect 19760 18164 19766 18216
rect 20162 18204 20168 18216
rect 20123 18176 20168 18204
rect 20162 18164 20168 18176
rect 20220 18164 20226 18216
rect 20625 18207 20683 18213
rect 20625 18173 20637 18207
rect 20671 18173 20683 18207
rect 20625 18167 20683 18173
rect 20892 18207 20950 18213
rect 20892 18173 20904 18207
rect 20938 18204 20950 18207
rect 22557 18207 22615 18213
rect 22557 18204 22569 18207
rect 20938 18176 22569 18204
rect 20938 18173 20950 18176
rect 20892 18167 20950 18173
rect 22557 18173 22569 18176
rect 22603 18204 22615 18207
rect 22646 18204 22652 18216
rect 22603 18176 22652 18204
rect 22603 18173 22615 18176
rect 22557 18167 22615 18173
rect 19150 18136 19156 18148
rect 18708 18108 19156 18136
rect 15620 18096 15626 18108
rect 19150 18096 19156 18108
rect 19208 18136 19214 18148
rect 20640 18136 20668 18167
rect 22646 18164 22652 18176
rect 22704 18164 22710 18216
rect 20990 18136 20996 18148
rect 19208 18108 20996 18136
rect 19208 18096 19214 18108
rect 20990 18096 20996 18108
rect 21048 18096 21054 18148
rect 21358 18096 21364 18148
rect 21416 18136 21422 18148
rect 21416 18108 22232 18136
rect 21416 18096 21422 18108
rect 4062 18068 4068 18080
rect 2179 18040 3832 18068
rect 4023 18040 4068 18068
rect 2179 18037 2191 18040
rect 2133 18031 2191 18037
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 6178 18068 6184 18080
rect 6139 18040 6184 18068
rect 6178 18028 6184 18040
rect 6236 18028 6242 18080
rect 6914 18068 6920 18080
rect 6875 18040 6920 18068
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 8566 18071 8624 18077
rect 8566 18037 8578 18071
rect 8612 18068 8624 18071
rect 9217 18071 9275 18077
rect 9217 18068 9229 18071
rect 8612 18040 9229 18068
rect 8612 18037 8624 18040
rect 8566 18031 8624 18037
rect 9217 18037 9229 18040
rect 9263 18068 9275 18071
rect 9306 18068 9312 18080
rect 9263 18040 9312 18068
rect 9263 18037 9275 18040
rect 9217 18031 9275 18037
rect 9306 18028 9312 18040
rect 9364 18068 9370 18080
rect 11050 18071 11108 18077
rect 11050 18068 11062 18071
rect 9364 18040 11062 18068
rect 9364 18028 9370 18040
rect 11050 18037 11062 18040
rect 11096 18037 11108 18071
rect 11050 18031 11108 18037
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 13173 18071 13231 18077
rect 13173 18068 13185 18071
rect 12768 18040 13185 18068
rect 12768 18028 12774 18040
rect 13173 18037 13185 18040
rect 13219 18037 13231 18071
rect 14274 18068 14280 18080
rect 14235 18040 14280 18068
rect 13173 18031 13231 18037
rect 14274 18028 14280 18040
rect 14332 18028 14338 18080
rect 14369 18071 14427 18077
rect 14369 18037 14381 18071
rect 14415 18068 14427 18071
rect 14826 18068 14832 18080
rect 14415 18040 14832 18068
rect 14415 18037 14427 18040
rect 14369 18031 14427 18037
rect 14826 18028 14832 18040
rect 14884 18028 14890 18080
rect 17218 18068 17224 18080
rect 17179 18040 17224 18068
rect 17218 18028 17224 18040
rect 17276 18028 17282 18080
rect 17402 18068 17408 18080
rect 17363 18040 17408 18068
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 17773 18071 17831 18077
rect 17773 18037 17785 18071
rect 17819 18068 17831 18071
rect 18230 18068 18236 18080
rect 17819 18040 18236 18068
rect 17819 18037 17831 18040
rect 17773 18031 17831 18037
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 20073 18071 20131 18077
rect 20073 18037 20085 18071
rect 20119 18068 20131 18071
rect 20438 18068 20444 18080
rect 20119 18040 20444 18068
rect 20119 18037 20131 18040
rect 20073 18031 20131 18037
rect 20438 18028 20444 18040
rect 20496 18028 20502 18080
rect 22002 18068 22008 18080
rect 21963 18040 22008 18068
rect 22002 18028 22008 18040
rect 22060 18028 22066 18080
rect 22204 18077 22232 18108
rect 22189 18071 22247 18077
rect 22189 18037 22201 18071
rect 22235 18037 22247 18071
rect 22189 18031 22247 18037
rect 22554 18028 22560 18080
rect 22612 18068 22618 18080
rect 22649 18071 22707 18077
rect 22649 18068 22661 18071
rect 22612 18040 22661 18068
rect 22612 18028 22618 18040
rect 22649 18037 22661 18040
rect 22695 18037 22707 18071
rect 22649 18031 22707 18037
rect 1104 17978 23460 18000
rect 1104 17926 8446 17978
rect 8498 17926 8510 17978
rect 8562 17926 8574 17978
rect 8626 17926 8638 17978
rect 8690 17926 15910 17978
rect 15962 17926 15974 17978
rect 16026 17926 16038 17978
rect 16090 17926 16102 17978
rect 16154 17926 23460 17978
rect 1104 17904 23460 17926
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 3881 17867 3939 17873
rect 3881 17864 3893 17867
rect 3108 17836 3893 17864
rect 3108 17824 3114 17836
rect 3881 17833 3893 17836
rect 3927 17833 3939 17867
rect 3881 17827 3939 17833
rect 4801 17867 4859 17873
rect 4801 17833 4813 17867
rect 4847 17864 4859 17867
rect 5074 17864 5080 17876
rect 4847 17836 5080 17864
rect 4847 17833 4859 17836
rect 4801 17827 4859 17833
rect 5074 17824 5080 17836
rect 5132 17824 5138 17876
rect 6822 17864 6828 17876
rect 5184 17836 6828 17864
rect 2400 17799 2458 17805
rect 2400 17765 2412 17799
rect 2446 17796 2458 17799
rect 3418 17796 3424 17808
rect 2446 17768 3424 17796
rect 2446 17765 2458 17768
rect 2400 17759 2458 17765
rect 3418 17756 3424 17768
rect 3476 17796 3482 17808
rect 3786 17796 3792 17808
rect 3476 17768 3792 17796
rect 3476 17756 3482 17768
rect 3786 17756 3792 17768
rect 3844 17756 3850 17808
rect 1762 17688 1768 17740
rect 1820 17728 1826 17740
rect 4249 17731 4307 17737
rect 4249 17728 4261 17731
rect 1820 17700 4261 17728
rect 1820 17688 1826 17700
rect 4249 17697 4261 17700
rect 4295 17697 4307 17731
rect 4249 17691 4307 17697
rect 2130 17660 2136 17672
rect 2091 17632 2136 17660
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 3234 17620 3240 17672
rect 3292 17660 3298 17672
rect 4341 17663 4399 17669
rect 4341 17660 4353 17663
rect 3292 17632 4353 17660
rect 3292 17620 3298 17632
rect 4341 17629 4353 17632
rect 4387 17629 4399 17663
rect 4341 17623 4399 17629
rect 4430 17620 4436 17672
rect 4488 17660 4494 17672
rect 4525 17663 4583 17669
rect 4525 17660 4537 17663
rect 4488 17632 4537 17660
rect 4488 17620 4494 17632
rect 4525 17629 4537 17632
rect 4571 17660 4583 17663
rect 5184 17660 5212 17836
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 7190 17824 7196 17876
rect 7248 17864 7254 17876
rect 9585 17867 9643 17873
rect 9585 17864 9597 17867
rect 7248 17836 9597 17864
rect 7248 17824 7254 17836
rect 9585 17833 9597 17836
rect 9631 17833 9643 17867
rect 9585 17827 9643 17833
rect 11238 17824 11244 17876
rect 11296 17864 11302 17876
rect 12253 17867 12311 17873
rect 12253 17864 12265 17867
rect 11296 17836 12265 17864
rect 11296 17824 11302 17836
rect 12253 17833 12265 17836
rect 12299 17833 12311 17867
rect 12253 17827 12311 17833
rect 13541 17867 13599 17873
rect 13541 17833 13553 17867
rect 13587 17864 13599 17867
rect 13814 17864 13820 17876
rect 13587 17836 13820 17864
rect 13587 17833 13599 17836
rect 13541 17827 13599 17833
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 15286 17824 15292 17876
rect 15344 17864 15350 17876
rect 15749 17867 15807 17873
rect 15749 17864 15761 17867
rect 15344 17836 15761 17864
rect 15344 17824 15350 17836
rect 15749 17833 15761 17836
rect 15795 17833 15807 17867
rect 15749 17827 15807 17833
rect 17497 17867 17555 17873
rect 17497 17833 17509 17867
rect 17543 17864 17555 17867
rect 18690 17864 18696 17876
rect 17543 17836 18696 17864
rect 17543 17833 17555 17836
rect 17497 17827 17555 17833
rect 18690 17824 18696 17836
rect 18748 17824 18754 17876
rect 19613 17867 19671 17873
rect 19613 17833 19625 17867
rect 19659 17864 19671 17867
rect 19702 17864 19708 17876
rect 19659 17836 19708 17864
rect 19659 17833 19671 17836
rect 19613 17827 19671 17833
rect 19702 17824 19708 17836
rect 19760 17824 19766 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 22925 17867 22983 17873
rect 22925 17864 22937 17867
rect 20772 17836 22937 17864
rect 20772 17824 20778 17836
rect 22925 17833 22937 17836
rect 22971 17833 22983 17867
rect 22925 17827 22983 17833
rect 5936 17799 5994 17805
rect 5936 17765 5948 17799
rect 5982 17796 5994 17799
rect 5982 17768 7880 17796
rect 5982 17765 5994 17768
rect 5936 17759 5994 17765
rect 6086 17688 6092 17740
rect 6144 17728 6150 17740
rect 6181 17731 6239 17737
rect 6181 17728 6193 17731
rect 6144 17700 6193 17728
rect 6144 17688 6150 17700
rect 6181 17697 6193 17700
rect 6227 17697 6239 17731
rect 6181 17691 6239 17697
rect 6641 17731 6699 17737
rect 6641 17697 6653 17731
rect 6687 17728 6699 17731
rect 7282 17728 7288 17740
rect 6687 17700 7288 17728
rect 6687 17697 6699 17700
rect 6641 17691 6699 17697
rect 7282 17688 7288 17700
rect 7340 17688 7346 17740
rect 7852 17728 7880 17768
rect 7926 17756 7932 17808
rect 7984 17796 7990 17808
rect 8030 17799 8088 17805
rect 8030 17796 8042 17799
rect 7984 17768 8042 17796
rect 7984 17756 7990 17768
rect 8030 17765 8042 17768
rect 8076 17796 8088 17799
rect 8076 17768 9628 17796
rect 8076 17765 8088 17768
rect 8030 17759 8088 17765
rect 9493 17731 9551 17737
rect 7852 17700 8892 17728
rect 8294 17660 8300 17672
rect 4571 17632 5212 17660
rect 8255 17632 8300 17660
rect 4571 17629 4583 17632
rect 4525 17623 4583 17629
rect 8294 17620 8300 17632
rect 8352 17620 8358 17672
rect 8864 17660 8892 17700
rect 9493 17697 9505 17731
rect 9539 17697 9551 17731
rect 9600 17728 9628 17768
rect 11054 17756 11060 17808
rect 11112 17796 11118 17808
rect 11158 17799 11216 17805
rect 11158 17796 11170 17799
rect 11112 17768 11170 17796
rect 11112 17756 11118 17768
rect 11158 17765 11170 17768
rect 11204 17765 11216 17799
rect 11158 17759 11216 17765
rect 14274 17756 14280 17808
rect 14332 17796 14338 17808
rect 14614 17799 14672 17805
rect 14614 17796 14626 17799
rect 14332 17768 14626 17796
rect 14332 17756 14338 17768
rect 14614 17765 14626 17768
rect 14660 17796 14672 17799
rect 14918 17796 14924 17808
rect 14660 17768 14924 17796
rect 14660 17765 14672 17768
rect 14614 17759 14672 17765
rect 14918 17756 14924 17768
rect 14976 17756 14982 17808
rect 16574 17756 16580 17808
rect 16632 17796 16638 17808
rect 16954 17799 17012 17805
rect 16954 17796 16966 17799
rect 16632 17768 16966 17796
rect 16632 17756 16638 17768
rect 16954 17765 16966 17768
rect 17000 17765 17012 17799
rect 16954 17759 17012 17765
rect 17218 17756 17224 17808
rect 17276 17796 17282 17808
rect 19518 17796 19524 17808
rect 17276 17768 19524 17796
rect 17276 17756 17282 17768
rect 9600 17700 9720 17728
rect 9493 17691 9551 17697
rect 8864 17632 9260 17660
rect 3513 17595 3571 17601
rect 3513 17561 3525 17595
rect 3559 17592 3571 17595
rect 4062 17592 4068 17604
rect 3559 17564 4068 17592
rect 3559 17561 3571 17564
rect 3513 17555 3571 17561
rect 4062 17552 4068 17564
rect 4120 17552 4126 17604
rect 6917 17595 6975 17601
rect 6917 17561 6929 17595
rect 6963 17592 6975 17595
rect 7190 17592 7196 17604
rect 6963 17564 7196 17592
rect 6963 17561 6975 17564
rect 6917 17555 6975 17561
rect 7190 17552 7196 17564
rect 7248 17552 7254 17604
rect 9125 17595 9183 17601
rect 9125 17592 9137 17595
rect 8312 17564 9137 17592
rect 6362 17484 6368 17536
rect 6420 17524 6426 17536
rect 6457 17527 6515 17533
rect 6457 17524 6469 17527
rect 6420 17496 6469 17524
rect 6420 17484 6426 17496
rect 6457 17493 6469 17496
rect 6503 17493 6515 17527
rect 6457 17487 6515 17493
rect 7006 17484 7012 17536
rect 7064 17524 7070 17536
rect 8312 17524 8340 17564
rect 9125 17561 9137 17564
rect 9171 17561 9183 17595
rect 9232 17592 9260 17632
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 9508 17660 9536 17691
rect 9692 17669 9720 17700
rect 12066 17688 12072 17740
rect 12124 17728 12130 17740
rect 12345 17731 12403 17737
rect 12345 17728 12357 17731
rect 12124 17700 12357 17728
rect 12124 17688 12130 17700
rect 12345 17697 12357 17700
rect 12391 17697 12403 17731
rect 12345 17691 12403 17697
rect 13173 17731 13231 17737
rect 13173 17697 13185 17731
rect 13219 17728 13231 17731
rect 13354 17728 13360 17740
rect 13219 17700 13360 17728
rect 13219 17697 13231 17700
rect 13173 17691 13231 17697
rect 13354 17688 13360 17700
rect 13412 17688 13418 17740
rect 14366 17728 14372 17740
rect 14327 17700 14372 17728
rect 14366 17688 14372 17700
rect 14424 17688 14430 17740
rect 16390 17688 16396 17740
rect 16448 17728 16454 17740
rect 17313 17731 17371 17737
rect 16448 17700 17264 17728
rect 16448 17688 16454 17700
rect 9456 17632 9536 17660
rect 9677 17663 9735 17669
rect 9456 17620 9462 17632
rect 9677 17629 9689 17663
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 11425 17663 11483 17669
rect 11425 17629 11437 17663
rect 11471 17660 11483 17663
rect 11514 17660 11520 17672
rect 11471 17632 11520 17660
rect 11471 17629 11483 17632
rect 11425 17623 11483 17629
rect 11514 17620 11520 17632
rect 11572 17620 11578 17672
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17629 12219 17663
rect 12894 17660 12900 17672
rect 12855 17632 12900 17660
rect 12161 17623 12219 17629
rect 10045 17595 10103 17601
rect 10045 17592 10057 17595
rect 9232 17564 10057 17592
rect 9125 17555 9183 17561
rect 10045 17561 10057 17564
rect 10091 17592 10103 17595
rect 10410 17592 10416 17604
rect 10091 17564 10416 17592
rect 10091 17561 10103 17564
rect 10045 17555 10103 17561
rect 10410 17552 10416 17564
rect 10468 17552 10474 17604
rect 12176 17592 12204 17623
rect 12894 17620 12900 17632
rect 12952 17620 12958 17672
rect 13078 17660 13084 17672
rect 13039 17632 13084 17660
rect 13078 17620 13084 17632
rect 13136 17620 13142 17672
rect 17236 17669 17264 17700
rect 17313 17697 17325 17731
rect 17359 17728 17371 17731
rect 17402 17728 17408 17740
rect 17359 17700 17408 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 17402 17688 17408 17700
rect 17460 17688 17466 17740
rect 17604 17737 17632 17768
rect 19518 17756 19524 17768
rect 19576 17756 19582 17808
rect 21628 17799 21686 17805
rect 21628 17765 21640 17799
rect 21674 17796 21686 17799
rect 22554 17796 22560 17808
rect 21674 17768 22560 17796
rect 21674 17765 21686 17768
rect 21628 17759 21686 17765
rect 22554 17756 22560 17768
rect 22612 17756 22618 17808
rect 17589 17731 17647 17737
rect 17589 17697 17601 17731
rect 17635 17697 17647 17731
rect 17589 17691 17647 17697
rect 18316 17731 18374 17737
rect 18316 17697 18328 17731
rect 18362 17728 18374 17731
rect 19058 17728 19064 17740
rect 18362 17700 19064 17728
rect 18362 17697 18374 17700
rect 18316 17691 18374 17697
rect 19058 17688 19064 17700
rect 19116 17688 19122 17740
rect 20726 17731 20784 17737
rect 20726 17728 20738 17731
rect 19444 17700 20738 17728
rect 17221 17663 17279 17669
rect 17221 17629 17233 17663
rect 17267 17629 17279 17663
rect 17221 17623 17279 17629
rect 17678 17620 17684 17672
rect 17736 17660 17742 17672
rect 18049 17663 18107 17669
rect 18049 17660 18061 17663
rect 17736 17632 18061 17660
rect 17736 17620 17742 17632
rect 18049 17629 18061 17632
rect 18095 17629 18107 17663
rect 18049 17623 18107 17629
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 19444 17660 19472 17700
rect 20726 17697 20738 17700
rect 20772 17697 20784 17731
rect 21082 17728 21088 17740
rect 21043 17700 21088 17728
rect 20726 17691 20784 17697
rect 21082 17688 21088 17700
rect 21140 17688 21146 17740
rect 21450 17728 21456 17740
rect 21376 17700 21456 17728
rect 20990 17660 20996 17672
rect 19392 17632 19472 17660
rect 20951 17632 20996 17660
rect 19392 17620 19398 17632
rect 12176 17564 13768 17592
rect 7064 17496 8340 17524
rect 8941 17527 8999 17533
rect 7064 17484 7070 17496
rect 8941 17493 8953 17527
rect 8987 17524 8999 17527
rect 9306 17524 9312 17536
rect 8987 17496 9312 17524
rect 8987 17493 8999 17496
rect 8941 17487 8999 17493
rect 9306 17484 9312 17496
rect 9364 17484 9370 17536
rect 12713 17527 12771 17533
rect 12713 17493 12725 17527
rect 12759 17524 12771 17527
rect 13538 17524 13544 17536
rect 12759 17496 13544 17524
rect 12759 17493 12771 17496
rect 12713 17487 12771 17493
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 13740 17533 13768 17564
rect 15470 17552 15476 17604
rect 15528 17592 15534 17604
rect 19444 17601 19472 17632
rect 20990 17620 20996 17632
rect 21048 17660 21054 17672
rect 21376 17669 21404 17700
rect 21450 17688 21456 17700
rect 21508 17688 21514 17740
rect 22094 17688 22100 17740
rect 22152 17728 22158 17740
rect 23017 17731 23075 17737
rect 23017 17728 23029 17731
rect 22152 17700 23029 17728
rect 22152 17688 22158 17700
rect 23017 17697 23029 17700
rect 23063 17697 23075 17731
rect 23017 17691 23075 17697
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 21048 17632 21373 17660
rect 21048 17620 21054 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 15841 17595 15899 17601
rect 15841 17592 15853 17595
rect 15528 17564 15853 17592
rect 15528 17552 15534 17564
rect 15841 17561 15853 17564
rect 15887 17561 15899 17595
rect 15841 17555 15899 17561
rect 17773 17595 17831 17601
rect 17773 17561 17785 17595
rect 17819 17592 17831 17595
rect 19429 17595 19487 17601
rect 17819 17564 18092 17592
rect 17819 17561 17831 17564
rect 17773 17555 17831 17561
rect 13725 17527 13783 17533
rect 13725 17493 13737 17527
rect 13771 17524 13783 17527
rect 17494 17524 17500 17536
rect 13771 17496 17500 17524
rect 13771 17493 13783 17496
rect 13725 17487 13783 17493
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 17586 17484 17592 17536
rect 17644 17524 17650 17536
rect 17865 17527 17923 17533
rect 17865 17524 17877 17527
rect 17644 17496 17877 17524
rect 17644 17484 17650 17496
rect 17865 17493 17877 17496
rect 17911 17493 17923 17527
rect 18064 17524 18092 17564
rect 19429 17561 19441 17595
rect 19475 17561 19487 17595
rect 19429 17555 19487 17561
rect 22646 17552 22652 17604
rect 22704 17592 22710 17604
rect 22741 17595 22799 17601
rect 22741 17592 22753 17595
rect 22704 17564 22753 17592
rect 22704 17552 22710 17564
rect 22741 17561 22753 17564
rect 22787 17561 22799 17595
rect 22741 17555 22799 17561
rect 19334 17524 19340 17536
rect 18064 17496 19340 17524
rect 17865 17487 17923 17493
rect 19334 17484 19340 17496
rect 19392 17484 19398 17536
rect 21269 17527 21327 17533
rect 21269 17493 21281 17527
rect 21315 17524 21327 17527
rect 22554 17524 22560 17536
rect 21315 17496 22560 17524
rect 21315 17493 21327 17496
rect 21269 17487 21327 17493
rect 22554 17484 22560 17496
rect 22612 17484 22618 17536
rect 1104 17434 23460 17456
rect 1104 17382 4714 17434
rect 4766 17382 4778 17434
rect 4830 17382 4842 17434
rect 4894 17382 4906 17434
rect 4958 17382 12178 17434
rect 12230 17382 12242 17434
rect 12294 17382 12306 17434
rect 12358 17382 12370 17434
rect 12422 17382 19642 17434
rect 19694 17382 19706 17434
rect 19758 17382 19770 17434
rect 19822 17382 19834 17434
rect 19886 17382 23460 17434
rect 1104 17360 23460 17382
rect 1762 17320 1768 17332
rect 1723 17292 1768 17320
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 3237 17323 3295 17329
rect 3237 17289 3249 17323
rect 3283 17320 3295 17323
rect 3326 17320 3332 17332
rect 3283 17292 3332 17320
rect 3283 17289 3295 17292
rect 3237 17283 3295 17289
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 5810 17280 5816 17332
rect 5868 17320 5874 17332
rect 6457 17323 6515 17329
rect 6457 17320 6469 17323
rect 5868 17292 6469 17320
rect 5868 17280 5874 17292
rect 6457 17289 6469 17292
rect 6503 17289 6515 17323
rect 6457 17283 6515 17289
rect 8205 17323 8263 17329
rect 8205 17289 8217 17323
rect 8251 17320 8263 17323
rect 9582 17320 9588 17332
rect 8251 17292 9588 17320
rect 8251 17289 8263 17292
rect 8205 17283 8263 17289
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 13354 17320 13360 17332
rect 13315 17292 13360 17320
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 14918 17320 14924 17332
rect 14879 17292 14924 17320
rect 14918 17280 14924 17292
rect 14976 17280 14982 17332
rect 16577 17323 16635 17329
rect 16577 17289 16589 17323
rect 16623 17320 16635 17323
rect 17678 17320 17684 17332
rect 16623 17292 17684 17320
rect 16623 17289 16635 17292
rect 16577 17283 16635 17289
rect 17678 17280 17684 17292
rect 17736 17280 17742 17332
rect 19058 17320 19064 17332
rect 19019 17292 19064 17320
rect 19058 17280 19064 17292
rect 19116 17280 19122 17332
rect 19978 17320 19984 17332
rect 19939 17292 19984 17320
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 21082 17320 21088 17332
rect 21039 17292 21088 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 22186 17320 22192 17332
rect 21192 17292 22192 17320
rect 4614 17212 4620 17264
rect 4672 17252 4678 17264
rect 4672 17224 4844 17252
rect 4672 17212 4678 17224
rect 3234 17184 3240 17196
rect 3068 17156 3240 17184
rect 2889 17119 2947 17125
rect 2889 17085 2901 17119
rect 2935 17116 2947 17119
rect 3068 17116 3096 17156
rect 3234 17144 3240 17156
rect 3292 17144 3298 17196
rect 4816 17193 4844 17224
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 10045 17255 10103 17261
rect 10045 17252 10057 17255
rect 9732 17224 10057 17252
rect 9732 17212 9738 17224
rect 10045 17221 10057 17224
rect 10091 17221 10103 17255
rect 10045 17215 10103 17221
rect 4801 17187 4859 17193
rect 4801 17153 4813 17187
rect 4847 17153 4859 17187
rect 4801 17147 4859 17153
rect 6822 17144 6828 17196
rect 6880 17184 6886 17196
rect 7009 17187 7067 17193
rect 7009 17184 7021 17187
rect 6880 17156 7021 17184
rect 6880 17144 6886 17156
rect 7009 17153 7021 17156
rect 7055 17153 7067 17187
rect 7009 17147 7067 17153
rect 7466 17144 7472 17196
rect 7524 17184 7530 17196
rect 7653 17187 7711 17193
rect 7653 17184 7665 17187
rect 7524 17156 7665 17184
rect 7524 17144 7530 17156
rect 7653 17153 7665 17156
rect 7699 17184 7711 17187
rect 10689 17187 10747 17193
rect 7699 17156 8432 17184
rect 7699 17153 7711 17156
rect 7653 17147 7711 17153
rect 2935 17088 3096 17116
rect 3145 17119 3203 17125
rect 2935 17085 2947 17088
rect 2889 17079 2947 17085
rect 3145 17085 3157 17119
rect 3191 17085 3203 17119
rect 3145 17079 3203 17085
rect 3160 17048 3188 17079
rect 4062 17076 4068 17128
rect 4120 17116 4126 17128
rect 4350 17119 4408 17125
rect 4350 17116 4362 17119
rect 4120 17088 4362 17116
rect 4120 17076 4126 17088
rect 4350 17085 4362 17088
rect 4396 17085 4408 17119
rect 4350 17079 4408 17085
rect 4617 17119 4675 17125
rect 4617 17085 4629 17119
rect 4663 17085 4675 17119
rect 4617 17079 4675 17085
rect 5068 17119 5126 17125
rect 5068 17085 5080 17119
rect 5114 17116 5126 17119
rect 6178 17116 6184 17128
rect 5114 17088 6184 17116
rect 5114 17085 5126 17088
rect 5068 17079 5126 17085
rect 4632 17048 4660 17079
rect 6178 17076 6184 17088
rect 6236 17076 6242 17128
rect 7282 17076 7288 17128
rect 7340 17116 7346 17128
rect 8202 17116 8208 17128
rect 7340 17088 8208 17116
rect 7340 17076 7346 17088
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17085 8355 17119
rect 8404 17116 8432 17156
rect 10689 17153 10701 17187
rect 10735 17184 10747 17187
rect 11790 17184 11796 17196
rect 10735 17156 11796 17184
rect 10735 17153 10747 17156
rect 10689 17147 10747 17153
rect 11790 17144 11796 17156
rect 11848 17144 11854 17196
rect 13372 17184 13400 17280
rect 14826 17252 14832 17264
rect 14787 17224 14832 17252
rect 14826 17212 14832 17224
rect 14884 17212 14890 17264
rect 16482 17212 16488 17264
rect 16540 17252 16546 17264
rect 17405 17255 17463 17261
rect 17405 17252 17417 17255
rect 16540 17224 17417 17252
rect 16540 17212 16546 17224
rect 17405 17221 17417 17224
rect 17451 17221 17463 17255
rect 17405 17215 17463 17221
rect 13372 17156 13584 17184
rect 8553 17119 8611 17125
rect 8553 17116 8565 17119
rect 8404 17088 8565 17116
rect 8297 17079 8355 17085
rect 8553 17085 8565 17088
rect 8599 17085 8611 17119
rect 9769 17119 9827 17125
rect 9769 17116 9781 17119
rect 8553 17079 8611 17085
rect 8680 17088 9781 17116
rect 6917 17051 6975 17057
rect 6917 17048 6929 17051
rect 3160 17020 4660 17048
rect 6196 17020 6929 17048
rect 4080 16992 4108 17020
rect 6196 16992 6224 17020
rect 6917 17017 6929 17020
rect 6963 17017 6975 17051
rect 6917 17011 6975 17017
rect 7745 17051 7803 17057
rect 7745 17017 7757 17051
rect 7791 17048 7803 17051
rect 8312 17048 8340 17079
rect 8680 17060 8708 17088
rect 9769 17085 9781 17088
rect 9815 17085 9827 17119
rect 9769 17079 9827 17085
rect 10318 17076 10324 17128
rect 10376 17116 10382 17128
rect 10413 17119 10471 17125
rect 10413 17116 10425 17119
rect 10376 17088 10425 17116
rect 10376 17076 10382 17088
rect 10413 17085 10425 17088
rect 10459 17085 10471 17119
rect 10413 17079 10471 17085
rect 11241 17119 11299 17125
rect 11241 17085 11253 17119
rect 11287 17116 11299 17119
rect 11330 17116 11336 17128
rect 11287 17088 11336 17116
rect 11287 17085 11299 17088
rect 11241 17079 11299 17085
rect 7791 17020 8248 17048
rect 8312 17020 8616 17048
rect 7791 17017 7803 17020
rect 7745 17011 7803 17017
rect 4062 16940 4068 16992
rect 4120 16940 4126 16992
rect 6178 16980 6184 16992
rect 6091 16952 6184 16980
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 6822 16980 6828 16992
rect 6783 16952 6828 16980
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 7834 16940 7840 16992
rect 7892 16980 7898 16992
rect 8220 16980 8248 17020
rect 8294 16980 8300 16992
rect 7892 16952 7937 16980
rect 8220 16952 8300 16980
rect 7892 16940 7898 16952
rect 8294 16940 8300 16952
rect 8352 16940 8358 16992
rect 8588 16980 8616 17020
rect 8662 17008 8668 17060
rect 8720 17008 8726 17060
rect 11256 17048 11284 17079
rect 11330 17076 11336 17088
rect 11388 17076 11394 17128
rect 11974 17116 11980 17128
rect 11935 17088 11980 17116
rect 11974 17076 11980 17088
rect 12032 17076 12038 17128
rect 12244 17119 12302 17125
rect 12244 17085 12256 17119
rect 12290 17116 12302 17119
rect 13078 17116 13084 17128
rect 12290 17088 13084 17116
rect 12290 17085 12302 17088
rect 12244 17079 12302 17085
rect 13078 17076 13084 17088
rect 13136 17076 13142 17128
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17085 13507 17119
rect 13556 17116 13584 17156
rect 13705 17119 13763 17125
rect 13705 17116 13717 17119
rect 13556 17088 13717 17116
rect 13449 17079 13507 17085
rect 13705 17085 13717 17088
rect 13751 17085 13763 17119
rect 14844 17116 14872 17212
rect 16298 17184 16304 17196
rect 16259 17156 16304 17184
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 16034 17119 16092 17125
rect 16034 17116 16046 17119
rect 14844 17088 16046 17116
rect 13705 17079 13763 17085
rect 16034 17085 16046 17088
rect 16080 17085 16092 17119
rect 16034 17079 16092 17085
rect 16761 17119 16819 17125
rect 16761 17085 16773 17119
rect 16807 17116 16819 17119
rect 16850 17116 16856 17128
rect 16807 17088 16856 17116
rect 16807 17085 16819 17088
rect 16761 17079 16819 17085
rect 11514 17048 11520 17060
rect 9968 17020 11284 17048
rect 11427 17020 11520 17048
rect 8846 16980 8852 16992
rect 8588 16952 8852 16980
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 9677 16983 9735 16989
rect 9677 16949 9689 16983
rect 9723 16980 9735 16983
rect 9858 16980 9864 16992
rect 9723 16952 9864 16980
rect 9723 16949 9735 16952
rect 9677 16943 9735 16949
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 9968 16989 9996 17020
rect 9953 16983 10011 16989
rect 9953 16949 9965 16983
rect 9999 16949 10011 16983
rect 10502 16980 10508 16992
rect 10463 16952 10508 16980
rect 9953 16943 10011 16949
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11440 16989 11468 17020
rect 11514 17008 11520 17020
rect 11572 17048 11578 17060
rect 11992 17048 12020 17076
rect 13464 17048 13492 17079
rect 16850 17076 16856 17088
rect 16908 17076 16914 17128
rect 17313 17119 17371 17125
rect 17313 17085 17325 17119
rect 17359 17085 17371 17119
rect 17586 17116 17592 17128
rect 17547 17088 17592 17116
rect 17313 17079 17371 17085
rect 11572 17020 13492 17048
rect 17037 17051 17095 17057
rect 11572 17008 11578 17020
rect 17037 17017 17049 17051
rect 17083 17048 17095 17051
rect 17328 17048 17356 17079
rect 17586 17076 17592 17088
rect 17644 17076 17650 17128
rect 17678 17076 17684 17128
rect 17736 17125 17742 17128
rect 17736 17116 17746 17125
rect 19076 17116 19104 17280
rect 19334 17212 19340 17264
rect 19392 17252 19398 17264
rect 21192 17252 21220 17292
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 19392 17224 21220 17252
rect 22005 17255 22063 17261
rect 19392 17212 19398 17224
rect 22005 17221 22017 17255
rect 22051 17252 22063 17255
rect 22094 17252 22100 17264
rect 22051 17224 22100 17252
rect 22051 17221 22063 17224
rect 22005 17215 22063 17221
rect 22094 17212 22100 17224
rect 22152 17212 22158 17264
rect 19245 17187 19303 17193
rect 19245 17153 19257 17187
rect 19291 17184 19303 17187
rect 19610 17184 19616 17196
rect 19291 17156 19616 17184
rect 19291 17153 19303 17156
rect 19245 17147 19303 17153
rect 19610 17144 19616 17156
rect 19668 17184 19674 17196
rect 20438 17184 20444 17196
rect 19668 17156 20116 17184
rect 20399 17156 20444 17184
rect 19668 17144 19674 17156
rect 19521 17119 19579 17125
rect 19521 17116 19533 17119
rect 17736 17088 17781 17116
rect 19076 17088 19533 17116
rect 17736 17079 17746 17088
rect 19521 17085 19533 17088
rect 19567 17085 19579 17119
rect 19521 17079 19579 17085
rect 17736 17076 17742 17079
rect 17083 17020 17356 17048
rect 17083 17017 17095 17020
rect 17037 17011 17095 17017
rect 11425 16983 11483 16989
rect 11425 16980 11437 16983
rect 11204 16952 11437 16980
rect 11204 16940 11210 16952
rect 11425 16949 11437 16952
rect 11471 16949 11483 16983
rect 11425 16943 11483 16949
rect 15194 16940 15200 16992
rect 15252 16980 15258 16992
rect 16206 16980 16212 16992
rect 15252 16952 16212 16980
rect 15252 16940 15258 16952
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 17126 16980 17132 16992
rect 17087 16952 17132 16980
rect 17126 16940 17132 16952
rect 17184 16940 17190 16992
rect 17328 16980 17356 17020
rect 17770 17008 17776 17060
rect 17828 17048 17834 17060
rect 17948 17051 18006 17057
rect 17948 17048 17960 17051
rect 17828 17020 17960 17048
rect 17828 17008 17834 17020
rect 17948 17017 17960 17020
rect 17994 17048 18006 17051
rect 19429 17051 19487 17057
rect 19429 17048 19441 17051
rect 17994 17020 19441 17048
rect 17994 17017 18006 17020
rect 17948 17011 18006 17017
rect 19429 17017 19441 17020
rect 19475 17017 19487 17051
rect 20088 17048 20116 17156
rect 20438 17144 20444 17156
rect 20496 17144 20502 17196
rect 20530 17144 20536 17196
rect 20588 17184 20594 17196
rect 20588 17156 20633 17184
rect 20588 17144 20594 17156
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 21545 17187 21603 17193
rect 21545 17184 21557 17187
rect 20772 17156 21557 17184
rect 20772 17144 20778 17156
rect 21545 17153 21557 17156
rect 21591 17153 21603 17187
rect 21545 17147 21603 17153
rect 22462 17144 22468 17196
rect 22520 17184 22526 17196
rect 22649 17187 22707 17193
rect 22649 17184 22661 17187
rect 22520 17156 22661 17184
rect 22520 17144 22526 17156
rect 22649 17153 22661 17156
rect 22695 17153 22707 17187
rect 22649 17147 22707 17153
rect 22738 17144 22744 17196
rect 22796 17184 22802 17196
rect 22796 17156 22841 17184
rect 22796 17144 22802 17156
rect 20346 17116 20352 17128
rect 20307 17088 20352 17116
rect 20346 17076 20352 17088
rect 20404 17076 20410 17128
rect 20438 17048 20444 17060
rect 20088 17020 20444 17048
rect 19429 17011 19487 17017
rect 20438 17008 20444 17020
rect 20496 17048 20502 17060
rect 20548 17048 20576 17144
rect 21358 17116 21364 17128
rect 21319 17088 21364 17116
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 21818 17116 21824 17128
rect 21779 17088 21824 17116
rect 21818 17076 21824 17088
rect 21876 17076 21882 17128
rect 22554 17116 22560 17128
rect 22515 17088 22560 17116
rect 22554 17076 22560 17088
rect 22612 17076 22618 17128
rect 20496 17020 20576 17048
rect 21453 17051 21511 17057
rect 20496 17008 20502 17020
rect 21453 17017 21465 17051
rect 21499 17048 21511 17051
rect 21910 17048 21916 17060
rect 21499 17020 21916 17048
rect 21499 17017 21511 17020
rect 21453 17011 21511 17017
rect 21910 17008 21916 17020
rect 21968 17008 21974 17060
rect 19242 16980 19248 16992
rect 17328 16952 19248 16980
rect 19242 16940 19248 16952
rect 19300 16940 19306 16992
rect 19886 16980 19892 16992
rect 19847 16952 19892 16980
rect 19886 16940 19892 16952
rect 19944 16940 19950 16992
rect 22186 16980 22192 16992
rect 22147 16952 22192 16980
rect 22186 16940 22192 16952
rect 22244 16940 22250 16992
rect 1104 16890 23460 16912
rect 1104 16838 8446 16890
rect 8498 16838 8510 16890
rect 8562 16838 8574 16890
rect 8626 16838 8638 16890
rect 8690 16838 15910 16890
rect 15962 16838 15974 16890
rect 16026 16838 16038 16890
rect 16090 16838 16102 16890
rect 16154 16838 23460 16890
rect 1104 16816 23460 16838
rect 2961 16779 3019 16785
rect 2961 16745 2973 16779
rect 3007 16776 3019 16779
rect 3234 16776 3240 16788
rect 3007 16748 3240 16776
rect 3007 16745 3019 16748
rect 2961 16739 3019 16745
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 4801 16779 4859 16785
rect 4801 16745 4813 16779
rect 4847 16776 4859 16779
rect 6822 16776 6828 16788
rect 4847 16748 6828 16776
rect 4847 16745 4859 16748
rect 4801 16739 4859 16745
rect 2774 16708 2780 16720
rect 1596 16680 2780 16708
rect 1596 16649 1624 16680
rect 2774 16668 2780 16680
rect 2832 16668 2838 16720
rect 4816 16708 4844 16739
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7009 16779 7067 16785
rect 7009 16776 7021 16779
rect 6972 16748 7021 16776
rect 6972 16736 6978 16748
rect 7009 16745 7021 16748
rect 7055 16745 7067 16779
rect 7466 16776 7472 16788
rect 7427 16748 7472 16776
rect 7009 16739 7067 16745
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 7834 16736 7840 16788
rect 7892 16776 7898 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 7892 16748 9137 16776
rect 7892 16736 7898 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9125 16739 9183 16745
rect 9677 16779 9735 16785
rect 9677 16745 9689 16779
rect 9723 16745 9735 16779
rect 9677 16739 9735 16745
rect 12529 16779 12587 16785
rect 12529 16745 12541 16779
rect 12575 16776 12587 16779
rect 13078 16776 13084 16788
rect 12575 16748 13084 16776
rect 12575 16745 12587 16748
rect 12529 16739 12587 16745
rect 4356 16680 4844 16708
rect 5936 16711 5994 16717
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16609 1639 16643
rect 1581 16603 1639 16609
rect 1848 16643 1906 16649
rect 1848 16609 1860 16643
rect 1894 16640 1906 16643
rect 4356 16640 4384 16680
rect 5936 16677 5948 16711
rect 5982 16708 5994 16711
rect 6178 16708 6184 16720
rect 5982 16680 6184 16708
rect 5982 16677 5994 16680
rect 5936 16671 5994 16677
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 6457 16711 6515 16717
rect 6457 16677 6469 16711
rect 6503 16708 6515 16711
rect 6546 16708 6552 16720
rect 6503 16680 6552 16708
rect 6503 16677 6515 16680
rect 6457 16671 6515 16677
rect 6546 16668 6552 16680
rect 6604 16668 6610 16720
rect 8478 16708 8484 16720
rect 7944 16680 8484 16708
rect 1894 16612 4384 16640
rect 4433 16643 4491 16649
rect 1894 16609 1906 16612
rect 1848 16603 1906 16609
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4479 16612 4568 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4540 16572 4568 16612
rect 4614 16600 4620 16652
rect 4672 16640 4678 16652
rect 4709 16643 4767 16649
rect 4709 16640 4721 16643
rect 4672 16612 4721 16640
rect 4672 16600 4678 16612
rect 4709 16609 4721 16612
rect 4755 16609 4767 16643
rect 6362 16640 6368 16652
rect 4709 16603 4767 16609
rect 4816 16612 6368 16640
rect 4816 16572 4844 16612
rect 6362 16600 6368 16612
rect 6420 16600 6426 16652
rect 6917 16643 6975 16649
rect 6917 16609 6929 16643
rect 6963 16640 6975 16643
rect 7006 16640 7012 16652
rect 6963 16612 7012 16640
rect 6963 16609 6975 16612
rect 6917 16603 6975 16609
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 7944 16640 7972 16680
rect 8478 16668 8484 16680
rect 8536 16668 8542 16720
rect 8604 16711 8662 16717
rect 8604 16677 8616 16711
rect 8650 16708 8662 16711
rect 8938 16708 8944 16720
rect 8650 16680 8944 16708
rect 8650 16677 8662 16680
rect 8604 16671 8662 16677
rect 8938 16668 8944 16680
rect 8996 16668 9002 16720
rect 9692 16708 9720 16739
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 14458 16736 14464 16788
rect 14516 16776 14522 16788
rect 15023 16779 15081 16785
rect 15023 16776 15035 16779
rect 14516 16748 15035 16776
rect 14516 16736 14522 16748
rect 15023 16745 15035 16748
rect 15069 16745 15081 16779
rect 15023 16739 15081 16745
rect 15933 16779 15991 16785
rect 15933 16745 15945 16779
rect 15979 16776 15991 16779
rect 16206 16776 16212 16788
rect 15979 16748 16212 16776
rect 15979 16745 15991 16748
rect 15933 16739 15991 16745
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 17589 16779 17647 16785
rect 17589 16745 17601 16779
rect 17635 16776 17647 16779
rect 17770 16776 17776 16788
rect 17635 16748 17776 16776
rect 17635 16745 17647 16748
rect 17589 16739 17647 16745
rect 17770 16736 17776 16748
rect 17828 16736 17834 16788
rect 19794 16776 19800 16788
rect 17880 16748 19800 16776
rect 9766 16708 9772 16720
rect 9679 16680 9772 16708
rect 9766 16668 9772 16680
rect 9824 16708 9830 16720
rect 11394 16711 11452 16717
rect 11394 16708 11406 16711
rect 9824 16680 11406 16708
rect 9824 16668 9830 16680
rect 11394 16677 11406 16680
rect 11440 16677 11452 16711
rect 11790 16708 11796 16720
rect 11394 16671 11452 16677
rect 11532 16680 11796 16708
rect 7392 16612 7972 16640
rect 6178 16572 6184 16584
rect 4540 16544 4844 16572
rect 6139 16544 6184 16572
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 6825 16575 6883 16581
rect 6825 16541 6837 16575
rect 6871 16572 6883 16575
rect 7190 16572 7196 16584
rect 6871 16544 7196 16572
rect 6871 16541 6883 16544
rect 6825 16535 6883 16541
rect 7190 16532 7196 16544
rect 7248 16532 7254 16584
rect 7392 16513 7420 16612
rect 8018 16600 8024 16652
rect 8076 16640 8082 16652
rect 9585 16643 9643 16649
rect 9585 16640 9597 16643
rect 8076 16612 9597 16640
rect 8076 16600 8082 16612
rect 9585 16609 9597 16612
rect 9631 16609 9643 16643
rect 9585 16603 9643 16609
rect 10801 16643 10859 16649
rect 10801 16609 10813 16643
rect 10847 16640 10859 16643
rect 11532 16640 11560 16680
rect 11790 16668 11796 16680
rect 11848 16668 11854 16720
rect 13630 16708 13636 16720
rect 13591 16680 13636 16708
rect 13630 16668 13636 16680
rect 13688 16668 13694 16720
rect 14550 16708 14556 16720
rect 14511 16680 14556 16708
rect 14550 16668 14556 16680
rect 14608 16668 14614 16720
rect 16942 16668 16948 16720
rect 17000 16708 17006 16720
rect 17138 16711 17196 16717
rect 17138 16708 17150 16711
rect 17000 16680 17150 16708
rect 17000 16668 17006 16680
rect 17138 16677 17150 16680
rect 17184 16677 17196 16711
rect 17138 16671 17196 16677
rect 17494 16668 17500 16720
rect 17552 16708 17558 16720
rect 17880 16708 17908 16748
rect 19794 16736 19800 16748
rect 19852 16736 19858 16788
rect 19886 16736 19892 16788
rect 19944 16776 19950 16788
rect 20809 16779 20867 16785
rect 20809 16776 20821 16779
rect 19944 16748 20821 16776
rect 19944 16736 19950 16748
rect 20809 16745 20821 16748
rect 20855 16745 20867 16779
rect 20809 16739 20867 16745
rect 17552 16680 17908 16708
rect 17552 16668 17558 16680
rect 18046 16668 18052 16720
rect 18104 16708 18110 16720
rect 19426 16708 19432 16720
rect 18104 16680 19432 16708
rect 18104 16668 18110 16680
rect 19426 16668 19432 16680
rect 19484 16668 19490 16720
rect 21720 16711 21778 16717
rect 21720 16677 21732 16711
rect 21766 16708 21778 16711
rect 22002 16708 22008 16720
rect 21766 16680 22008 16708
rect 21766 16677 21778 16680
rect 21720 16671 21778 16677
rect 22002 16668 22008 16680
rect 22060 16668 22066 16720
rect 10847 16612 11560 16640
rect 10847 16609 10859 16612
rect 10801 16603 10859 16609
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 12989 16643 13047 16649
rect 12989 16640 13001 16643
rect 11756 16612 13001 16640
rect 11756 16600 11762 16612
rect 12989 16609 13001 16612
rect 13035 16609 13047 16643
rect 13170 16640 13176 16652
rect 13131 16612 13176 16640
rect 12989 16603 13047 16609
rect 13170 16600 13176 16612
rect 13228 16600 13234 16652
rect 15470 16640 15476 16652
rect 15431 16612 15476 16640
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 15565 16643 15623 16649
rect 15565 16609 15577 16643
rect 15611 16640 15623 16643
rect 15654 16640 15660 16652
rect 15611 16612 15660 16640
rect 15611 16609 15623 16612
rect 15565 16603 15623 16609
rect 15654 16600 15660 16612
rect 15712 16600 15718 16652
rect 16298 16600 16304 16652
rect 16356 16640 16362 16652
rect 17405 16643 17463 16649
rect 17405 16640 17417 16643
rect 16356 16612 17417 16640
rect 16356 16600 16362 16612
rect 17405 16609 17417 16612
rect 17451 16609 17463 16643
rect 17405 16603 17463 16609
rect 18713 16643 18771 16649
rect 18713 16609 18725 16643
rect 18759 16640 18771 16643
rect 18874 16640 18880 16652
rect 18759 16612 18880 16640
rect 18759 16609 18771 16612
rect 18713 16603 18771 16609
rect 18874 16600 18880 16612
rect 18932 16600 18938 16652
rect 19058 16640 19064 16652
rect 19019 16612 19064 16640
rect 19058 16600 19064 16612
rect 19116 16600 19122 16652
rect 19245 16643 19303 16649
rect 19245 16609 19257 16643
rect 19291 16640 19303 16643
rect 19978 16640 19984 16652
rect 19291 16612 19840 16640
rect 19939 16612 19984 16640
rect 19291 16609 19303 16612
rect 19245 16603 19303 16609
rect 8846 16572 8852 16584
rect 8807 16544 8852 16572
rect 8846 16532 8852 16544
rect 8904 16572 8910 16584
rect 11057 16575 11115 16581
rect 8904 16544 9674 16572
rect 8904 16532 8910 16544
rect 7377 16507 7435 16513
rect 7377 16473 7389 16507
rect 7423 16473 7435 16507
rect 7377 16467 7435 16473
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 4249 16439 4307 16445
rect 4249 16436 4261 16439
rect 4120 16408 4261 16436
rect 4120 16396 4126 16408
rect 4249 16405 4261 16408
rect 4295 16405 4307 16439
rect 4522 16436 4528 16448
rect 4483 16408 4528 16436
rect 4249 16399 4307 16405
rect 4522 16396 4528 16408
rect 4580 16396 4586 16448
rect 5442 16396 5448 16448
rect 5500 16436 5506 16448
rect 6365 16439 6423 16445
rect 6365 16436 6377 16439
rect 5500 16408 6377 16436
rect 5500 16396 5506 16408
rect 6365 16405 6377 16408
rect 6411 16405 6423 16439
rect 6365 16399 6423 16405
rect 8110 16396 8116 16448
rect 8168 16436 8174 16448
rect 9401 16439 9459 16445
rect 9401 16436 9413 16439
rect 8168 16408 9413 16436
rect 8168 16396 8174 16408
rect 9401 16405 9413 16408
rect 9447 16405 9459 16439
rect 9646 16436 9674 16544
rect 11057 16541 11069 16575
rect 11103 16572 11115 16575
rect 11146 16572 11152 16584
rect 11103 16544 11152 16572
rect 11103 16541 11115 16544
rect 11057 16535 11115 16541
rect 10778 16436 10784 16448
rect 9646 16408 10784 16436
rect 9401 16399 9459 16405
rect 10778 16396 10784 16408
rect 10836 16436 10842 16448
rect 11072 16436 11100 16535
rect 11146 16532 11152 16544
rect 11204 16532 11210 16584
rect 12894 16572 12900 16584
rect 12855 16544 12900 16572
rect 12894 16532 12900 16544
rect 12952 16532 12958 16584
rect 14458 16572 14464 16584
rect 14419 16544 14464 16572
rect 14458 16532 14464 16544
rect 14516 16532 14522 16584
rect 14642 16572 14648 16584
rect 14603 16544 14648 16572
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 15381 16575 15439 16581
rect 15381 16541 15393 16575
rect 15427 16541 15439 16575
rect 18966 16572 18972 16584
rect 18927 16544 18972 16572
rect 15381 16535 15439 16541
rect 15396 16504 15424 16535
rect 18966 16532 18972 16544
rect 19024 16532 19030 16584
rect 19426 16572 19432 16584
rect 19076 16544 19432 16572
rect 15396 16476 16068 16504
rect 16040 16445 16068 16476
rect 10836 16408 11100 16436
rect 16025 16439 16083 16445
rect 10836 16396 10842 16408
rect 16025 16405 16037 16439
rect 16071 16436 16083 16439
rect 16298 16436 16304 16448
rect 16071 16408 16304 16436
rect 16071 16405 16083 16408
rect 16025 16399 16083 16405
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 17402 16396 17408 16448
rect 17460 16436 17466 16448
rect 19076 16436 19104 16544
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 19334 16464 19340 16516
rect 19392 16504 19398 16516
rect 19613 16507 19671 16513
rect 19613 16504 19625 16507
rect 19392 16476 19625 16504
rect 19392 16464 19398 16476
rect 19613 16473 19625 16476
rect 19659 16473 19671 16507
rect 19812 16504 19840 16612
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 20073 16643 20131 16649
rect 20073 16609 20085 16643
rect 20119 16640 20131 16643
rect 20530 16640 20536 16652
rect 20119 16612 20536 16640
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 21450 16640 21456 16652
rect 21411 16612 21456 16640
rect 21450 16600 21456 16612
rect 21508 16600 21514 16652
rect 23106 16640 23112 16652
rect 23067 16612 23112 16640
rect 23106 16600 23112 16612
rect 23164 16600 23170 16652
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16572 20315 16575
rect 20714 16572 20720 16584
rect 20303 16544 20720 16572
rect 20303 16541 20315 16544
rect 20257 16535 20315 16541
rect 20714 16532 20720 16544
rect 20772 16532 20778 16584
rect 20898 16572 20904 16584
rect 20859 16544 20904 16572
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16541 21051 16575
rect 20993 16535 21051 16541
rect 20441 16507 20499 16513
rect 20441 16504 20453 16507
rect 19812 16476 20453 16504
rect 19613 16467 19671 16473
rect 20441 16473 20453 16476
rect 20487 16473 20499 16507
rect 20732 16504 20760 16532
rect 21008 16504 21036 16535
rect 20732 16476 21036 16504
rect 20441 16467 20499 16473
rect 17460 16408 19104 16436
rect 19429 16439 19487 16445
rect 17460 16396 17466 16408
rect 19429 16405 19441 16439
rect 19475 16436 19487 16439
rect 21450 16436 21456 16448
rect 19475 16408 21456 16436
rect 19475 16405 19487 16408
rect 19429 16399 19487 16405
rect 21450 16396 21456 16408
rect 21508 16396 21514 16448
rect 22830 16436 22836 16448
rect 22791 16408 22836 16436
rect 22830 16396 22836 16408
rect 22888 16396 22894 16448
rect 22922 16396 22928 16448
rect 22980 16436 22986 16448
rect 22980 16408 23025 16436
rect 22980 16396 22986 16408
rect 1104 16346 23460 16368
rect 1104 16294 4714 16346
rect 4766 16294 4778 16346
rect 4830 16294 4842 16346
rect 4894 16294 4906 16346
rect 4958 16294 12178 16346
rect 12230 16294 12242 16346
rect 12294 16294 12306 16346
rect 12358 16294 12370 16346
rect 12422 16294 19642 16346
rect 19694 16294 19706 16346
rect 19758 16294 19770 16346
rect 19822 16294 19834 16346
rect 19886 16294 23460 16346
rect 1104 16272 23460 16294
rect 3418 16232 3424 16244
rect 3379 16204 3424 16232
rect 3418 16192 3424 16204
rect 3476 16192 3482 16244
rect 6273 16235 6331 16241
rect 6273 16201 6285 16235
rect 6319 16232 6331 16235
rect 7558 16232 7564 16244
rect 6319 16204 7564 16232
rect 6319 16201 6331 16204
rect 6273 16195 6331 16201
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 8389 16235 8447 16241
rect 8389 16232 8401 16235
rect 8352 16204 8401 16232
rect 8352 16192 8358 16204
rect 8389 16201 8401 16204
rect 8435 16201 8447 16235
rect 14369 16235 14427 16241
rect 8389 16195 8447 16201
rect 9416 16204 14320 16232
rect 4614 16124 4620 16176
rect 4672 16164 4678 16176
rect 4709 16167 4767 16173
rect 4709 16164 4721 16167
rect 4672 16136 4721 16164
rect 4672 16124 4678 16136
rect 4709 16133 4721 16136
rect 4755 16133 4767 16167
rect 6914 16164 6920 16176
rect 4709 16127 4767 16133
rect 5276 16136 5764 16164
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16096 4123 16099
rect 5276 16096 5304 16136
rect 4111 16068 5304 16096
rect 5353 16099 5411 16105
rect 4111 16065 4123 16068
rect 4065 16059 4123 16065
rect 5353 16065 5365 16099
rect 5399 16096 5411 16099
rect 5442 16096 5448 16108
rect 5399 16068 5448 16096
rect 5399 16065 5411 16068
rect 5353 16059 5411 16065
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 5736 16105 5764 16136
rect 6380 16136 6920 16164
rect 5721 16099 5779 16105
rect 5721 16065 5733 16099
rect 5767 16096 5779 16099
rect 5994 16096 6000 16108
rect 5767 16068 6000 16096
rect 5767 16065 5779 16068
rect 5721 16059 5779 16065
rect 5994 16056 6000 16068
rect 6052 16056 6058 16108
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 16028 2099 16031
rect 2774 16028 2780 16040
rect 2087 16000 2780 16028
rect 2087 15997 2099 16000
rect 2041 15991 2099 15997
rect 2774 15988 2780 16000
rect 2832 15988 2838 16040
rect 4249 16031 4307 16037
rect 4249 15997 4261 16031
rect 4295 16028 4307 16031
rect 4522 16028 4528 16040
rect 4295 16000 4528 16028
rect 4295 15997 4307 16000
rect 4249 15991 4307 15997
rect 4522 15988 4528 16000
rect 4580 15988 4586 16040
rect 6380 16028 6408 16136
rect 6914 16124 6920 16136
rect 6972 16124 6978 16176
rect 6457 16099 6515 16105
rect 6457 16065 6469 16099
rect 6503 16096 6515 16099
rect 8938 16096 8944 16108
rect 6503 16068 7052 16096
rect 6503 16065 6515 16068
rect 6457 16059 6515 16065
rect 4632 16000 6408 16028
rect 1578 15960 1584 15972
rect 1539 15932 1584 15960
rect 1578 15920 1584 15932
rect 1636 15920 1642 15972
rect 1762 15920 1768 15972
rect 1820 15960 1826 15972
rect 2286 15963 2344 15969
rect 2286 15960 2298 15963
rect 1820 15932 2298 15960
rect 1820 15920 1826 15932
rect 2286 15929 2298 15932
rect 2332 15929 2344 15963
rect 2286 15923 2344 15929
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 4154 15892 4160 15904
rect 4115 15864 4160 15892
rect 4154 15852 4160 15864
rect 4212 15852 4218 15904
rect 4632 15901 4660 16000
rect 6730 15988 6736 16040
rect 6788 16028 6794 16040
rect 6917 16031 6975 16037
rect 6917 16028 6929 16031
rect 6788 16000 6929 16028
rect 6788 15988 6794 16000
rect 6917 15997 6929 16000
rect 6963 15997 6975 16031
rect 7024 16028 7052 16068
rect 8312 16068 8944 16096
rect 8018 16028 8024 16040
rect 7024 16000 8024 16028
rect 6917 15991 6975 15997
rect 8018 15988 8024 16000
rect 8076 15988 8082 16040
rect 5077 15963 5135 15969
rect 5077 15929 5089 15963
rect 5123 15960 5135 15963
rect 6362 15960 6368 15972
rect 5123 15932 6368 15960
rect 5123 15929 5135 15932
rect 5077 15923 5135 15929
rect 6362 15920 6368 15932
rect 6420 15920 6426 15972
rect 6641 15963 6699 15969
rect 6641 15929 6653 15963
rect 6687 15929 6699 15963
rect 6641 15923 6699 15929
rect 6825 15963 6883 15969
rect 6825 15929 6837 15963
rect 6871 15960 6883 15963
rect 7006 15960 7012 15972
rect 6871 15932 7012 15960
rect 6871 15929 6883 15932
rect 6825 15923 6883 15929
rect 4617 15895 4675 15901
rect 4617 15861 4629 15895
rect 4663 15861 4675 15895
rect 4617 15855 4675 15861
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 5810 15892 5816 15904
rect 5224 15864 5269 15892
rect 5771 15864 5816 15892
rect 5224 15852 5230 15864
rect 5810 15852 5816 15864
rect 5868 15852 5874 15904
rect 5902 15852 5908 15904
rect 5960 15892 5966 15904
rect 6656 15892 6684 15923
rect 7006 15920 7012 15932
rect 7064 15920 7070 15972
rect 7184 15963 7242 15969
rect 7184 15929 7196 15963
rect 7230 15960 7242 15963
rect 8202 15960 8208 15972
rect 7230 15932 8208 15960
rect 7230 15929 7242 15932
rect 7184 15923 7242 15929
rect 7199 15892 7227 15923
rect 8202 15920 8208 15932
rect 8260 15920 8266 15972
rect 8312 15901 8340 16068
rect 8938 16056 8944 16068
rect 8996 16056 9002 16108
rect 9122 16056 9128 16108
rect 9180 16096 9186 16108
rect 9416 16105 9444 16204
rect 12176 16176 12204 16204
rect 14292 16176 14320 16204
rect 14369 16201 14381 16235
rect 14415 16232 14427 16235
rect 14550 16232 14556 16244
rect 14415 16204 14556 16232
rect 14415 16201 14427 16204
rect 14369 16195 14427 16201
rect 14550 16192 14556 16204
rect 14608 16192 14614 16244
rect 16761 16235 16819 16241
rect 16761 16201 16773 16235
rect 16807 16232 16819 16235
rect 17310 16232 17316 16244
rect 16807 16204 17316 16232
rect 16807 16201 16819 16204
rect 16761 16195 16819 16201
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 18874 16192 18880 16244
rect 18932 16232 18938 16244
rect 18969 16235 19027 16241
rect 18969 16232 18981 16235
rect 18932 16204 18981 16232
rect 18932 16192 18938 16204
rect 18969 16201 18981 16204
rect 19015 16232 19027 16235
rect 19015 16204 19754 16232
rect 19015 16201 19027 16204
rect 18969 16195 19027 16201
rect 12158 16124 12164 16176
rect 12216 16124 12222 16176
rect 14274 16164 14280 16176
rect 14187 16136 14280 16164
rect 14274 16124 14280 16136
rect 14332 16164 14338 16176
rect 19610 16164 19616 16176
rect 14332 16136 14964 16164
rect 14332 16124 14338 16136
rect 9401 16099 9459 16105
rect 9401 16096 9413 16099
rect 9180 16068 9413 16096
rect 9180 16056 9186 16068
rect 9401 16065 9413 16068
rect 9447 16065 9459 16099
rect 9401 16059 9459 16065
rect 9858 16056 9864 16108
rect 9916 16096 9922 16108
rect 10137 16099 10195 16105
rect 9916 16068 9961 16096
rect 9916 16056 9922 16068
rect 10137 16065 10149 16099
rect 10183 16096 10195 16099
rect 10318 16096 10324 16108
rect 10183 16068 10324 16096
rect 10183 16065 10195 16068
rect 10137 16059 10195 16065
rect 10318 16056 10324 16068
rect 10376 16056 10382 16108
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16096 11943 16099
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 11931 16068 12296 16096
rect 11931 16065 11943 16068
rect 11885 16059 11943 16065
rect 11974 15988 11980 16040
rect 12032 16028 12038 16040
rect 12161 16031 12219 16037
rect 12161 16028 12173 16031
rect 12032 16000 12173 16028
rect 12032 15988 12038 16000
rect 12161 15997 12173 16000
rect 12207 15997 12219 16031
rect 12268 16028 12296 16068
rect 13556 16068 13737 16096
rect 12894 16028 12900 16040
rect 12268 16000 12900 16028
rect 12161 15991 12219 15997
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 12428 15963 12486 15969
rect 11072 15932 12112 15960
rect 5960 15864 6005 15892
rect 6656 15864 7227 15892
rect 8297 15895 8355 15901
rect 5960 15852 5966 15864
rect 8297 15861 8309 15895
rect 8343 15861 8355 15895
rect 8754 15892 8760 15904
rect 8715 15864 8760 15892
rect 8297 15855 8355 15861
rect 8754 15852 8760 15864
rect 8812 15852 8818 15904
rect 8846 15852 8852 15904
rect 8904 15892 8910 15904
rect 9306 15892 9312 15904
rect 8904 15864 8949 15892
rect 9219 15864 9312 15892
rect 8904 15852 8910 15864
rect 9306 15852 9312 15864
rect 9364 15892 9370 15904
rect 9867 15895 9925 15901
rect 9867 15892 9879 15895
rect 9364 15864 9879 15892
rect 9364 15852 9370 15864
rect 9867 15861 9879 15864
rect 9913 15892 9925 15895
rect 11072 15892 11100 15932
rect 11238 15892 11244 15904
rect 9913 15864 11100 15892
rect 11199 15864 11244 15892
rect 9913 15861 9925 15864
rect 9867 15855 9925 15861
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 11330 15852 11336 15904
rect 11388 15892 11394 15904
rect 12084 15901 12112 15932
rect 12428 15929 12440 15963
rect 12474 15960 12486 15963
rect 12618 15960 12624 15972
rect 12474 15932 12624 15960
rect 12474 15929 12486 15932
rect 12428 15923 12486 15929
rect 12618 15920 12624 15932
rect 12676 15960 12682 15972
rect 13170 15960 13176 15972
rect 12676 15932 13176 15960
rect 12676 15920 12682 15932
rect 13170 15920 13176 15932
rect 13228 15920 13234 15972
rect 12069 15895 12127 15901
rect 11388 15864 11433 15892
rect 11388 15852 11394 15864
rect 12069 15861 12081 15895
rect 12115 15892 12127 15895
rect 12710 15892 12716 15904
rect 12115 15864 12716 15892
rect 12115 15861 12127 15864
rect 12069 15855 12127 15861
rect 12710 15852 12716 15864
rect 12768 15852 12774 15904
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13556 15901 13584 16068
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 14642 16096 14648 16108
rect 14603 16068 14648 16096
rect 13725 16059 13783 16065
rect 14642 16056 14648 16068
rect 14700 16056 14706 16108
rect 14936 16105 14964 16136
rect 18616 16136 19616 16164
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15427 16099 15485 16105
rect 15427 16065 15439 16099
rect 15473 16096 15485 16099
rect 15746 16096 15752 16108
rect 15473 16068 15752 16096
rect 15473 16065 15485 16068
rect 15427 16059 15485 16065
rect 15746 16056 15752 16068
rect 15804 16056 15810 16108
rect 15654 16028 15660 16040
rect 15028 16000 15660 16028
rect 13909 15963 13967 15969
rect 13909 15929 13921 15963
rect 13955 15960 13967 15963
rect 14090 15960 14096 15972
rect 13955 15932 14096 15960
rect 13955 15929 13967 15932
rect 13909 15923 13967 15929
rect 14090 15920 14096 15932
rect 14148 15960 14154 15972
rect 15028 15960 15056 16000
rect 15654 15988 15660 16000
rect 15712 15988 15718 16040
rect 16945 16031 17003 16037
rect 16945 15997 16957 16031
rect 16991 16028 17003 16031
rect 17126 16028 17132 16040
rect 16991 16000 17132 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17126 15988 17132 16000
rect 17184 15988 17190 16040
rect 17494 16028 17500 16040
rect 17455 16000 17500 16028
rect 17494 15988 17500 16000
rect 17552 15988 17558 16040
rect 17586 15988 17592 16040
rect 17644 16028 17650 16040
rect 17862 16037 17868 16040
rect 17856 16028 17868 16037
rect 17644 16000 17689 16028
rect 17775 16000 17868 16028
rect 17644 15988 17650 16000
rect 17856 15991 17868 16000
rect 17920 16028 17926 16040
rect 18616 16028 18644 16136
rect 19610 16124 19616 16136
rect 19668 16124 19674 16176
rect 19518 16096 19524 16108
rect 19479 16068 19524 16096
rect 19518 16056 19524 16068
rect 19576 16056 19582 16108
rect 19726 16096 19754 16204
rect 19978 16192 19984 16244
rect 20036 16232 20042 16244
rect 20165 16235 20223 16241
rect 20165 16232 20177 16235
rect 20036 16204 20177 16232
rect 20036 16192 20042 16204
rect 20165 16201 20177 16204
rect 20211 16201 20223 16235
rect 20165 16195 20223 16201
rect 20898 16192 20904 16244
rect 20956 16232 20962 16244
rect 20993 16235 21051 16241
rect 20993 16232 21005 16235
rect 20956 16204 21005 16232
rect 20956 16192 20962 16204
rect 20993 16201 21005 16204
rect 21039 16201 21051 16235
rect 21818 16232 21824 16244
rect 21779 16204 21824 16232
rect 20993 16195 21051 16201
rect 21818 16192 21824 16204
rect 21876 16232 21882 16244
rect 22925 16235 22983 16241
rect 21876 16204 22094 16232
rect 21876 16192 21882 16204
rect 19794 16124 19800 16176
rect 19852 16164 19858 16176
rect 22066 16164 22094 16204
rect 22925 16201 22937 16235
rect 22971 16232 22983 16235
rect 23106 16232 23112 16244
rect 22971 16204 23112 16232
rect 22971 16201 22983 16204
rect 22925 16195 22983 16201
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 19852 16136 20576 16164
rect 22066 16136 22508 16164
rect 19852 16124 19858 16136
rect 20070 16096 20076 16108
rect 19726 16068 20076 16096
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 20438 16096 20444 16108
rect 20399 16068 20444 16096
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20548 16105 20576 16136
rect 20533 16099 20591 16105
rect 20533 16065 20545 16099
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16096 21327 16099
rect 22370 16096 22376 16108
rect 21315 16068 22094 16096
rect 22331 16068 22376 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 17920 16000 18644 16028
rect 19153 16031 19211 16037
rect 17862 15988 17868 15991
rect 17920 15988 17926 16000
rect 19153 15997 19165 16031
rect 19199 16028 19211 16031
rect 19334 16028 19340 16040
rect 19199 16000 19340 16028
rect 19199 15997 19211 16000
rect 19153 15991 19211 15997
rect 19334 15988 19340 16000
rect 19392 15988 19398 16040
rect 19705 16031 19763 16037
rect 19705 15997 19717 16031
rect 19751 16028 19763 16031
rect 20714 16028 20720 16040
rect 19751 16000 20720 16028
rect 19751 15997 19763 16000
rect 19705 15991 19763 15997
rect 20714 15988 20720 16000
rect 20772 15988 20778 16040
rect 21450 16028 21456 16040
rect 21411 16000 21456 16028
rect 21450 15988 21456 16000
rect 21508 15988 21514 16040
rect 18506 15960 18512 15972
rect 14148 15932 15056 15960
rect 17144 15932 18512 15960
rect 14148 15920 14154 15932
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 13412 15864 13553 15892
rect 13412 15852 13418 15864
rect 13541 15861 13553 15864
rect 13587 15861 13599 15895
rect 13541 15855 13599 15861
rect 13722 15852 13728 15904
rect 13780 15892 13786 15904
rect 14001 15895 14059 15901
rect 14001 15892 14013 15895
rect 13780 15864 14013 15892
rect 13780 15852 13786 15864
rect 14001 15861 14013 15864
rect 14047 15861 14059 15895
rect 14001 15855 14059 15861
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14829 15895 14887 15901
rect 14829 15892 14841 15895
rect 14240 15864 14841 15892
rect 14240 15852 14246 15864
rect 14829 15861 14841 15864
rect 14875 15892 14887 15895
rect 15378 15892 15384 15904
rect 15436 15901 15442 15904
rect 17144 15901 17172 15932
rect 18506 15920 18512 15932
rect 18564 15920 18570 15972
rect 21361 15963 21419 15969
rect 21361 15960 21373 15963
rect 19352 15932 21373 15960
rect 14875 15864 15384 15892
rect 14875 15861 14887 15864
rect 14829 15855 14887 15861
rect 15378 15852 15384 15864
rect 15436 15892 15445 15901
rect 17129 15895 17187 15901
rect 15436 15864 15481 15892
rect 15436 15855 15445 15864
rect 17129 15861 17141 15895
rect 17175 15861 17187 15895
rect 17129 15855 17187 15861
rect 15436 15852 15442 15855
rect 17218 15852 17224 15904
rect 17276 15892 17282 15904
rect 17313 15895 17371 15901
rect 17313 15892 17325 15895
rect 17276 15864 17325 15892
rect 17276 15852 17282 15864
rect 17313 15861 17325 15864
rect 17359 15861 17371 15895
rect 17313 15855 17371 15861
rect 17586 15852 17592 15904
rect 17644 15892 17650 15904
rect 18874 15892 18880 15904
rect 17644 15864 18880 15892
rect 17644 15852 17650 15864
rect 18874 15852 18880 15864
rect 18932 15852 18938 15904
rect 19352 15901 19380 15932
rect 21361 15929 21373 15932
rect 21407 15929 21419 15963
rect 22066 15960 22094 16068
rect 22370 16056 22376 16068
rect 22428 16056 22434 16108
rect 22480 16105 22508 16136
rect 22465 16099 22523 16105
rect 22465 16065 22477 16099
rect 22511 16065 22523 16099
rect 22465 16059 22523 16065
rect 22186 15988 22192 16040
rect 22244 16028 22250 16040
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 22244 16000 22569 16028
rect 22244 15988 22250 16000
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 22738 15960 22744 15972
rect 22066 15932 22744 15960
rect 21361 15923 21419 15929
rect 22738 15920 22744 15932
rect 22796 15920 22802 15972
rect 19337 15895 19395 15901
rect 19337 15861 19349 15895
rect 19383 15861 19395 15895
rect 19337 15855 19395 15861
rect 19794 15852 19800 15904
rect 19852 15892 19858 15904
rect 19852 15864 19897 15892
rect 19852 15852 19858 15864
rect 20070 15852 20076 15904
rect 20128 15892 20134 15904
rect 20625 15895 20683 15901
rect 20625 15892 20637 15895
rect 20128 15864 20637 15892
rect 20128 15852 20134 15864
rect 20625 15861 20637 15864
rect 20671 15861 20683 15895
rect 20625 15855 20683 15861
rect 1104 15802 23460 15824
rect 1104 15750 8446 15802
rect 8498 15750 8510 15802
rect 8562 15750 8574 15802
rect 8626 15750 8638 15802
rect 8690 15750 15910 15802
rect 15962 15750 15974 15802
rect 16026 15750 16038 15802
rect 16090 15750 16102 15802
rect 16154 15750 23460 15802
rect 1104 15728 23460 15750
rect 2774 15688 2780 15700
rect 2746 15648 2780 15688
rect 2832 15688 2838 15700
rect 3510 15688 3516 15700
rect 2832 15660 3516 15688
rect 2832 15648 2838 15660
rect 3510 15648 3516 15660
rect 3568 15688 3574 15700
rect 4062 15688 4068 15700
rect 3568 15660 4068 15688
rect 3568 15648 3574 15660
rect 4062 15648 4068 15660
rect 4120 15688 4126 15700
rect 6733 15691 6791 15697
rect 4120 15660 5580 15688
rect 4120 15648 4126 15660
rect 2746 15620 2774 15648
rect 5442 15620 5448 15632
rect 1504 15592 2774 15620
rect 3252 15592 5448 15620
rect 1504 15561 1532 15592
rect 1762 15561 1768 15564
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15521 1547 15555
rect 1756 15552 1768 15561
rect 1723 15524 1768 15552
rect 1489 15515 1547 15521
rect 1756 15515 1768 15524
rect 1762 15512 1768 15515
rect 1820 15512 1826 15564
rect 3252 15552 3280 15592
rect 5442 15580 5448 15592
rect 5500 15580 5506 15632
rect 5552 15620 5580 15660
rect 6733 15657 6745 15691
rect 6779 15657 6791 15691
rect 8202 15688 8208 15700
rect 8163 15660 8208 15688
rect 6733 15651 6791 15657
rect 6748 15620 6776 15651
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 8754 15688 8760 15700
rect 8527 15660 8760 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 8754 15648 8760 15660
rect 8812 15648 8818 15700
rect 9401 15691 9459 15697
rect 9401 15657 9413 15691
rect 9447 15688 9459 15691
rect 9674 15688 9680 15700
rect 9447 15660 9680 15688
rect 9447 15657 9459 15660
rect 9401 15651 9459 15657
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 9858 15688 9864 15700
rect 9819 15660 9864 15688
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 10100 15660 10333 15688
rect 10100 15648 10106 15660
rect 10321 15657 10333 15660
rect 10367 15688 10379 15691
rect 10502 15688 10508 15700
rect 10367 15660 10508 15688
rect 10367 15657 10379 15660
rect 10321 15651 10379 15657
rect 10502 15648 10508 15660
rect 10560 15648 10566 15700
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 11238 15688 11244 15700
rect 10652 15660 11244 15688
rect 10652 15648 10658 15660
rect 11238 15648 11244 15660
rect 11296 15688 11302 15700
rect 12161 15691 12219 15697
rect 11296 15660 11652 15688
rect 11296 15648 11302 15660
rect 6822 15620 6828 15632
rect 5552 15592 6132 15620
rect 6735 15592 6828 15620
rect 3068 15524 3280 15552
rect 3329 15555 3387 15561
rect 3068 15493 3096 15524
rect 3329 15521 3341 15555
rect 3375 15552 3387 15555
rect 3694 15552 3700 15564
rect 3375 15524 3700 15552
rect 3375 15521 3387 15524
rect 3329 15515 3387 15521
rect 3694 15512 3700 15524
rect 3752 15512 3758 15564
rect 3881 15555 3939 15561
rect 3881 15521 3893 15555
rect 3927 15552 3939 15555
rect 3970 15552 3976 15564
rect 3927 15524 3976 15552
rect 3927 15521 3939 15524
rect 3881 15515 3939 15521
rect 3970 15512 3976 15524
rect 4028 15512 4034 15564
rect 4148 15555 4206 15561
rect 4148 15521 4160 15555
rect 4194 15552 4206 15555
rect 4522 15552 4528 15564
rect 4194 15524 4528 15552
rect 4194 15521 4206 15524
rect 4148 15515 4206 15521
rect 4522 15512 4528 15524
rect 4580 15512 4586 15564
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15552 5411 15555
rect 5552 15552 5580 15592
rect 5399 15524 5580 15552
rect 5620 15555 5678 15561
rect 5399 15521 5411 15524
rect 5353 15515 5411 15521
rect 5620 15521 5632 15555
rect 5666 15552 5678 15555
rect 5994 15552 6000 15564
rect 5666 15524 6000 15552
rect 5666 15521 5678 15524
rect 5620 15515 5678 15521
rect 5994 15512 6000 15524
rect 6052 15512 6058 15564
rect 6104 15552 6132 15592
rect 6822 15580 6828 15592
rect 6880 15620 6886 15632
rect 7070 15623 7128 15629
rect 7070 15620 7082 15623
rect 6880 15592 7082 15620
rect 6880 15580 6886 15592
rect 7070 15589 7082 15592
rect 7116 15589 7128 15623
rect 7070 15583 7128 15589
rect 9493 15623 9551 15629
rect 9493 15589 9505 15623
rect 9539 15620 9551 15623
rect 11330 15620 11336 15632
rect 9539 15592 11336 15620
rect 9539 15589 9551 15592
rect 9493 15583 9551 15589
rect 11330 15580 11336 15592
rect 11388 15580 11394 15632
rect 6104 15524 6776 15552
rect 6748 15496 6776 15524
rect 7558 15512 7564 15564
rect 7616 15552 7622 15564
rect 8297 15555 8355 15561
rect 8297 15552 8309 15555
rect 7616 15524 8309 15552
rect 7616 15512 7622 15524
rect 8297 15521 8309 15524
rect 8343 15521 8355 15555
rect 8297 15515 8355 15521
rect 8573 15555 8631 15561
rect 8573 15521 8585 15555
rect 8619 15521 8631 15555
rect 11048 15555 11106 15561
rect 11048 15552 11060 15555
rect 8573 15515 8631 15521
rect 10152 15524 11060 15552
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15453 3111 15487
rect 3234 15484 3240 15496
rect 3195 15456 3240 15484
rect 3053 15447 3111 15453
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 6825 15487 6883 15493
rect 6825 15484 6837 15487
rect 6788 15456 6837 15484
rect 6788 15444 6794 15456
rect 6825 15453 6837 15456
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 7926 15444 7932 15496
rect 7984 15484 7990 15496
rect 8588 15484 8616 15515
rect 7984 15456 8616 15484
rect 9309 15487 9367 15493
rect 7984 15444 7990 15456
rect 9309 15453 9321 15487
rect 9355 15484 9367 15487
rect 9766 15484 9772 15496
rect 9355 15456 9772 15484
rect 9355 15453 9367 15456
rect 9309 15447 9367 15453
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 10152 15493 10180 15524
rect 11048 15521 11060 15524
rect 11094 15552 11106 15555
rect 11514 15552 11520 15564
rect 11094 15524 11520 15552
rect 11094 15521 11106 15524
rect 11048 15515 11106 15521
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 11624 15552 11652 15660
rect 12161 15657 12173 15691
rect 12207 15688 12219 15691
rect 12618 15688 12624 15700
rect 12207 15660 12624 15688
rect 12207 15657 12219 15660
rect 12161 15651 12219 15657
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 12710 15648 12716 15700
rect 12768 15697 12774 15700
rect 12768 15688 12777 15697
rect 14090 15688 14096 15700
rect 12768 15660 13983 15688
rect 14051 15660 14096 15688
rect 12768 15651 12777 15660
rect 12768 15648 12774 15651
rect 13955 15620 13983 15660
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 15654 15648 15660 15700
rect 15712 15688 15718 15700
rect 15841 15691 15899 15697
rect 15841 15688 15853 15691
rect 15712 15660 15853 15688
rect 15712 15648 15718 15660
rect 15841 15657 15853 15660
rect 15887 15657 15899 15691
rect 15841 15651 15899 15657
rect 17497 15691 17555 15697
rect 17497 15657 17509 15691
rect 17543 15688 17555 15691
rect 17862 15688 17868 15700
rect 17543 15660 17868 15688
rect 17543 15657 17555 15660
rect 17497 15651 17555 15657
rect 14182 15620 14188 15632
rect 13955 15592 14188 15620
rect 14182 15580 14188 15592
rect 14240 15580 14246 15632
rect 14458 15580 14464 15632
rect 14516 15620 14522 15632
rect 15482 15623 15540 15629
rect 15482 15620 15494 15623
rect 14516 15592 15494 15620
rect 14516 15580 14522 15592
rect 15482 15589 15494 15592
rect 15528 15589 15540 15623
rect 15856 15620 15884 15651
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 18966 15648 18972 15700
rect 19024 15688 19030 15700
rect 19613 15691 19671 15697
rect 19024 15660 19069 15688
rect 19024 15648 19030 15660
rect 19613 15657 19625 15691
rect 19659 15688 19671 15691
rect 19794 15688 19800 15700
rect 19659 15660 19800 15688
rect 19659 15657 19671 15660
rect 19613 15651 19671 15657
rect 16114 15620 16120 15632
rect 15856 15592 16120 15620
rect 15482 15583 15540 15589
rect 16114 15580 16120 15592
rect 16172 15580 16178 15632
rect 16298 15580 16304 15632
rect 16356 15620 16362 15632
rect 16954 15623 17012 15629
rect 16954 15620 16966 15623
rect 16356 15592 16966 15620
rect 16356 15580 16362 15592
rect 16954 15589 16966 15592
rect 17000 15589 17012 15623
rect 16954 15583 17012 15589
rect 18632 15623 18690 15629
rect 18632 15589 18644 15623
rect 18678 15620 18690 15623
rect 19628 15620 19656 15651
rect 19794 15648 19800 15660
rect 19852 15648 19858 15700
rect 22738 15688 22744 15700
rect 22699 15660 22744 15688
rect 22738 15648 22744 15660
rect 22796 15648 22802 15700
rect 18678 15592 19656 15620
rect 18678 15589 18690 15592
rect 18632 15583 18690 15589
rect 20254 15580 20260 15632
rect 20312 15620 20318 15632
rect 20530 15620 20536 15632
rect 20312 15592 20536 15620
rect 20312 15580 20318 15592
rect 20530 15580 20536 15592
rect 20588 15580 20594 15632
rect 20714 15580 20720 15632
rect 20772 15629 20778 15632
rect 20772 15620 20784 15629
rect 21536 15623 21594 15629
rect 20772 15592 20817 15620
rect 20772 15583 20784 15592
rect 21536 15589 21548 15623
rect 21582 15620 21594 15623
rect 22278 15620 22284 15632
rect 21582 15592 22284 15620
rect 21582 15589 21594 15592
rect 21536 15583 21594 15589
rect 20772 15580 20778 15583
rect 22278 15580 22284 15592
rect 22336 15620 22342 15632
rect 22830 15620 22836 15632
rect 22336 15592 22836 15620
rect 22336 15580 22342 15592
rect 22830 15580 22836 15592
rect 22888 15580 22894 15632
rect 12989 15555 13047 15561
rect 12989 15552 13001 15555
rect 11624 15524 13001 15552
rect 12989 15521 13001 15524
rect 13035 15521 13047 15555
rect 12989 15515 13047 15521
rect 15749 15555 15807 15561
rect 15749 15521 15761 15555
rect 15795 15552 15807 15555
rect 16390 15552 16396 15564
rect 15795 15524 16396 15552
rect 15795 15521 15807 15524
rect 15749 15515 15807 15521
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 17405 15555 17463 15561
rect 17405 15521 17417 15555
rect 17451 15552 17463 15555
rect 17494 15552 17500 15564
rect 17451 15524 17500 15552
rect 17451 15521 17463 15524
rect 17405 15515 17463 15521
rect 17494 15512 17500 15524
rect 17552 15552 17558 15564
rect 17552 15524 19012 15552
rect 17552 15512 17558 15524
rect 10137 15487 10195 15493
rect 10137 15453 10149 15487
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15484 10287 15487
rect 10594 15484 10600 15496
rect 10275 15456 10600 15484
rect 10275 15453 10287 15456
rect 10229 15447 10287 15453
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 10778 15484 10784 15496
rect 10739 15456 10784 15484
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 12158 15444 12164 15496
rect 12216 15484 12222 15496
rect 12253 15487 12311 15493
rect 12253 15484 12265 15487
rect 12216 15456 12265 15484
rect 12216 15444 12222 15456
rect 12253 15453 12265 15456
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 12710 15444 12716 15496
rect 12768 15484 12774 15496
rect 13722 15484 13728 15496
rect 12768 15456 13728 15484
rect 12768 15444 12774 15456
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 17221 15487 17279 15493
rect 17221 15453 17233 15487
rect 17267 15484 17279 15487
rect 17586 15484 17592 15496
rect 17267 15456 17592 15484
rect 17267 15453 17279 15456
rect 17221 15447 17279 15453
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 18874 15484 18880 15496
rect 18835 15456 18880 15484
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 18984 15484 19012 15524
rect 19058 15512 19064 15564
rect 19116 15552 19122 15564
rect 19153 15555 19211 15561
rect 19153 15552 19165 15555
rect 19116 15524 19165 15552
rect 19116 15512 19122 15524
rect 19153 15521 19165 15524
rect 19199 15521 19211 15555
rect 19153 15515 19211 15521
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15521 19487 15555
rect 19429 15515 19487 15521
rect 19334 15484 19340 15496
rect 18984 15456 19340 15484
rect 19334 15444 19340 15456
rect 19392 15444 19398 15496
rect 8757 15419 8815 15425
rect 8757 15385 8769 15419
rect 8803 15416 8815 15419
rect 9214 15416 9220 15428
rect 8803 15388 9220 15416
rect 8803 15385 8815 15388
rect 8757 15379 8815 15385
rect 9214 15376 9220 15388
rect 9272 15376 9278 15428
rect 10796 15416 10824 15444
rect 14369 15419 14427 15425
rect 14369 15416 14381 15419
rect 10244 15388 10824 15416
rect 13648 15388 14381 15416
rect 2866 15348 2872 15360
rect 2827 15320 2872 15348
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 3697 15351 3755 15357
rect 3697 15317 3709 15351
rect 3743 15348 3755 15351
rect 3878 15348 3884 15360
rect 3743 15320 3884 15348
rect 3743 15317 3755 15320
rect 3697 15311 3755 15317
rect 3878 15308 3884 15320
rect 3936 15308 3942 15360
rect 5258 15348 5264 15360
rect 5219 15320 5264 15348
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 10134 15308 10140 15360
rect 10192 15348 10198 15360
rect 10244 15348 10272 15388
rect 10192 15320 10272 15348
rect 10689 15351 10747 15357
rect 10192 15308 10198 15320
rect 10689 15317 10701 15351
rect 10735 15348 10747 15351
rect 11698 15348 11704 15360
rect 10735 15320 11704 15348
rect 10735 15317 10747 15320
rect 10689 15311 10747 15317
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 11790 15308 11796 15360
rect 11848 15348 11854 15360
rect 13648 15348 13676 15388
rect 14369 15385 14381 15388
rect 14415 15385 14427 15419
rect 14369 15379 14427 15385
rect 11848 15320 13676 15348
rect 11848 15308 11854 15320
rect 18874 15308 18880 15360
rect 18932 15348 18938 15360
rect 19245 15351 19303 15357
rect 19245 15348 19257 15351
rect 18932 15320 19257 15348
rect 18932 15308 18938 15320
rect 19245 15317 19257 15320
rect 19291 15317 19303 15351
rect 19444 15348 19472 15515
rect 19978 15512 19984 15564
rect 20036 15552 20042 15564
rect 20993 15555 21051 15561
rect 20993 15552 21005 15555
rect 20036 15524 21005 15552
rect 20036 15512 20042 15524
rect 20993 15521 21005 15524
rect 21039 15521 21051 15555
rect 20993 15515 21051 15521
rect 21008 15484 21036 15515
rect 21174 15512 21180 15564
rect 21232 15552 21238 15564
rect 22925 15555 22983 15561
rect 22925 15552 22937 15555
rect 21232 15524 22937 15552
rect 21232 15512 21238 15524
rect 22925 15521 22937 15524
rect 22971 15521 22983 15555
rect 22925 15515 22983 15521
rect 21269 15487 21327 15493
rect 21269 15484 21281 15487
rect 21008 15456 21281 15484
rect 21269 15453 21281 15456
rect 21315 15453 21327 15487
rect 21269 15447 21327 15453
rect 20622 15348 20628 15360
rect 19444 15320 20628 15348
rect 19245 15311 19303 15317
rect 20622 15308 20628 15320
rect 20680 15348 20686 15360
rect 21085 15351 21143 15357
rect 21085 15348 21097 15351
rect 20680 15320 21097 15348
rect 20680 15308 20686 15320
rect 21085 15317 21097 15320
rect 21131 15317 21143 15351
rect 21284 15348 21312 15447
rect 21450 15348 21456 15360
rect 21284 15320 21456 15348
rect 21085 15311 21143 15317
rect 21450 15308 21456 15320
rect 21508 15308 21514 15360
rect 22554 15308 22560 15360
rect 22612 15348 22618 15360
rect 22649 15351 22707 15357
rect 22649 15348 22661 15351
rect 22612 15320 22661 15348
rect 22612 15308 22618 15320
rect 22649 15317 22661 15320
rect 22695 15317 22707 15351
rect 22649 15311 22707 15317
rect 1104 15258 23460 15280
rect 1104 15206 4714 15258
rect 4766 15206 4778 15258
rect 4830 15206 4842 15258
rect 4894 15206 4906 15258
rect 4958 15206 12178 15258
rect 12230 15206 12242 15258
rect 12294 15206 12306 15258
rect 12358 15206 12370 15258
rect 12422 15206 19642 15258
rect 19694 15206 19706 15258
rect 19758 15206 19770 15258
rect 19822 15206 19834 15258
rect 19886 15206 23460 15258
rect 1104 15184 23460 15206
rect 4522 15104 4528 15156
rect 4580 15144 4586 15156
rect 4893 15147 4951 15153
rect 4893 15144 4905 15147
rect 4580 15116 4905 15144
rect 4580 15104 4586 15116
rect 4893 15113 4905 15116
rect 4939 15113 4951 15147
rect 4893 15107 4951 15113
rect 4985 15147 5043 15153
rect 4985 15113 4997 15147
rect 5031 15144 5043 15147
rect 5166 15144 5172 15156
rect 5031 15116 5172 15144
rect 5031 15113 5043 15116
rect 4985 15107 5043 15113
rect 3510 15008 3516 15020
rect 3471 14980 3516 15008
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 4908 15008 4936 15107
rect 5166 15104 5172 15116
rect 5224 15104 5230 15156
rect 6362 15104 6368 15156
rect 6420 15144 6426 15156
rect 6457 15147 6515 15153
rect 6457 15144 6469 15147
rect 6420 15116 6469 15144
rect 6420 15104 6426 15116
rect 6457 15113 6469 15116
rect 6503 15113 6515 15147
rect 6457 15107 6515 15113
rect 8297 15147 8355 15153
rect 8297 15113 8309 15147
rect 8343 15144 8355 15147
rect 8846 15144 8852 15156
rect 8343 15116 8852 15144
rect 8343 15113 8355 15116
rect 8297 15107 8355 15113
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 9217 15147 9275 15153
rect 9217 15113 9229 15147
rect 9263 15144 9275 15147
rect 9858 15144 9864 15156
rect 9263 15116 9864 15144
rect 9263 15113 9275 15116
rect 9217 15107 9275 15113
rect 9858 15104 9864 15116
rect 9916 15104 9922 15156
rect 10042 15144 10048 15156
rect 10003 15116 10048 15144
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 11701 15147 11759 15153
rect 11701 15144 11713 15147
rect 10152 15116 11713 15144
rect 8110 15076 8116 15088
rect 6748 15048 7052 15076
rect 6748 15020 6776 15048
rect 5445 15011 5503 15017
rect 5445 15008 5457 15011
rect 4908 14980 5457 15008
rect 5445 14977 5457 14980
rect 5491 14977 5503 15011
rect 5445 14971 5503 14977
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 6730 15008 6736 15020
rect 5675 14980 6736 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 6914 14968 6920 15020
rect 6972 14968 6978 15020
rect 7024 15017 7052 15048
rect 7392 15048 8116 15076
rect 7392 15017 7420 15048
rect 8110 15036 8116 15048
rect 8168 15036 8174 15088
rect 10152 15076 10180 15116
rect 11701 15113 11713 15116
rect 11747 15113 11759 15147
rect 14458 15144 14464 15156
rect 14419 15116 14464 15144
rect 11701 15107 11759 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 15746 15144 15752 15156
rect 15707 15116 15752 15144
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 17037 15147 17095 15153
rect 17037 15144 17049 15147
rect 16040 15116 17049 15144
rect 11514 15076 11520 15088
rect 10060 15048 10180 15076
rect 11475 15048 11520 15076
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 14977 7067 15011
rect 7009 14971 7067 14977
rect 7377 15011 7435 15017
rect 7377 14977 7389 15011
rect 7423 14977 7435 15011
rect 7558 15008 7564 15020
rect 7519 14980 7564 15008
rect 7377 14971 7435 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 15008 8723 15011
rect 9214 15008 9220 15020
rect 8711 14980 9220 15008
rect 8711 14977 8723 14980
rect 8665 14971 8723 14977
rect 9214 14968 9220 14980
rect 9272 14968 9278 15020
rect 9398 14968 9404 15020
rect 9456 14968 9462 15020
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 9585 15011 9643 15017
rect 9585 14977 9597 15011
rect 9631 15008 9643 15011
rect 10060 15008 10088 15048
rect 11514 15036 11520 15048
rect 11572 15036 11578 15088
rect 11882 15036 11888 15088
rect 11940 15076 11946 15088
rect 11940 15048 13124 15076
rect 11940 15036 11946 15048
rect 9631 14980 10088 15008
rect 9631 14977 9643 14980
rect 9585 14971 9643 14977
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14940 2099 14943
rect 3142 14940 3148 14952
rect 2087 14912 3148 14940
rect 2087 14909 2099 14912
rect 2041 14903 2099 14909
rect 3142 14900 3148 14912
rect 3200 14940 3206 14952
rect 3528 14940 3556 14968
rect 3200 14912 3556 14940
rect 3200 14900 3206 14912
rect 5258 14900 5264 14952
rect 5316 14940 5322 14952
rect 5353 14943 5411 14949
rect 5353 14940 5365 14943
rect 5316 14912 5365 14940
rect 5316 14900 5322 14912
rect 5353 14909 5365 14912
rect 5399 14909 5411 14943
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 5353 14903 5411 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6932 14940 6960 14968
rect 7653 14943 7711 14949
rect 7653 14940 7665 14943
rect 6932 14912 7665 14940
rect 7653 14909 7665 14912
rect 7699 14940 7711 14943
rect 7926 14940 7932 14952
rect 7699 14912 7932 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 7926 14900 7932 14912
rect 7984 14900 7990 14952
rect 8113 14943 8171 14949
rect 8113 14940 8125 14943
rect 8036 14912 8125 14940
rect 2222 14832 2228 14884
rect 2280 14881 2286 14884
rect 2280 14875 2344 14881
rect 2280 14841 2298 14875
rect 2332 14841 2344 14875
rect 3780 14875 3838 14881
rect 3780 14872 3792 14875
rect 2280 14835 2344 14841
rect 3436 14844 3792 14872
rect 2280 14832 2286 14835
rect 3436 14813 3464 14844
rect 3780 14841 3792 14844
rect 3826 14872 3838 14875
rect 4062 14872 4068 14884
rect 3826 14844 4068 14872
rect 3826 14841 3838 14844
rect 3780 14835 3838 14841
rect 4062 14832 4068 14844
rect 4120 14832 4126 14884
rect 5994 14832 6000 14884
rect 6052 14872 6058 14884
rect 6917 14875 6975 14881
rect 6917 14872 6929 14875
rect 6052 14844 6929 14872
rect 6052 14832 6058 14844
rect 6917 14841 6929 14844
rect 6963 14841 6975 14875
rect 6917 14835 6975 14841
rect 8036 14813 8064 14912
rect 8113 14909 8125 14912
rect 8159 14909 8171 14943
rect 8113 14903 8171 14909
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14940 8907 14943
rect 9416 14940 9444 14968
rect 8895 14912 9444 14940
rect 8895 14909 8907 14912
rect 8849 14903 8907 14909
rect 8757 14875 8815 14881
rect 8757 14841 8769 14875
rect 8803 14872 8815 14875
rect 8803 14844 9352 14872
rect 8803 14841 8815 14844
rect 8757 14835 8815 14841
rect 3421 14807 3479 14813
rect 3421 14773 3433 14807
rect 3467 14773 3479 14807
rect 3421 14767 3479 14773
rect 8021 14807 8079 14813
rect 8021 14773 8033 14807
rect 8067 14773 8079 14807
rect 9324 14804 9352 14844
rect 9398 14832 9404 14884
rect 9456 14872 9462 14884
rect 9508 14872 9536 14971
rect 10134 14968 10140 15020
rect 10192 15008 10198 15020
rect 10192 14980 10237 15008
rect 10192 14968 10198 14980
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 13096 15017 13124 15048
rect 12253 15011 12311 15017
rect 12253 15008 12265 15011
rect 12032 14980 12265 15008
rect 12032 14968 12038 14980
rect 12253 14977 12265 14980
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 13081 15011 13139 15017
rect 13081 14977 13093 15011
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 15197 15011 15255 15017
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 16040 15008 16068 15116
rect 17037 15113 17049 15116
rect 17083 15113 17095 15147
rect 18138 15144 18144 15156
rect 18099 15116 18144 15144
rect 17037 15107 17095 15113
rect 18138 15104 18144 15116
rect 18196 15104 18202 15156
rect 18414 15104 18420 15156
rect 18472 15104 18478 15156
rect 19150 15104 19156 15156
rect 19208 15144 19214 15156
rect 20622 15144 20628 15156
rect 19208 15116 20628 15144
rect 19208 15104 19214 15116
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 20806 15104 20812 15156
rect 20864 15144 20870 15156
rect 21269 15147 21327 15153
rect 21269 15144 21281 15147
rect 20864 15116 21281 15144
rect 20864 15104 20870 15116
rect 21269 15113 21281 15116
rect 21315 15113 21327 15147
rect 21269 15107 21327 15113
rect 16114 15036 16120 15088
rect 16172 15076 16178 15088
rect 16172 15048 16344 15076
rect 16172 15036 16178 15048
rect 16206 15008 16212 15020
rect 15243 14980 16068 15008
rect 16167 14980 16212 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 16206 14968 16212 14980
rect 16264 14968 16270 15020
rect 16316 15017 16344 15048
rect 16390 15036 16396 15088
rect 16448 15076 16454 15088
rect 18432 15076 18460 15104
rect 22186 15076 22192 15088
rect 16448 15048 18460 15076
rect 22066 15048 22192 15076
rect 16448 15036 16454 15048
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 17770 14968 17776 15020
rect 17828 15008 17834 15020
rect 18417 15011 18475 15017
rect 18417 15008 18429 15011
rect 17828 14980 18429 15008
rect 17828 14968 17834 14980
rect 18417 14977 18429 14980
rect 18463 14977 18475 15011
rect 22066 15008 22094 15048
rect 22186 15036 22192 15048
rect 22244 15036 22250 15088
rect 22278 15008 22284 15020
rect 18417 14971 18475 14977
rect 19720 14980 20024 15008
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14940 9735 14943
rect 11330 14940 11336 14952
rect 9723 14912 11336 14940
rect 9723 14909 9735 14912
rect 9677 14903 9735 14909
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 11882 14900 11888 14952
rect 11940 14940 11946 14952
rect 12158 14940 12164 14952
rect 11940 14912 12164 14940
rect 11940 14900 11946 14912
rect 12158 14900 12164 14912
rect 12216 14900 12222 14952
rect 12526 14940 12532 14952
rect 12487 14912 12532 14940
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 13354 14949 13360 14952
rect 13348 14903 13360 14949
rect 13412 14940 13418 14952
rect 13412 14912 13448 14940
rect 13354 14900 13360 14903
rect 13412 14900 13418 14912
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 17218 14940 17224 14952
rect 15528 14912 15573 14940
rect 17179 14912 17224 14940
rect 15528 14900 15534 14912
rect 17218 14900 17224 14912
rect 17276 14900 17282 14952
rect 18046 14940 18052 14952
rect 18007 14912 18052 14940
rect 18046 14900 18052 14912
rect 18104 14940 18110 14952
rect 18325 14943 18383 14949
rect 18325 14940 18337 14943
rect 18104 14912 18337 14940
rect 18104 14900 18110 14912
rect 18325 14909 18337 14912
rect 18371 14909 18383 14943
rect 19720 14940 19748 14980
rect 19886 14940 19892 14952
rect 18325 14903 18383 14909
rect 18616 14912 19748 14940
rect 19847 14912 19892 14940
rect 10382 14875 10440 14881
rect 10382 14872 10394 14875
rect 9456 14844 10394 14872
rect 9456 14832 9462 14844
rect 10382 14841 10394 14844
rect 10428 14841 10440 14875
rect 10382 14835 10440 14841
rect 12713 14875 12771 14881
rect 12713 14841 12725 14875
rect 12759 14872 12771 14875
rect 12802 14872 12808 14884
rect 12759 14844 12808 14872
rect 12759 14841 12771 14844
rect 12713 14835 12771 14841
rect 12802 14832 12808 14844
rect 12860 14832 12866 14884
rect 13814 14832 13820 14884
rect 13872 14872 13878 14884
rect 13872 14844 14596 14872
rect 13872 14832 13878 14844
rect 10962 14804 10968 14816
rect 9324 14776 10968 14804
rect 8021 14767 8079 14773
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11054 14764 11060 14816
rect 11112 14804 11118 14816
rect 11606 14804 11612 14816
rect 11112 14776 11612 14804
rect 11112 14764 11118 14776
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 12069 14807 12127 14813
rect 12069 14804 12081 14807
rect 11848 14776 12081 14804
rect 11848 14764 11854 14776
rect 12069 14773 12081 14776
rect 12115 14773 12127 14807
rect 12069 14767 12127 14773
rect 12158 14764 12164 14816
rect 12216 14804 12222 14816
rect 12897 14807 12955 14813
rect 12216 14776 12261 14804
rect 12216 14764 12222 14776
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 13722 14804 13728 14816
rect 12943 14776 13728 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 13722 14764 13728 14776
rect 13780 14764 13786 14816
rect 14568 14813 14596 14844
rect 14642 14832 14648 14884
rect 14700 14872 14706 14884
rect 15013 14875 15071 14881
rect 15013 14872 15025 14875
rect 14700 14844 15025 14872
rect 14700 14832 14706 14844
rect 15013 14841 15025 14844
rect 15059 14841 15071 14875
rect 15013 14835 15071 14841
rect 16117 14875 16175 14881
rect 16117 14841 16129 14875
rect 16163 14872 16175 14875
rect 16577 14875 16635 14881
rect 16577 14872 16589 14875
rect 16163 14844 16589 14872
rect 16163 14841 16175 14844
rect 16117 14835 16175 14841
rect 16577 14841 16589 14844
rect 16623 14841 16635 14875
rect 16577 14835 16635 14841
rect 17037 14875 17095 14881
rect 17037 14841 17049 14875
rect 17083 14872 17095 14875
rect 17494 14872 17500 14884
rect 17083 14844 17500 14872
rect 17083 14841 17095 14844
rect 17037 14835 17095 14841
rect 17494 14832 17500 14844
rect 17552 14872 17558 14884
rect 17589 14875 17647 14881
rect 17589 14872 17601 14875
rect 17552 14844 17601 14872
rect 17552 14832 17558 14844
rect 17589 14841 17601 14844
rect 17635 14841 17647 14875
rect 17589 14835 17647 14841
rect 14553 14807 14611 14813
rect 14553 14773 14565 14807
rect 14599 14773 14611 14807
rect 14918 14804 14924 14816
rect 14879 14776 14924 14804
rect 14553 14767 14611 14773
rect 14918 14764 14924 14776
rect 14976 14764 14982 14816
rect 15562 14764 15568 14816
rect 15620 14804 15626 14816
rect 15657 14807 15715 14813
rect 15657 14804 15669 14807
rect 15620 14776 15669 14804
rect 15620 14764 15626 14776
rect 15657 14773 15669 14776
rect 15703 14804 15715 14807
rect 16298 14804 16304 14816
rect 15703 14776 16304 14804
rect 15703 14773 15715 14776
rect 15657 14767 15715 14773
rect 16298 14764 16304 14776
rect 16356 14764 16362 14816
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 18616 14804 18644 14912
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 19996 14940 20024 14980
rect 21560 14980 22094 15008
rect 22239 14980 22284 15008
rect 20714 14940 20720 14952
rect 19996 14912 20720 14940
rect 20714 14900 20720 14912
rect 20772 14900 20778 14952
rect 21560 14949 21588 14980
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 22465 15011 22523 15017
rect 22465 14977 22477 15011
rect 22511 15008 22523 15011
rect 22922 15008 22928 15020
rect 22511 14980 22928 15008
rect 22511 14977 22523 14980
rect 22465 14971 22523 14977
rect 22922 14968 22928 14980
rect 22980 14968 22986 15020
rect 21545 14943 21603 14949
rect 21545 14909 21557 14943
rect 21591 14909 21603 14943
rect 21545 14903 21603 14909
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 22557 14943 22615 14949
rect 22557 14940 22569 14943
rect 22152 14912 22569 14940
rect 22152 14900 22158 14912
rect 22557 14909 22569 14912
rect 22603 14909 22615 14943
rect 22557 14903 22615 14909
rect 18684 14875 18742 14881
rect 18684 14841 18696 14875
rect 18730 14872 18742 14875
rect 19242 14872 19248 14884
rect 18730 14844 19248 14872
rect 18730 14841 18742 14844
rect 18684 14835 18742 14841
rect 19242 14832 19248 14844
rect 19300 14832 19306 14884
rect 19978 14872 19984 14884
rect 19812 14844 19984 14872
rect 18472 14776 18644 14804
rect 18472 14764 18478 14776
rect 18874 14764 18880 14816
rect 18932 14804 18938 14816
rect 19518 14804 19524 14816
rect 18932 14776 19524 14804
rect 18932 14764 18938 14776
rect 19518 14764 19524 14776
rect 19576 14764 19582 14816
rect 19812 14813 19840 14844
rect 19978 14832 19984 14844
rect 20036 14872 20042 14884
rect 20134 14875 20192 14881
rect 20134 14872 20146 14875
rect 20036 14844 20146 14872
rect 20036 14832 20042 14844
rect 20134 14841 20146 14844
rect 20180 14841 20192 14875
rect 20134 14835 20192 14841
rect 19797 14807 19855 14813
rect 19797 14773 19809 14807
rect 19843 14773 19855 14807
rect 19797 14767 19855 14773
rect 19886 14764 19892 14816
rect 19944 14804 19950 14816
rect 20438 14804 20444 14816
rect 19944 14776 20444 14804
rect 19944 14764 19950 14776
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 21358 14804 21364 14816
rect 21319 14776 21364 14804
rect 21358 14764 21364 14776
rect 21416 14764 21422 14816
rect 22005 14807 22063 14813
rect 22005 14773 22017 14807
rect 22051 14804 22063 14807
rect 22462 14804 22468 14816
rect 22051 14776 22468 14804
rect 22051 14773 22063 14776
rect 22005 14767 22063 14773
rect 22462 14764 22468 14776
rect 22520 14764 22526 14816
rect 22925 14807 22983 14813
rect 22925 14773 22937 14807
rect 22971 14804 22983 14807
rect 23569 14807 23627 14813
rect 23569 14804 23581 14807
rect 22971 14776 23581 14804
rect 22971 14773 22983 14776
rect 22925 14767 22983 14773
rect 23569 14773 23581 14776
rect 23615 14773 23627 14807
rect 23569 14767 23627 14773
rect 1104 14714 23460 14736
rect 1104 14662 8446 14714
rect 8498 14662 8510 14714
rect 8562 14662 8574 14714
rect 8626 14662 8638 14714
rect 8690 14662 15910 14714
rect 15962 14662 15974 14714
rect 16026 14662 16038 14714
rect 16090 14662 16102 14714
rect 16154 14662 23460 14714
rect 1104 14640 23460 14662
rect 4065 14603 4123 14609
rect 4065 14569 4077 14603
rect 4111 14600 4123 14603
rect 4154 14600 4160 14612
rect 4111 14572 4160 14600
rect 4111 14569 4123 14572
rect 4065 14563 4123 14569
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 5994 14600 6000 14612
rect 5955 14572 6000 14600
rect 5994 14560 6000 14572
rect 6052 14560 6058 14612
rect 6917 14603 6975 14609
rect 6917 14569 6929 14603
rect 6963 14600 6975 14603
rect 7282 14600 7288 14612
rect 6963 14572 7288 14600
rect 6963 14569 6975 14572
rect 6917 14563 6975 14569
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 12529 14603 12587 14609
rect 9140 14572 12388 14600
rect 2866 14492 2872 14544
rect 2924 14541 2930 14544
rect 2924 14532 2936 14541
rect 4884 14535 4942 14541
rect 2924 14504 2969 14532
rect 2924 14495 2936 14504
rect 4884 14501 4896 14535
rect 4930 14532 4942 14535
rect 5258 14532 5264 14544
rect 4930 14504 5264 14532
rect 4930 14501 4942 14504
rect 4884 14495 4942 14501
rect 2924 14492 2930 14495
rect 5258 14492 5264 14504
rect 5316 14492 5322 14544
rect 7190 14492 7196 14544
rect 7248 14532 7254 14544
rect 7438 14535 7496 14541
rect 7438 14532 7450 14535
rect 7248 14504 7450 14532
rect 7248 14492 7254 14504
rect 7438 14501 7450 14504
rect 7484 14501 7496 14535
rect 7438 14495 7496 14501
rect 3142 14464 3148 14476
rect 3103 14436 3148 14464
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 3878 14464 3884 14476
rect 3839 14436 3884 14464
rect 3878 14424 3884 14436
rect 3936 14424 3942 14476
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6270 14464 6276 14476
rect 6227 14436 6276 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6270 14424 6276 14436
rect 6328 14424 6334 14476
rect 7101 14467 7159 14473
rect 7101 14433 7113 14467
rect 7147 14464 7159 14467
rect 8754 14464 8760 14476
rect 7147 14436 8616 14464
rect 8715 14436 8760 14464
rect 7147 14433 7159 14436
rect 7101 14427 7159 14433
rect 3160 14396 3188 14424
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 3160 14368 4629 14396
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 6730 14396 6736 14408
rect 6691 14368 6736 14396
rect 4617 14359 4675 14365
rect 6730 14356 6736 14368
rect 6788 14356 6794 14408
rect 7190 14396 7196 14408
rect 7151 14368 7196 14396
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 8588 14396 8616 14436
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 9140 14473 9168 14572
rect 11149 14535 11207 14541
rect 11149 14532 11161 14535
rect 9784 14504 11161 14532
rect 9125 14467 9183 14473
rect 9125 14433 9137 14467
rect 9171 14433 9183 14467
rect 9125 14427 9183 14433
rect 8846 14396 8852 14408
rect 8588 14368 8852 14396
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 9784 14396 9812 14504
rect 11149 14501 11161 14504
rect 11195 14501 11207 14535
rect 11149 14495 11207 14501
rect 11238 14492 11244 14544
rect 11296 14532 11302 14544
rect 11974 14532 11980 14544
rect 11296 14504 11341 14532
rect 11532 14504 11980 14532
rect 11296 14492 11302 14504
rect 10525 14467 10583 14473
rect 10525 14433 10537 14467
rect 10571 14464 10583 14467
rect 10571 14436 11192 14464
rect 10571 14433 10583 14436
rect 10525 14427 10583 14433
rect 10778 14396 10784 14408
rect 8956 14368 9812 14396
rect 10739 14368 10784 14396
rect 8956 14337 8984 14368
rect 10778 14356 10784 14368
rect 10836 14356 10842 14408
rect 11054 14396 11060 14408
rect 11015 14368 11060 14396
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 11164 14396 11192 14436
rect 11532 14396 11560 14504
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 12069 14535 12127 14541
rect 12069 14501 12081 14535
rect 12115 14532 12127 14535
rect 12250 14532 12256 14544
rect 12115 14504 12256 14532
rect 12115 14501 12127 14504
rect 12069 14495 12127 14501
rect 12250 14492 12256 14504
rect 12308 14492 12314 14544
rect 12360 14532 12388 14572
rect 12529 14569 12541 14603
rect 12575 14569 12587 14603
rect 13814 14600 13820 14612
rect 13775 14572 13820 14600
rect 12529 14563 12587 14569
rect 12544 14532 12572 14563
rect 13814 14560 13820 14572
rect 13872 14560 13878 14612
rect 14185 14603 14243 14609
rect 14185 14569 14197 14603
rect 14231 14569 14243 14603
rect 14185 14563 14243 14569
rect 12360 14504 12572 14532
rect 14200 14532 14228 14563
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 14369 14603 14427 14609
rect 14369 14600 14381 14603
rect 14332 14572 14381 14600
rect 14332 14560 14338 14572
rect 14369 14569 14381 14572
rect 14415 14569 14427 14603
rect 14369 14563 14427 14569
rect 15470 14560 15476 14612
rect 15528 14600 15534 14612
rect 17586 14600 17592 14612
rect 15528 14572 17592 14600
rect 15528 14560 15534 14572
rect 17586 14560 17592 14572
rect 17644 14600 17650 14612
rect 17954 14600 17960 14612
rect 17644 14572 17960 14600
rect 17644 14560 17650 14572
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 19334 14600 19340 14612
rect 18340 14572 19340 14600
rect 16574 14532 16580 14544
rect 14200 14504 14780 14532
rect 11606 14424 11612 14476
rect 11664 14464 11670 14476
rect 12897 14467 12955 14473
rect 11664 14436 11928 14464
rect 11664 14424 11670 14436
rect 11164 14368 11560 14396
rect 11698 14356 11704 14408
rect 11756 14396 11762 14408
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 11756 14368 11805 14396
rect 11756 14356 11762 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 11900 14396 11928 14436
rect 12897 14433 12909 14467
rect 12943 14433 12955 14467
rect 14550 14464 14556 14476
rect 14511 14436 14556 14464
rect 12897 14427 12955 14433
rect 11977 14399 12035 14405
rect 11977 14396 11989 14399
rect 11900 14368 11989 14396
rect 11793 14359 11851 14365
rect 11977 14365 11989 14368
rect 12023 14365 12035 14399
rect 12526 14396 12532 14408
rect 12439 14368 12532 14396
rect 11977 14359 12035 14365
rect 8941 14331 8999 14337
rect 8941 14297 8953 14331
rect 8987 14297 8999 14331
rect 9398 14328 9404 14340
rect 9359 14300 9404 14328
rect 8941 14291 8999 14297
rect 9398 14288 9404 14300
rect 9456 14288 9462 14340
rect 12158 14328 12164 14340
rect 10796 14300 12164 14328
rect 1765 14263 1823 14269
rect 1765 14229 1777 14263
rect 1811 14260 1823 14263
rect 2222 14260 2228 14272
rect 1811 14232 2228 14260
rect 1811 14229 1823 14232
rect 1765 14223 1823 14229
rect 2222 14220 2228 14232
rect 2280 14260 2286 14272
rect 3970 14260 3976 14272
rect 2280 14232 3976 14260
rect 2280 14220 2286 14232
rect 3970 14220 3976 14232
rect 4028 14220 4034 14272
rect 8478 14220 8484 14272
rect 8536 14260 8542 14272
rect 8573 14263 8631 14269
rect 8573 14260 8585 14263
rect 8536 14232 8585 14260
rect 8536 14220 8542 14232
rect 8573 14229 8585 14232
rect 8619 14229 8631 14263
rect 8573 14223 8631 14229
rect 9309 14263 9367 14269
rect 9309 14229 9321 14263
rect 9355 14260 9367 14263
rect 10796 14260 10824 14300
rect 12158 14288 12164 14300
rect 12216 14288 12222 14340
rect 12452 14337 12480 14368
rect 12526 14356 12532 14368
rect 12584 14396 12590 14408
rect 12912 14396 12940 14427
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 14752 14473 14780 14504
rect 14936 14504 16580 14532
rect 14737 14467 14795 14473
rect 14737 14433 14749 14467
rect 14783 14433 14795 14467
rect 14737 14427 14795 14433
rect 12584 14368 12940 14396
rect 12989 14399 13047 14405
rect 12584 14356 12590 14368
rect 12989 14365 13001 14399
rect 13035 14365 13047 14399
rect 12989 14359 13047 14365
rect 13173 14399 13231 14405
rect 13173 14365 13185 14399
rect 13219 14396 13231 14399
rect 13354 14396 13360 14408
rect 13219 14368 13360 14396
rect 13219 14365 13231 14368
rect 13173 14359 13231 14365
rect 12437 14331 12495 14337
rect 12437 14297 12449 14331
rect 12483 14297 12495 14331
rect 13004 14328 13032 14359
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 13633 14399 13691 14405
rect 13633 14365 13645 14399
rect 13679 14365 13691 14399
rect 13633 14359 13691 14365
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14396 13783 14399
rect 14936 14396 14964 14504
rect 16574 14492 16580 14504
rect 16632 14492 16638 14544
rect 18340 14541 18368 14572
rect 19334 14560 19340 14572
rect 19392 14560 19398 14612
rect 19978 14600 19984 14612
rect 19939 14572 19984 14600
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20254 14560 20260 14612
rect 20312 14600 20318 14612
rect 20349 14603 20407 14609
rect 20349 14600 20361 14603
rect 20312 14572 20361 14600
rect 20312 14560 20318 14572
rect 20349 14569 20361 14572
rect 20395 14569 20407 14603
rect 20349 14563 20407 14569
rect 20714 14560 20720 14612
rect 20772 14600 20778 14612
rect 20809 14603 20867 14609
rect 20809 14600 20821 14603
rect 20772 14572 20821 14600
rect 20772 14560 20778 14572
rect 20809 14569 20821 14572
rect 20855 14600 20867 14603
rect 22186 14600 22192 14612
rect 20855 14572 22192 14600
rect 20855 14569 20867 14572
rect 20809 14563 20867 14569
rect 22186 14560 22192 14572
rect 22244 14560 22250 14612
rect 22370 14560 22376 14612
rect 22428 14600 22434 14612
rect 22741 14603 22799 14609
rect 22741 14600 22753 14603
rect 22428 14572 22753 14600
rect 22428 14560 22434 14572
rect 22741 14569 22753 14572
rect 22787 14569 22799 14603
rect 22741 14563 22799 14569
rect 18325 14535 18383 14541
rect 18325 14501 18337 14535
rect 18371 14501 18383 14535
rect 18325 14495 18383 14501
rect 18509 14535 18567 14541
rect 18509 14501 18521 14535
rect 18555 14532 18567 14535
rect 22094 14532 22100 14544
rect 18555 14504 22100 14532
rect 18555 14501 18567 14504
rect 18509 14495 18567 14501
rect 22094 14492 22100 14504
rect 22152 14492 22158 14544
rect 22296 14504 22968 14532
rect 15280 14467 15338 14473
rect 15280 14433 15292 14467
rect 15326 14464 15338 14467
rect 15746 14464 15752 14476
rect 15326 14436 15752 14464
rect 15326 14433 15338 14436
rect 15280 14427 15338 14433
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 16758 14473 16764 14476
rect 16752 14427 16764 14473
rect 16816 14464 16822 14476
rect 16816 14436 16852 14464
rect 16758 14424 16764 14427
rect 16816 14424 16822 14436
rect 18046 14424 18052 14476
rect 18104 14464 18110 14476
rect 18601 14467 18659 14473
rect 18601 14464 18613 14467
rect 18104 14436 18613 14464
rect 18104 14424 18110 14436
rect 18601 14433 18613 14436
rect 18647 14433 18659 14467
rect 18601 14427 18659 14433
rect 18785 14467 18843 14473
rect 18785 14433 18797 14467
rect 18831 14433 18843 14467
rect 18785 14427 18843 14433
rect 19153 14467 19211 14473
rect 19153 14433 19165 14467
rect 19199 14464 19211 14467
rect 19245 14467 19303 14473
rect 19245 14464 19257 14467
rect 19199 14436 19257 14464
rect 19199 14433 19211 14436
rect 19153 14427 19211 14433
rect 19245 14433 19257 14436
rect 19291 14464 19303 14467
rect 19426 14464 19432 14476
rect 19291 14436 19432 14464
rect 19291 14433 19303 14436
rect 19245 14427 19303 14433
rect 13771 14368 14964 14396
rect 13771 14365 13783 14368
rect 13725 14359 13783 14365
rect 12437 14291 12495 14297
rect 12932 14300 13032 14328
rect 13648 14328 13676 14359
rect 15010 14356 15016 14408
rect 15068 14396 15074 14408
rect 15068 14368 15113 14396
rect 15068 14356 15074 14368
rect 16206 14356 16212 14408
rect 16264 14396 16270 14408
rect 16485 14399 16543 14405
rect 16485 14396 16497 14399
rect 16264 14368 16497 14396
rect 16264 14356 16270 14368
rect 16485 14365 16497 14368
rect 16531 14365 16543 14399
rect 16485 14359 16543 14365
rect 17862 14356 17868 14408
rect 17920 14356 17926 14408
rect 13814 14328 13820 14340
rect 13648 14300 13820 14328
rect 11606 14260 11612 14272
rect 9355 14232 10824 14260
rect 11567 14232 11612 14260
rect 9355 14229 9367 14232
rect 9309 14223 9367 14229
rect 11606 14220 11612 14232
rect 11664 14260 11670 14272
rect 12932 14260 12960 14300
rect 13814 14288 13820 14300
rect 13872 14288 13878 14340
rect 17880 14328 17908 14356
rect 18800 14328 18828 14427
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 19978 14464 19984 14476
rect 19628 14436 19984 14464
rect 19628 14396 19656 14436
rect 19978 14424 19984 14436
rect 20036 14424 20042 14476
rect 21174 14464 21180 14476
rect 20548 14436 21180 14464
rect 19794 14396 19800 14408
rect 18984 14368 19656 14396
rect 19755 14368 19800 14396
rect 18984 14337 19012 14368
rect 19794 14356 19800 14368
rect 19852 14356 19858 14408
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14365 19947 14399
rect 19889 14359 19947 14365
rect 17880 14300 18828 14328
rect 18969 14331 19027 14337
rect 18969 14297 18981 14331
rect 19015 14297 19027 14331
rect 18969 14291 19027 14297
rect 19242 14288 19248 14340
rect 19300 14328 19306 14340
rect 19904 14328 19932 14359
rect 19300 14300 19932 14328
rect 19300 14288 19306 14300
rect 11664 14232 12960 14260
rect 11664 14220 11670 14232
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 14921 14263 14979 14269
rect 14921 14260 14933 14263
rect 14884 14232 14933 14260
rect 14884 14220 14890 14232
rect 14921 14229 14933 14232
rect 14967 14229 14979 14263
rect 14921 14223 14979 14229
rect 16393 14263 16451 14269
rect 16393 14229 16405 14263
rect 16439 14260 16451 14263
rect 16758 14260 16764 14272
rect 16439 14232 16764 14260
rect 16439 14229 16451 14232
rect 16393 14223 16451 14229
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 17865 14263 17923 14269
rect 17865 14260 17877 14263
rect 17460 14232 17877 14260
rect 17460 14220 17466 14232
rect 17865 14229 17877 14232
rect 17911 14229 17923 14263
rect 17865 14223 17923 14229
rect 18049 14263 18107 14269
rect 18049 14229 18061 14263
rect 18095 14260 18107 14263
rect 19150 14260 19156 14272
rect 18095 14232 19156 14260
rect 18095 14229 18107 14232
rect 18049 14223 18107 14229
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 19429 14263 19487 14269
rect 19429 14229 19441 14263
rect 19475 14260 19487 14263
rect 20548 14260 20576 14436
rect 21174 14424 21180 14436
rect 21232 14424 21238 14476
rect 21634 14424 21640 14476
rect 21692 14464 21698 14476
rect 22296 14464 22324 14504
rect 21692 14436 22324 14464
rect 22393 14467 22451 14473
rect 21692 14424 21698 14436
rect 22393 14433 22405 14467
rect 22439 14464 22451 14467
rect 22554 14464 22560 14476
rect 22439 14436 22560 14464
rect 22439 14433 22451 14436
rect 22393 14427 22451 14433
rect 22554 14424 22560 14436
rect 22612 14424 22618 14476
rect 22646 14424 22652 14476
rect 22704 14464 22710 14476
rect 22940 14473 22968 14504
rect 22925 14467 22983 14473
rect 22704 14436 22749 14464
rect 22704 14424 22710 14436
rect 22925 14433 22937 14467
rect 22971 14433 22983 14467
rect 22925 14427 22983 14433
rect 20625 14399 20683 14405
rect 20625 14365 20637 14399
rect 20671 14365 20683 14399
rect 20625 14359 20683 14365
rect 20717 14399 20775 14405
rect 20717 14365 20729 14399
rect 20763 14396 20775 14399
rect 21082 14396 21088 14408
rect 20763 14368 21088 14396
rect 20763 14365 20775 14368
rect 20717 14359 20775 14365
rect 20640 14328 20668 14359
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 21177 14331 21235 14337
rect 20640 14300 20760 14328
rect 19475 14232 20576 14260
rect 20732 14260 20760 14300
rect 21177 14297 21189 14331
rect 21223 14328 21235 14331
rect 21223 14300 21680 14328
rect 21223 14297 21235 14300
rect 21177 14291 21235 14297
rect 20898 14260 20904 14272
rect 20732 14232 20904 14260
rect 19475 14229 19487 14232
rect 19429 14223 19487 14229
rect 20898 14220 20904 14232
rect 20956 14260 20962 14272
rect 21269 14263 21327 14269
rect 21269 14260 21281 14263
rect 20956 14232 21281 14260
rect 20956 14220 20962 14232
rect 21269 14229 21281 14232
rect 21315 14229 21327 14263
rect 21652 14260 21680 14300
rect 22738 14260 22744 14272
rect 21652 14232 22744 14260
rect 21269 14223 21327 14229
rect 22738 14220 22744 14232
rect 22796 14220 22802 14272
rect 1104 14170 23460 14192
rect 1104 14118 4714 14170
rect 4766 14118 4778 14170
rect 4830 14118 4842 14170
rect 4894 14118 4906 14170
rect 4958 14118 12178 14170
rect 12230 14118 12242 14170
rect 12294 14118 12306 14170
rect 12358 14118 12370 14170
rect 12422 14118 19642 14170
rect 19694 14118 19706 14170
rect 19758 14118 19770 14170
rect 19822 14118 19834 14170
rect 19886 14118 23460 14170
rect 1104 14096 23460 14118
rect 1397 14059 1455 14065
rect 1397 14025 1409 14059
rect 1443 14056 1455 14059
rect 1762 14056 1768 14068
rect 1443 14028 1768 14056
rect 1443 14025 1455 14028
rect 1397 14019 1455 14025
rect 1762 14016 1768 14028
rect 1820 14056 1826 14068
rect 1820 14028 3188 14056
rect 1820 14016 1826 14028
rect 2792 13960 3096 13988
rect 2792 13920 2820 13960
rect 2700 13892 2820 13920
rect 2521 13855 2579 13861
rect 2521 13821 2533 13855
rect 2567 13852 2579 13855
rect 2700 13852 2728 13892
rect 2866 13880 2872 13932
rect 2924 13920 2930 13932
rect 2961 13923 3019 13929
rect 2961 13920 2973 13923
rect 2924 13892 2973 13920
rect 2924 13880 2930 13892
rect 2961 13889 2973 13892
rect 3007 13889 3019 13923
rect 2961 13883 3019 13889
rect 2567 13824 2728 13852
rect 2567 13821 2579 13824
rect 2521 13815 2579 13821
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 3068 13852 3096 13960
rect 3160 13929 3188 14028
rect 3234 14016 3240 14068
rect 3292 14056 3298 14068
rect 3605 14059 3663 14065
rect 3605 14056 3617 14059
rect 3292 14028 3617 14056
rect 3292 14016 3298 14028
rect 3605 14025 3617 14028
rect 3651 14025 3663 14059
rect 3605 14019 3663 14025
rect 3694 14016 3700 14068
rect 3752 14056 3758 14068
rect 4709 14059 4767 14065
rect 3752 14028 3797 14056
rect 3752 14016 3758 14028
rect 4709 14025 4721 14059
rect 4755 14056 4767 14059
rect 5810 14056 5816 14068
rect 4755 14028 5816 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 5902 14016 5908 14068
rect 5960 14056 5966 14068
rect 5997 14059 6055 14065
rect 5997 14056 6009 14059
rect 5960 14028 6009 14056
rect 5960 14016 5966 14028
rect 5997 14025 6009 14028
rect 6043 14025 6055 14059
rect 5997 14019 6055 14025
rect 8754 14016 8760 14068
rect 8812 14056 8818 14068
rect 9677 14059 9735 14065
rect 9677 14056 9689 14059
rect 8812 14028 9689 14056
rect 8812 14016 8818 14028
rect 9677 14025 9689 14028
rect 9723 14025 9735 14059
rect 9677 14019 9735 14025
rect 10962 14016 10968 14068
rect 11020 14056 11026 14068
rect 11514 14056 11520 14068
rect 11020 14028 11520 14056
rect 11020 14016 11026 14028
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 11701 14059 11759 14065
rect 11701 14025 11713 14059
rect 11747 14056 11759 14059
rect 11974 14056 11980 14068
rect 11747 14028 11980 14056
rect 11747 14025 11759 14028
rect 11701 14019 11759 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 13265 14059 13323 14065
rect 13265 14056 13277 14059
rect 12084 14028 13277 14056
rect 5721 13991 5779 13997
rect 5721 13957 5733 13991
rect 5767 13957 5779 13991
rect 5721 13951 5779 13957
rect 9585 13991 9643 13997
rect 9585 13957 9597 13991
rect 9631 13988 9643 13991
rect 9631 13960 10180 13988
rect 9631 13957 9643 13960
rect 9585 13951 9643 13957
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13889 3203 13923
rect 3145 13883 3203 13889
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 4157 13923 4215 13929
rect 4157 13920 4169 13923
rect 4028 13892 4169 13920
rect 4028 13880 4034 13892
rect 4157 13889 4169 13892
rect 4203 13889 4215 13923
rect 4157 13883 4215 13889
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4430 13920 4436 13932
rect 4387 13892 4436 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4430 13880 4436 13892
rect 4488 13880 4494 13932
rect 5166 13920 5172 13932
rect 5079 13892 5172 13920
rect 5166 13880 5172 13892
rect 5224 13920 5230 13932
rect 5442 13920 5448 13932
rect 5224 13892 5448 13920
rect 5224 13880 5230 13892
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 4062 13852 4068 13864
rect 2832 13824 2877 13852
rect 3068 13824 3924 13852
rect 4023 13824 4068 13852
rect 2832 13812 2838 13824
rect 2958 13744 2964 13796
rect 3016 13784 3022 13796
rect 3237 13787 3295 13793
rect 3237 13784 3249 13787
rect 3016 13756 3249 13784
rect 3016 13744 3022 13756
rect 3237 13753 3249 13756
rect 3283 13753 3295 13787
rect 3896 13784 3924 13824
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4522 13852 4528 13864
rect 4483 13824 4528 13852
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 5261 13855 5319 13861
rect 5261 13821 5273 13855
rect 5307 13852 5319 13855
rect 5534 13852 5540 13864
rect 5307 13824 5540 13852
rect 5307 13821 5319 13824
rect 5261 13815 5319 13821
rect 5534 13812 5540 13824
rect 5592 13812 5598 13864
rect 5736 13852 5764 13951
rect 9033 13923 9091 13929
rect 8680 13892 8984 13920
rect 5813 13855 5871 13861
rect 5813 13852 5825 13855
rect 5736 13824 5825 13852
rect 5813 13821 5825 13824
rect 5859 13821 5871 13855
rect 5813 13815 5871 13821
rect 8478 13812 8484 13864
rect 8536 13861 8542 13864
rect 8536 13852 8548 13861
rect 8680 13852 8708 13892
rect 8536 13824 8708 13852
rect 8536 13815 8548 13824
rect 8536 13812 8542 13815
rect 8754 13812 8760 13864
rect 8812 13852 8818 13864
rect 8956 13852 8984 13892
rect 9033 13889 9045 13923
rect 9079 13920 9091 13923
rect 9306 13920 9312 13932
rect 9079 13892 9312 13920
rect 9079 13889 9091 13892
rect 9033 13883 9091 13889
rect 9306 13880 9312 13892
rect 9364 13880 9370 13932
rect 10152 13929 10180 13960
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13920 10379 13923
rect 10870 13920 10876 13932
rect 10367 13892 10876 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 10870 13880 10876 13892
rect 10928 13920 10934 13932
rect 11149 13923 11207 13929
rect 11149 13920 11161 13923
rect 10928 13892 11161 13920
rect 10928 13880 10934 13892
rect 11149 13889 11161 13892
rect 11195 13920 11207 13923
rect 12084 13920 12112 14028
rect 13265 14025 13277 14028
rect 13311 14025 13323 14059
rect 13265 14019 13323 14025
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 13541 14059 13599 14065
rect 13541 14056 13553 14059
rect 13412 14028 13553 14056
rect 13412 14016 13418 14028
rect 13541 14025 13553 14028
rect 13587 14025 13599 14059
rect 13541 14019 13599 14025
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 15749 14059 15807 14065
rect 15749 14056 15761 14059
rect 13872 14028 15761 14056
rect 13872 14016 13878 14028
rect 15749 14025 15761 14028
rect 15795 14025 15807 14059
rect 18598 14056 18604 14068
rect 15749 14019 15807 14025
rect 15856 14028 18604 14056
rect 14277 13991 14335 13997
rect 14277 13957 14289 13991
rect 14323 13988 14335 13991
rect 14550 13988 14556 14000
rect 14323 13960 14556 13988
rect 14323 13957 14335 13960
rect 14277 13951 14335 13957
rect 14550 13948 14556 13960
rect 14608 13988 14614 14000
rect 15470 13988 15476 14000
rect 14608 13960 15476 13988
rect 14608 13948 14614 13960
rect 15470 13948 15476 13960
rect 15528 13948 15534 14000
rect 13078 13920 13084 13932
rect 11195 13892 12112 13920
rect 13039 13892 13084 13920
rect 11195 13889 11207 13892
rect 11149 13883 11207 13889
rect 13078 13880 13084 13892
rect 13136 13920 13142 13932
rect 13354 13920 13360 13932
rect 13136 13892 13360 13920
rect 13136 13880 13142 13892
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 15856 13920 15884 14028
rect 18598 14016 18604 14028
rect 18656 14016 18662 14068
rect 19242 14056 19248 14068
rect 19203 14028 19248 14056
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 19705 14059 19763 14065
rect 19705 14025 19717 14059
rect 19751 14056 19763 14059
rect 22186 14056 22192 14068
rect 19751 14028 22094 14056
rect 22147 14028 22192 14056
rect 19751 14025 19763 14028
rect 19705 14019 19763 14025
rect 16117 13991 16175 13997
rect 16117 13957 16129 13991
rect 16163 13988 16175 13991
rect 16390 13988 16396 14000
rect 16163 13960 16396 13988
rect 16163 13957 16175 13960
rect 16117 13951 16175 13957
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 16592 13960 17908 13988
rect 16592 13929 16620 13960
rect 15580 13892 15884 13920
rect 16577 13923 16635 13929
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 8812 13824 8857 13852
rect 8956 13824 9137 13852
rect 8812 13812 8818 13824
rect 9125 13821 9137 13824
rect 9171 13821 9183 13855
rect 9125 13815 9183 13821
rect 10965 13855 11023 13861
rect 10965 13821 10977 13855
rect 11011 13852 11023 13855
rect 11698 13852 11704 13864
rect 11011 13824 11704 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 12802 13812 12808 13864
rect 12860 13861 12866 13864
rect 12860 13852 12872 13861
rect 12860 13824 12905 13852
rect 12860 13815 12872 13824
rect 12860 13812 12866 13815
rect 12986 13812 12992 13864
rect 13044 13852 13050 13864
rect 13722 13852 13728 13864
rect 13044 13824 13400 13852
rect 13683 13824 13728 13852
rect 13044 13812 13050 13824
rect 6546 13784 6552 13796
rect 3896 13756 6552 13784
rect 3237 13747 3295 13753
rect 6546 13744 6552 13756
rect 6604 13744 6610 13796
rect 9217 13787 9275 13793
rect 9217 13784 9229 13787
rect 8588 13756 9229 13784
rect 5353 13719 5411 13725
rect 5353 13685 5365 13719
rect 5399 13716 5411 13719
rect 6178 13716 6184 13728
rect 5399 13688 6184 13716
rect 5399 13685 5411 13688
rect 5353 13679 5411 13685
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 7377 13719 7435 13725
rect 7377 13685 7389 13719
rect 7423 13716 7435 13719
rect 7650 13716 7656 13728
rect 7423 13688 7656 13716
rect 7423 13685 7435 13688
rect 7377 13679 7435 13685
rect 7650 13676 7656 13688
rect 7708 13716 7714 13728
rect 8588 13716 8616 13756
rect 9217 13753 9229 13756
rect 9263 13753 9275 13787
rect 11330 13784 11336 13796
rect 11291 13756 11336 13784
rect 9217 13747 9275 13753
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 13372 13793 13400 13824
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 15580 13861 15608 13892
rect 16577 13889 16589 13923
rect 16623 13889 16635 13923
rect 16577 13883 16635 13889
rect 16666 13880 16672 13932
rect 16724 13920 16730 13932
rect 17402 13920 17408 13932
rect 16724 13892 16769 13920
rect 17363 13892 17408 13920
rect 16724 13880 16730 13892
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 17494 13880 17500 13932
rect 17552 13920 17558 13932
rect 17880 13920 17908 13960
rect 19426 13948 19432 14000
rect 19484 13988 19490 14000
rect 20254 13988 20260 14000
rect 19484 13960 20260 13988
rect 19484 13948 19490 13960
rect 20254 13948 20260 13960
rect 20312 13948 20318 14000
rect 22066 13988 22094 14028
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 22278 13988 22284 14000
rect 22066 13960 22284 13988
rect 22278 13948 22284 13960
rect 22336 13948 22342 14000
rect 17552 13892 17597 13920
rect 17880 13892 18000 13920
rect 17552 13880 17558 13892
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 15841 13855 15899 13861
rect 15841 13821 15853 13855
rect 15887 13852 15899 13855
rect 16482 13852 16488 13864
rect 15887 13824 16488 13852
rect 15887 13821 15899 13824
rect 15841 13815 15899 13821
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 17126 13812 17132 13864
rect 17184 13852 17190 13864
rect 17512 13852 17540 13880
rect 17770 13852 17776 13864
rect 17184 13824 17540 13852
rect 17683 13824 17776 13852
rect 17184 13812 17190 13824
rect 17770 13812 17776 13824
rect 17828 13852 17834 13864
rect 17865 13855 17923 13861
rect 17865 13852 17877 13855
rect 17828 13824 17877 13852
rect 17828 13812 17834 13824
rect 17865 13821 17877 13824
rect 17911 13821 17923 13855
rect 17972 13852 18000 13892
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 20070 13920 20076 13932
rect 19208 13892 20076 13920
rect 19208 13880 19214 13892
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 20441 13923 20499 13929
rect 20441 13889 20453 13923
rect 20487 13920 20499 13923
rect 20487 13892 20760 13920
rect 20487 13889 20499 13892
rect 20441 13883 20499 13889
rect 20732 13864 20760 13892
rect 22554 13880 22560 13932
rect 22612 13920 22618 13932
rect 22741 13923 22799 13929
rect 22741 13920 22753 13923
rect 22612 13892 22753 13920
rect 22612 13880 22618 13892
rect 22741 13889 22753 13892
rect 22787 13889 22799 13923
rect 22741 13883 22799 13889
rect 19242 13852 19248 13864
rect 17972 13824 19248 13852
rect 17865 13815 17923 13821
rect 19242 13812 19248 13824
rect 19300 13812 19306 13864
rect 19429 13855 19487 13861
rect 19429 13821 19441 13855
rect 19475 13852 19487 13855
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19475 13824 19533 13852
rect 19475 13821 19487 13824
rect 19429 13815 19487 13821
rect 19521 13821 19533 13824
rect 19567 13852 19579 13855
rect 20346 13852 20352 13864
rect 19567 13824 20352 13852
rect 19567 13821 19579 13824
rect 19521 13815 19579 13821
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 20625 13855 20683 13861
rect 20625 13821 20637 13855
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 13357 13787 13415 13793
rect 13357 13753 13369 13787
rect 13403 13753 13415 13787
rect 13357 13747 13415 13753
rect 16577 13787 16635 13793
rect 16577 13753 16589 13787
rect 16623 13784 16635 13787
rect 18132 13787 18190 13793
rect 16623 13756 18092 13784
rect 16623 13753 16635 13756
rect 16577 13747 16635 13753
rect 7708 13688 8616 13716
rect 7708 13676 7714 13688
rect 9858 13676 9864 13728
rect 9916 13716 9922 13728
rect 10045 13719 10103 13725
rect 10045 13716 10057 13719
rect 9916 13688 10057 13716
rect 9916 13676 9922 13688
rect 10045 13685 10057 13688
rect 10091 13685 10103 13719
rect 10502 13716 10508 13728
rect 10463 13688 10508 13716
rect 10045 13679 10103 13685
rect 10502 13676 10508 13688
rect 10560 13676 10566 13728
rect 10778 13676 10784 13728
rect 10836 13716 10842 13728
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 10836 13688 10885 13716
rect 10836 13676 10842 13688
rect 10873 13685 10885 13688
rect 10919 13685 10931 13719
rect 16942 13716 16948 13728
rect 16903 13688 16948 13716
rect 10873 13679 10931 13685
rect 16942 13676 16948 13688
rect 17000 13676 17006 13728
rect 17310 13716 17316 13728
rect 17271 13688 17316 13716
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 17494 13676 17500 13728
rect 17552 13716 17558 13728
rect 17773 13719 17831 13725
rect 17773 13716 17785 13719
rect 17552 13688 17785 13716
rect 17552 13676 17558 13688
rect 17773 13685 17785 13688
rect 17819 13685 17831 13719
rect 18064 13716 18092 13756
rect 18132 13753 18144 13787
rect 18178 13784 18190 13787
rect 18322 13784 18328 13796
rect 18178 13756 18328 13784
rect 18178 13753 18190 13756
rect 18132 13747 18190 13753
rect 18322 13744 18328 13756
rect 18380 13744 18386 13796
rect 20162 13784 20168 13796
rect 20123 13756 20168 13784
rect 20162 13744 20168 13756
rect 20220 13744 20226 13796
rect 20257 13787 20315 13793
rect 20257 13753 20269 13787
rect 20303 13784 20315 13787
rect 20438 13784 20444 13796
rect 20303 13756 20444 13784
rect 20303 13753 20315 13756
rect 20257 13747 20315 13753
rect 20438 13744 20444 13756
rect 20496 13744 20502 13796
rect 20640 13784 20668 13815
rect 20714 13812 20720 13864
rect 20772 13812 20778 13864
rect 20898 13861 20904 13864
rect 20892 13852 20904 13861
rect 20859 13824 20904 13852
rect 20892 13815 20904 13824
rect 20898 13812 20904 13815
rect 20956 13812 20962 13864
rect 22649 13855 22707 13861
rect 22649 13821 22661 13855
rect 22695 13852 22707 13855
rect 23569 13855 23627 13861
rect 23569 13852 23581 13855
rect 22695 13824 23581 13852
rect 22695 13821 22707 13824
rect 22649 13815 22707 13821
rect 23569 13821 23581 13824
rect 23615 13821 23627 13855
rect 23569 13815 23627 13821
rect 21450 13784 21456 13796
rect 20640 13756 21456 13784
rect 21450 13744 21456 13756
rect 21508 13744 21514 13796
rect 21818 13784 21824 13796
rect 21560 13756 21824 13784
rect 19797 13719 19855 13725
rect 19797 13716 19809 13719
rect 18064 13688 19809 13716
rect 17773 13679 17831 13685
rect 19797 13685 19809 13688
rect 19843 13685 19855 13719
rect 20456 13716 20484 13744
rect 21560 13716 21588 13756
rect 21818 13744 21824 13756
rect 21876 13784 21882 13796
rect 21876 13756 22140 13784
rect 21876 13744 21882 13756
rect 20456 13688 21588 13716
rect 19797 13679 19855 13685
rect 21634 13676 21640 13728
rect 21692 13716 21698 13728
rect 22005 13719 22063 13725
rect 22005 13716 22017 13719
rect 21692 13688 22017 13716
rect 21692 13676 21698 13688
rect 22005 13685 22017 13688
rect 22051 13685 22063 13719
rect 22112 13716 22140 13756
rect 22462 13744 22468 13796
rect 22520 13784 22526 13796
rect 22557 13787 22615 13793
rect 22557 13784 22569 13787
rect 22520 13756 22569 13784
rect 22520 13744 22526 13756
rect 22557 13753 22569 13756
rect 22603 13753 22615 13787
rect 22557 13747 22615 13753
rect 23017 13719 23075 13725
rect 23017 13716 23029 13719
rect 22112 13688 23029 13716
rect 22005 13679 22063 13685
rect 23017 13685 23029 13688
rect 23063 13685 23075 13719
rect 23017 13679 23075 13685
rect 1104 13626 23460 13648
rect 1104 13574 8446 13626
rect 8498 13574 8510 13626
rect 8562 13574 8574 13626
rect 8626 13574 8638 13626
rect 8690 13574 15910 13626
rect 15962 13574 15974 13626
rect 16026 13574 16038 13626
rect 16090 13574 16102 13626
rect 16154 13574 23460 13626
rect 1104 13552 23460 13574
rect 3329 13515 3387 13521
rect 3329 13481 3341 13515
rect 3375 13512 3387 13515
rect 3881 13515 3939 13521
rect 3881 13512 3893 13515
rect 3375 13484 3893 13512
rect 3375 13481 3387 13484
rect 3329 13475 3387 13481
rect 3881 13481 3893 13484
rect 3927 13481 3939 13515
rect 6178 13512 6184 13524
rect 6139 13484 6184 13512
rect 3881 13475 3939 13481
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 6546 13512 6552 13524
rect 6507 13484 6552 13512
rect 6546 13472 6552 13484
rect 6604 13472 6610 13524
rect 7926 13472 7932 13524
rect 7984 13512 7990 13524
rect 8757 13515 8815 13521
rect 7984 13484 8432 13512
rect 7984 13472 7990 13484
rect 5166 13444 5172 13456
rect 3252 13416 5172 13444
rect 3252 13376 3280 13416
rect 5166 13404 5172 13416
rect 5224 13404 5230 13456
rect 7650 13453 7656 13456
rect 7644 13444 7656 13453
rect 7611 13416 7656 13444
rect 7644 13407 7656 13416
rect 7650 13404 7656 13407
rect 7708 13404 7714 13456
rect 8294 13404 8300 13456
rect 8352 13404 8358 13456
rect 8404 13444 8432 13484
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9030 13512 9036 13524
rect 8803 13484 9036 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 9030 13472 9036 13484
rect 9088 13512 9094 13524
rect 9401 13515 9459 13521
rect 9401 13512 9413 13515
rect 9088 13484 9413 13512
rect 9088 13472 9094 13484
rect 9401 13481 9413 13484
rect 9447 13481 9459 13515
rect 9858 13512 9864 13524
rect 9819 13484 9864 13512
rect 9401 13475 9459 13481
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 11790 13512 11796 13524
rect 10183 13484 11796 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 11790 13472 11796 13484
rect 11848 13472 11854 13524
rect 12437 13515 12495 13521
rect 12437 13481 12449 13515
rect 12483 13512 12495 13515
rect 12802 13512 12808 13524
rect 12483 13484 12808 13512
rect 12483 13481 12495 13484
rect 12437 13475 12495 13481
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 15102 13512 15108 13524
rect 13955 13484 15108 13512
rect 9493 13447 9551 13453
rect 9493 13444 9505 13447
rect 8404 13416 9505 13444
rect 9493 13413 9505 13416
rect 9539 13413 9551 13447
rect 11606 13444 11612 13456
rect 9493 13407 9551 13413
rect 9968 13416 11612 13444
rect 4246 13376 4252 13388
rect 3068 13348 3280 13376
rect 4207 13348 4252 13376
rect 3068 13317 3096 13348
rect 4246 13336 4252 13348
rect 4304 13336 4310 13388
rect 4976 13379 5034 13385
rect 4976 13345 4988 13379
rect 5022 13376 5034 13379
rect 5442 13376 5448 13388
rect 5022 13348 5448 13376
rect 5022 13345 5034 13348
rect 4976 13339 5034 13345
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 7193 13379 7251 13385
rect 7193 13345 7205 13379
rect 7239 13376 7251 13379
rect 8312 13376 8340 13404
rect 9968 13385 9996 13416
rect 11606 13404 11612 13416
rect 11664 13404 11670 13456
rect 13955 13453 13983 13484
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17405 13515 17463 13521
rect 17405 13512 17417 13515
rect 17368 13484 17417 13512
rect 17368 13472 17374 13484
rect 17405 13481 17417 13484
rect 17451 13481 17463 13515
rect 17405 13475 17463 13481
rect 13940 13447 13998 13453
rect 13940 13413 13952 13447
rect 13986 13413 13998 13447
rect 13940 13407 13998 13413
rect 14636 13447 14694 13453
rect 14636 13413 14648 13447
rect 14682 13444 14694 13447
rect 14918 13444 14924 13456
rect 14682 13416 14924 13444
rect 14682 13413 14694 13416
rect 14636 13407 14694 13413
rect 14918 13404 14924 13416
rect 14976 13404 14982 13456
rect 17420 13444 17448 13475
rect 18322 13472 18328 13524
rect 18380 13512 18386 13524
rect 18598 13512 18604 13524
rect 18380 13484 18604 13512
rect 18380 13472 18386 13484
rect 18598 13472 18604 13484
rect 18656 13512 18662 13524
rect 18656 13484 22600 13512
rect 18656 13472 18662 13484
rect 17742 13447 17800 13453
rect 17742 13444 17754 13447
rect 17420 13416 17754 13444
rect 17742 13413 17754 13416
rect 17788 13413 17800 13447
rect 17742 13407 17800 13413
rect 18690 13404 18696 13456
rect 18748 13444 18754 13456
rect 18969 13447 19027 13453
rect 18969 13444 18981 13447
rect 18748 13416 18981 13444
rect 18748 13404 18754 13416
rect 18969 13413 18981 13416
rect 19015 13413 19027 13447
rect 18969 13407 19027 13413
rect 19076 13416 20024 13444
rect 7239 13348 8340 13376
rect 9953 13379 10011 13385
rect 7239 13345 7251 13348
rect 7193 13339 7251 13345
rect 9953 13345 9965 13379
rect 9999 13345 10011 13379
rect 10594 13376 10600 13388
rect 10555 13348 10600 13376
rect 9953 13339 10011 13345
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 11146 13336 11152 13388
rect 11204 13376 11210 13388
rect 11313 13379 11371 13385
rect 11313 13376 11325 13379
rect 11204 13348 11325 13376
rect 11204 13336 11210 13348
rect 11313 13345 11325 13348
rect 11359 13345 11371 13379
rect 12526 13376 12532 13388
rect 12487 13348 12532 13376
rect 11313 13339 11371 13345
rect 12526 13336 12532 13348
rect 12584 13336 12590 13388
rect 13446 13336 13452 13388
rect 13504 13376 13510 13388
rect 14185 13379 14243 13385
rect 14185 13376 14197 13379
rect 13504 13348 14197 13376
rect 13504 13336 13510 13348
rect 14185 13345 14197 13348
rect 14231 13376 14243 13379
rect 14369 13379 14427 13385
rect 14369 13376 14381 13379
rect 14231 13348 14381 13376
rect 14231 13345 14243 13348
rect 14185 13339 14243 13345
rect 14369 13345 14381 13348
rect 14415 13376 14427 13379
rect 15010 13376 15016 13388
rect 14415 13348 15016 13376
rect 14415 13345 14427 13348
rect 14369 13339 14427 13345
rect 15010 13336 15016 13348
rect 15068 13376 15074 13388
rect 16022 13376 16028 13388
rect 15068 13348 16028 13376
rect 15068 13336 15074 13348
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16292 13379 16350 13385
rect 16292 13345 16304 13379
rect 16338 13376 16350 13379
rect 17402 13376 17408 13388
rect 16338 13348 17408 13376
rect 16338 13345 16350 13348
rect 16292 13339 16350 13345
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 18322 13336 18328 13388
rect 18380 13376 18386 13388
rect 19076 13376 19104 13416
rect 19996 13385 20024 13416
rect 18380 13348 19104 13376
rect 19153 13379 19211 13385
rect 18380 13336 18386 13348
rect 18708 13320 18736 13348
rect 19153 13345 19165 13379
rect 19199 13345 19211 13379
rect 19153 13339 19211 13345
rect 19337 13379 19395 13385
rect 19337 13345 19349 13379
rect 19383 13376 19395 13379
rect 19797 13379 19855 13385
rect 19797 13376 19809 13379
rect 19383 13348 19809 13376
rect 19383 13345 19395 13348
rect 19337 13339 19395 13345
rect 19797 13345 19809 13348
rect 19843 13345 19855 13379
rect 19797 13339 19855 13345
rect 19981 13379 20039 13385
rect 19981 13345 19993 13379
rect 20027 13345 20039 13379
rect 20806 13376 20812 13388
rect 19981 13339 20039 13345
rect 20502 13348 20812 13376
rect 3053 13311 3111 13317
rect 3053 13277 3065 13311
rect 3099 13277 3111 13311
rect 3234 13308 3240 13320
rect 3195 13280 3240 13308
rect 3053 13271 3111 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 4338 13308 4344 13320
rect 4299 13280 4344 13308
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 4430 13268 4436 13320
rect 4488 13308 4494 13320
rect 4488 13280 4533 13308
rect 4488 13268 4494 13280
rect 4614 13268 4620 13320
rect 4672 13308 4678 13320
rect 4709 13311 4767 13317
rect 4709 13308 4721 13311
rect 4672 13280 4721 13308
rect 4672 13268 4678 13280
rect 4709 13277 4721 13280
rect 4755 13277 4767 13311
rect 6638 13308 6644 13320
rect 6599 13280 6644 13308
rect 4709 13271 4767 13277
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 6788 13280 6833 13308
rect 6788 13268 6794 13280
rect 7282 13268 7288 13320
rect 7340 13308 7346 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7340 13280 7389 13308
rect 7340 13268 7346 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 9306 13308 9312 13320
rect 9267 13280 9312 13308
rect 7377 13271 7435 13277
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 10686 13308 10692 13320
rect 10647 13280 10692 13308
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 10870 13308 10876 13320
rect 10831 13280 10876 13308
rect 10870 13268 10876 13280
rect 10928 13268 10934 13320
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13277 11115 13311
rect 17494 13308 17500 13320
rect 17455 13280 17500 13308
rect 11057 13271 11115 13277
rect 3697 13243 3755 13249
rect 3697 13209 3709 13243
rect 3743 13240 3755 13243
rect 4522 13240 4528 13252
rect 3743 13212 4528 13240
rect 3743 13209 3755 13212
rect 3697 13203 3755 13209
rect 4522 13200 4528 13212
rect 4580 13200 4586 13252
rect 10410 13200 10416 13252
rect 10468 13240 10474 13252
rect 11072 13240 11100 13271
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 18690 13268 18696 13320
rect 18748 13268 18754 13320
rect 19168 13308 19196 13339
rect 20502 13317 20530 13348
rect 20806 13336 20812 13348
rect 20864 13336 20870 13388
rect 22002 13336 22008 13388
rect 22060 13336 22066 13388
rect 22370 13376 22376 13388
rect 22331 13348 22376 13376
rect 22370 13336 22376 13348
rect 22428 13336 22434 13388
rect 20308 13311 20366 13317
rect 20308 13308 20320 13311
rect 18892 13280 19196 13308
rect 19996 13280 20320 13308
rect 12710 13240 12716 13252
rect 10468 13212 11100 13240
rect 12671 13212 12716 13240
rect 10468 13200 10474 13212
rect 12710 13200 12716 13212
rect 12768 13200 12774 13252
rect 17126 13200 17132 13252
rect 17184 13240 17190 13252
rect 17310 13240 17316 13252
rect 17184 13212 17316 13240
rect 17184 13200 17190 13212
rect 17310 13200 17316 13212
rect 17368 13200 17374 13252
rect 18892 13184 18920 13280
rect 5902 13132 5908 13184
rect 5960 13172 5966 13184
rect 6089 13175 6147 13181
rect 6089 13172 6101 13175
rect 5960 13144 6101 13172
rect 5960 13132 5966 13144
rect 6089 13141 6101 13144
rect 6135 13141 6147 13175
rect 6089 13135 6147 13141
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7009 13175 7067 13181
rect 7009 13172 7021 13175
rect 6972 13144 7021 13172
rect 6972 13132 6978 13144
rect 7009 13141 7021 13144
rect 7055 13141 7067 13175
rect 7009 13135 7067 13141
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 12805 13175 12863 13181
rect 10284 13144 10329 13172
rect 10284 13132 10290 13144
rect 12805 13141 12817 13175
rect 12851 13172 12863 13175
rect 14642 13172 14648 13184
rect 12851 13144 14648 13172
rect 12851 13141 12863 13144
rect 12805 13135 12863 13141
rect 14642 13132 14648 13144
rect 14700 13132 14706 13184
rect 15746 13172 15752 13184
rect 15659 13144 15752 13172
rect 15746 13132 15752 13144
rect 15804 13172 15810 13184
rect 16390 13172 16396 13184
rect 15804 13144 16396 13172
rect 15804 13132 15810 13144
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 18874 13172 18880 13184
rect 18835 13144 18880 13172
rect 18874 13132 18880 13144
rect 18932 13132 18938 13184
rect 19518 13132 19524 13184
rect 19576 13172 19582 13184
rect 19613 13175 19671 13181
rect 19613 13172 19625 13175
rect 19576 13144 19625 13172
rect 19576 13132 19582 13144
rect 19613 13141 19625 13144
rect 19659 13141 19671 13175
rect 19996 13172 20024 13280
rect 20308 13277 20320 13280
rect 20354 13277 20366 13311
rect 20308 13271 20366 13277
rect 20487 13311 20545 13317
rect 20487 13277 20499 13311
rect 20533 13277 20545 13311
rect 20487 13271 20545 13277
rect 20717 13311 20775 13317
rect 20717 13277 20729 13311
rect 20763 13308 20775 13311
rect 21082 13308 21088 13320
rect 20763 13280 21088 13308
rect 20763 13277 20775 13280
rect 20717 13271 20775 13277
rect 21082 13268 21088 13280
rect 21140 13308 21146 13320
rect 22020 13308 22048 13336
rect 22462 13308 22468 13320
rect 21140 13280 22048 13308
rect 22423 13280 22468 13308
rect 21140 13268 21146 13280
rect 22462 13268 22468 13280
rect 22520 13268 22526 13320
rect 22572 13317 22600 13484
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13277 22615 13311
rect 22830 13308 22836 13320
rect 22791 13280 22836 13308
rect 22557 13271 22615 13277
rect 22830 13268 22836 13280
rect 22888 13268 22894 13320
rect 22005 13243 22063 13249
rect 22005 13240 22017 13243
rect 21376 13212 22017 13240
rect 20438 13172 20444 13184
rect 19996 13144 20444 13172
rect 19613 13135 19671 13141
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 20806 13132 20812 13184
rect 20864 13172 20870 13184
rect 21376 13172 21404 13212
rect 22005 13209 22017 13212
rect 22051 13209 22063 13243
rect 22005 13203 22063 13209
rect 21818 13172 21824 13184
rect 20864 13144 21404 13172
rect 21779 13144 21824 13172
rect 20864 13132 20870 13144
rect 21818 13132 21824 13144
rect 21876 13132 21882 13184
rect 1104 13082 23460 13104
rect 1104 13030 4714 13082
rect 4766 13030 4778 13082
rect 4830 13030 4842 13082
rect 4894 13030 4906 13082
rect 4958 13030 12178 13082
rect 12230 13030 12242 13082
rect 12294 13030 12306 13082
rect 12358 13030 12370 13082
rect 12422 13030 19642 13082
rect 19694 13030 19706 13082
rect 19758 13030 19770 13082
rect 19822 13030 19834 13082
rect 19886 13030 23460 13082
rect 1104 13008 23460 13030
rect 3973 12971 4031 12977
rect 3973 12937 3985 12971
rect 4019 12968 4031 12971
rect 4338 12968 4344 12980
rect 4019 12940 4344 12968
rect 4019 12937 4031 12940
rect 3973 12931 4031 12937
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 5534 12968 5540 12980
rect 5495 12940 5540 12968
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 6457 12971 6515 12977
rect 6457 12937 6469 12971
rect 6503 12968 6515 12971
rect 6546 12968 6552 12980
rect 6503 12940 6552 12968
rect 6503 12937 6515 12940
rect 6457 12931 6515 12937
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 7926 12968 7932 12980
rect 7887 12940 7932 12968
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 10778 12968 10784 12980
rect 10739 12940 10784 12968
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 14737 12971 14795 12977
rect 14737 12937 14749 12971
rect 14783 12968 14795 12971
rect 14918 12968 14924 12980
rect 14783 12940 14924 12968
rect 14783 12937 14795 12940
rect 14737 12931 14795 12937
rect 14918 12928 14924 12940
rect 14976 12928 14982 12980
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 16485 12971 16543 12977
rect 16485 12968 16497 12971
rect 16080 12940 16497 12968
rect 16080 12928 16086 12940
rect 5442 12900 5448 12912
rect 5403 12872 5448 12900
rect 5442 12860 5448 12872
rect 5500 12900 5506 12912
rect 5500 12872 6040 12900
rect 5500 12860 5506 12872
rect 6012 12841 6040 12872
rect 9306 12860 9312 12912
rect 9364 12900 9370 12912
rect 9364 12872 11376 12900
rect 9364 12860 9370 12872
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6089 12835 6147 12841
rect 6089 12801 6101 12835
rect 6135 12832 6147 12835
rect 6730 12832 6736 12844
rect 6135 12804 6736 12832
rect 6135 12801 6147 12804
rect 6089 12795 6147 12801
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3878 12724 3884 12776
rect 3936 12764 3942 12776
rect 4065 12767 4123 12773
rect 4065 12764 4077 12767
rect 3936 12736 4077 12764
rect 3936 12724 3942 12736
rect 4065 12733 4077 12736
rect 4111 12764 4123 12767
rect 4614 12764 4620 12776
rect 4111 12736 4620 12764
rect 4111 12733 4123 12736
rect 4065 12727 4123 12733
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 5902 12764 5908 12776
rect 5863 12736 5908 12764
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 6104 12764 6132 12795
rect 6730 12792 6736 12804
rect 6788 12792 6794 12844
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12832 10103 12835
rect 10870 12832 10876 12844
rect 10091 12804 10876 12832
rect 10091 12801 10103 12804
rect 10045 12795 10103 12801
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11348 12841 11376 12872
rect 16224 12841 16252 12940
rect 16485 12937 16497 12940
rect 16531 12937 16543 12971
rect 16485 12931 16543 12937
rect 17770 12928 17776 12980
rect 17828 12968 17834 12980
rect 20162 12968 20168 12980
rect 17828 12940 20168 12968
rect 17828 12928 17834 12940
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20257 12971 20315 12977
rect 20257 12937 20269 12971
rect 20303 12968 20315 12971
rect 22554 12968 22560 12980
rect 20303 12940 22560 12968
rect 20303 12937 20315 12940
rect 20257 12931 20315 12937
rect 22554 12928 22560 12940
rect 22612 12928 22618 12980
rect 16500 12872 17264 12900
rect 16500 12844 16528 12872
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 13265 12835 13323 12841
rect 13265 12801 13277 12835
rect 13311 12832 13323 12835
rect 16209 12835 16267 12841
rect 13311 12804 13492 12832
rect 13311 12801 13323 12804
rect 13265 12795 13323 12801
rect 13464 12776 13492 12804
rect 16209 12801 16221 12835
rect 16255 12801 16267 12835
rect 16209 12795 16267 12801
rect 16482 12792 16488 12844
rect 16540 12792 16546 12844
rect 17126 12832 17132 12844
rect 17087 12804 17132 12832
rect 17126 12792 17132 12804
rect 17184 12792 17190 12844
rect 17236 12841 17264 12872
rect 19242 12860 19248 12912
rect 19300 12900 19306 12912
rect 20349 12903 20407 12909
rect 19300 12872 20300 12900
rect 19300 12860 19306 12872
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12801 17279 12835
rect 17221 12795 17279 12801
rect 19518 12792 19524 12844
rect 19576 12832 19582 12844
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 19576 12804 19809 12832
rect 19576 12792 19582 12804
rect 19797 12801 19809 12804
rect 19843 12801 19855 12835
rect 20272 12832 20300 12872
rect 20349 12869 20361 12903
rect 20395 12900 20407 12903
rect 20714 12900 20720 12912
rect 20395 12872 20720 12900
rect 20395 12869 20407 12872
rect 20349 12863 20407 12869
rect 20714 12860 20720 12872
rect 20772 12860 20778 12912
rect 22833 12903 22891 12909
rect 22833 12869 22845 12903
rect 22879 12900 22891 12903
rect 23474 12900 23480 12912
rect 22879 12872 23480 12900
rect 22879 12869 22891 12872
rect 22833 12863 22891 12869
rect 23474 12860 23480 12872
rect 23532 12860 23538 12912
rect 21910 12832 21916 12844
rect 20272 12804 20760 12832
rect 19797 12795 19855 12801
rect 6012 12736 6132 12764
rect 2860 12699 2918 12705
rect 2860 12665 2872 12699
rect 2906 12696 2918 12699
rect 3050 12696 3056 12708
rect 2906 12668 3056 12696
rect 2906 12665 2918 12668
rect 2860 12659 2918 12665
rect 3050 12656 3056 12668
rect 3108 12656 3114 12708
rect 4332 12699 4390 12705
rect 4332 12665 4344 12699
rect 4378 12696 4390 12699
rect 5258 12696 5264 12708
rect 4378 12668 5264 12696
rect 4378 12665 4390 12668
rect 4332 12659 4390 12665
rect 4246 12588 4252 12640
rect 4304 12628 4310 12640
rect 4347 12628 4375 12659
rect 5258 12656 5264 12668
rect 5316 12656 5322 12708
rect 4304 12600 4375 12628
rect 4304 12588 4310 12600
rect 4430 12588 4436 12640
rect 4488 12628 4494 12640
rect 6012 12628 6040 12736
rect 6638 12724 6644 12776
rect 6696 12764 6702 12776
rect 7570 12767 7628 12773
rect 7570 12764 7582 12767
rect 6696 12736 7582 12764
rect 6696 12724 6702 12736
rect 7570 12733 7582 12736
rect 7616 12733 7628 12767
rect 7570 12727 7628 12733
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 7282 12656 7288 12708
rect 7340 12696 7346 12708
rect 7852 12696 7880 12727
rect 8754 12724 8760 12776
rect 8812 12724 8818 12776
rect 9030 12724 9036 12776
rect 9088 12773 9094 12776
rect 9088 12764 9100 12773
rect 9309 12767 9367 12773
rect 9088 12736 9133 12764
rect 9088 12727 9100 12736
rect 9309 12733 9321 12767
rect 9355 12733 9367 12767
rect 11146 12764 11152 12776
rect 11107 12736 11152 12764
rect 9309 12727 9367 12733
rect 9088 12724 9094 12727
rect 8772 12696 8800 12724
rect 9324 12696 9352 12727
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 13354 12764 13360 12776
rect 13315 12736 13360 12764
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 13446 12724 13452 12776
rect 13504 12724 13510 12776
rect 15930 12764 15936 12776
rect 15988 12773 15994 12776
rect 14752 12736 15936 12764
rect 7340 12668 9352 12696
rect 13020 12699 13078 12705
rect 7340 12656 7346 12668
rect 13020 12665 13032 12699
rect 13066 12696 13078 12699
rect 13170 12696 13176 12708
rect 13066 12668 13176 12696
rect 13066 12665 13078 12668
rect 13020 12659 13078 12665
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 13624 12699 13682 12705
rect 13624 12665 13636 12699
rect 13670 12696 13682 12699
rect 14642 12696 14648 12708
rect 13670 12668 14648 12696
rect 13670 12665 13682 12668
rect 13624 12659 13682 12665
rect 14642 12656 14648 12668
rect 14700 12656 14706 12708
rect 4488 12600 6040 12628
rect 4488 12588 4494 12600
rect 8754 12588 8760 12640
rect 8812 12628 8818 12640
rect 9401 12631 9459 12637
rect 9401 12628 9413 12631
rect 8812 12600 9413 12628
rect 8812 12588 8818 12600
rect 9401 12597 9413 12600
rect 9447 12597 9459 12631
rect 9766 12628 9772 12640
rect 9727 12600 9772 12628
rect 9401 12591 9459 12597
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 9858 12588 9864 12640
rect 9916 12628 9922 12640
rect 9916 12600 9961 12628
rect 9916 12588 9922 12600
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 11885 12631 11943 12637
rect 11296 12600 11341 12628
rect 11296 12588 11302 12600
rect 11885 12597 11897 12631
rect 11931 12628 11943 12631
rect 14752 12628 14780 12736
rect 15930 12724 15936 12736
rect 15988 12727 16000 12773
rect 15988 12724 15994 12727
rect 16298 12724 16304 12776
rect 16356 12764 16362 12776
rect 16577 12767 16635 12773
rect 16356 12736 16401 12764
rect 16356 12724 16362 12736
rect 16577 12733 16589 12767
rect 16623 12764 16635 12767
rect 16623 12736 16657 12764
rect 16623 12733 16635 12736
rect 16577 12727 16635 12733
rect 16592 12696 16620 12727
rect 16758 12724 16764 12776
rect 16816 12764 16822 12776
rect 17313 12767 17371 12773
rect 17313 12764 17325 12767
rect 16816 12736 17325 12764
rect 16816 12724 16822 12736
rect 17313 12733 17325 12736
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 17773 12767 17831 12773
rect 17773 12764 17785 12767
rect 17552 12736 17785 12764
rect 17552 12724 17558 12736
rect 17773 12733 17785 12736
rect 17819 12733 17831 12767
rect 17773 12727 17831 12733
rect 18040 12767 18098 12773
rect 18040 12733 18052 12767
rect 18086 12764 18098 12767
rect 18874 12764 18880 12776
rect 18086 12736 18880 12764
rect 18086 12733 18098 12736
rect 18040 12727 18098 12733
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12733 20131 12767
rect 20073 12727 20131 12733
rect 17034 12696 17040 12708
rect 16408 12668 17040 12696
rect 11931 12600 14780 12628
rect 14829 12631 14887 12637
rect 11931 12597 11943 12600
rect 11885 12591 11943 12597
rect 14829 12597 14841 12631
rect 14875 12628 14887 12631
rect 15010 12628 15016 12640
rect 14875 12600 15016 12628
rect 14875 12597 14887 12600
rect 14829 12591 14887 12597
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 15746 12588 15752 12640
rect 15804 12628 15810 12640
rect 16408 12628 16436 12668
rect 17034 12656 17040 12668
rect 17092 12656 17098 12708
rect 17586 12696 17592 12708
rect 17144 12668 17592 12696
rect 15804 12600 16436 12628
rect 16761 12631 16819 12637
rect 15804 12588 15810 12600
rect 16761 12597 16773 12631
rect 16807 12628 16819 12631
rect 17144 12628 17172 12668
rect 17586 12656 17592 12668
rect 17644 12656 17650 12708
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 19705 12699 19763 12705
rect 19705 12696 19717 12699
rect 19484 12668 19717 12696
rect 19484 12656 19490 12668
rect 19705 12665 19717 12668
rect 19751 12696 19763 12699
rect 20088 12696 20116 12727
rect 19751 12668 20116 12696
rect 19751 12665 19763 12668
rect 19705 12659 19763 12665
rect 17678 12628 17684 12640
rect 16807 12600 17172 12628
rect 17639 12600 17684 12628
rect 16807 12597 16819 12600
rect 16761 12591 16819 12597
rect 17678 12588 17684 12600
rect 17736 12588 17742 12640
rect 19150 12628 19156 12640
rect 19111 12600 19156 12628
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 19242 12588 19248 12640
rect 19300 12628 19306 12640
rect 19610 12628 19616 12640
rect 19300 12600 19345 12628
rect 19571 12600 19616 12628
rect 19300 12588 19306 12600
rect 19610 12588 19616 12600
rect 19668 12588 19674 12640
rect 20732 12628 20760 12804
rect 21652 12804 21916 12832
rect 21652 12776 21680 12804
rect 21910 12792 21916 12804
rect 21968 12792 21974 12844
rect 22094 12792 22100 12844
rect 22152 12832 22158 12844
rect 22373 12835 22431 12841
rect 22373 12832 22385 12835
rect 22152 12804 22385 12832
rect 22152 12792 22158 12804
rect 22373 12801 22385 12804
rect 22419 12801 22431 12835
rect 22373 12795 22431 12801
rect 21473 12767 21531 12773
rect 21473 12733 21485 12767
rect 21519 12764 21531 12767
rect 21634 12764 21640 12776
rect 21519 12736 21640 12764
rect 21519 12733 21531 12736
rect 21473 12727 21531 12733
rect 21634 12724 21640 12736
rect 21692 12724 21698 12776
rect 21729 12767 21787 12773
rect 21729 12733 21741 12767
rect 21775 12733 21787 12767
rect 21729 12727 21787 12733
rect 21358 12656 21364 12708
rect 21416 12696 21422 12708
rect 21744 12696 21772 12727
rect 21416 12668 21772 12696
rect 22281 12699 22339 12705
rect 21416 12656 21422 12668
rect 22281 12665 22293 12699
rect 22327 12696 22339 12699
rect 22646 12696 22652 12708
rect 22327 12668 22652 12696
rect 22327 12665 22339 12668
rect 22281 12659 22339 12665
rect 22646 12656 22652 12668
rect 22704 12656 22710 12708
rect 21821 12631 21879 12637
rect 21821 12628 21833 12631
rect 20732 12600 21833 12628
rect 21821 12597 21833 12600
rect 21867 12597 21879 12631
rect 22370 12628 22376 12640
rect 22331 12600 22376 12628
rect 21821 12591 21879 12597
rect 22370 12588 22376 12600
rect 22428 12588 22434 12640
rect 1104 12538 23460 12560
rect 1104 12486 8446 12538
rect 8498 12486 8510 12538
rect 8562 12486 8574 12538
rect 8626 12486 8638 12538
rect 8690 12486 15910 12538
rect 15962 12486 15974 12538
rect 16026 12486 16038 12538
rect 16090 12486 16102 12538
rect 16154 12486 23460 12538
rect 1104 12464 23460 12486
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 3605 12427 3663 12433
rect 3605 12424 3617 12427
rect 3292 12396 3617 12424
rect 3292 12384 3298 12396
rect 3605 12393 3617 12396
rect 3651 12393 3663 12427
rect 4430 12424 4436 12436
rect 3605 12387 3663 12393
rect 3712 12396 4436 12424
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 3712 12356 3740 12396
rect 4430 12384 4436 12396
rect 4488 12384 4494 12436
rect 5258 12424 5264 12436
rect 5219 12396 5264 12424
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 6733 12427 6791 12433
rect 6733 12424 6745 12427
rect 6696 12396 6745 12424
rect 6696 12384 6702 12396
rect 6733 12393 6745 12396
rect 6779 12393 6791 12427
rect 6733 12387 6791 12393
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7374 12424 7380 12436
rect 6972 12396 7380 12424
rect 6972 12384 6978 12396
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 8297 12427 8355 12433
rect 8297 12424 8309 12427
rect 8076 12396 8309 12424
rect 8076 12384 8082 12396
rect 8297 12393 8309 12396
rect 8343 12424 8355 12427
rect 9401 12427 9459 12433
rect 9401 12424 9413 12427
rect 8343 12396 9413 12424
rect 8343 12393 8355 12396
rect 8297 12387 8355 12393
rect 9401 12393 9413 12396
rect 9447 12393 9459 12427
rect 9858 12424 9864 12436
rect 9819 12396 9864 12424
rect 9401 12387 9459 12393
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10229 12427 10287 12433
rect 10229 12393 10241 12427
rect 10275 12424 10287 12427
rect 10962 12424 10968 12436
rect 10275 12396 10968 12424
rect 10275 12393 10287 12396
rect 10229 12387 10287 12393
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 11238 12384 11244 12436
rect 11296 12424 11302 12436
rect 11974 12424 11980 12436
rect 11296 12396 11980 12424
rect 11296 12384 11302 12396
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 13725 12427 13783 12433
rect 13725 12424 13737 12427
rect 13688 12396 13737 12424
rect 13688 12384 13694 12396
rect 13725 12393 13737 12396
rect 13771 12424 13783 12427
rect 15746 12424 15752 12436
rect 13771 12396 15752 12424
rect 13771 12393 13783 12396
rect 13725 12387 13783 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 16669 12427 16727 12433
rect 16669 12393 16681 12427
rect 16715 12424 16727 12427
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 16715 12396 17877 12424
rect 16715 12393 16727 12396
rect 16669 12387 16727 12393
rect 17865 12393 17877 12396
rect 17911 12393 17923 12427
rect 17865 12387 17923 12393
rect 19153 12427 19211 12433
rect 19153 12393 19165 12427
rect 19199 12424 19211 12427
rect 19426 12424 19432 12436
rect 19199 12396 19432 12424
rect 19199 12393 19211 12396
rect 19153 12387 19211 12393
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 19610 12424 19616 12436
rect 19571 12396 19616 12424
rect 19610 12384 19616 12396
rect 19668 12384 19674 12436
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 2924 12328 3740 12356
rect 4148 12359 4206 12365
rect 2924 12316 2930 12328
rect 2976 12229 3004 12328
rect 4148 12325 4160 12359
rect 4194 12356 4206 12359
rect 4338 12356 4344 12368
rect 4194 12328 4344 12356
rect 4194 12325 4206 12328
rect 4148 12319 4206 12325
rect 4338 12316 4344 12328
rect 4396 12316 4402 12368
rect 5620 12359 5678 12365
rect 5620 12325 5632 12359
rect 5666 12356 5678 12359
rect 5902 12356 5908 12368
rect 5666 12328 5908 12356
rect 5666 12325 5678 12328
rect 5620 12319 5678 12325
rect 5902 12316 5908 12328
rect 5960 12316 5966 12368
rect 7184 12359 7242 12365
rect 7184 12325 7196 12359
rect 7230 12356 7242 12359
rect 7926 12356 7932 12368
rect 7230 12328 7932 12356
rect 7230 12325 7242 12328
rect 7184 12319 7242 12325
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 8846 12356 8852 12368
rect 8588 12328 8852 12356
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 3237 12291 3295 12297
rect 3237 12288 3249 12291
rect 3108 12260 3249 12288
rect 3108 12248 3114 12260
rect 3237 12257 3249 12260
rect 3283 12257 3295 12291
rect 3237 12251 3295 12257
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 8588 12297 8616 12328
rect 8846 12316 8852 12328
rect 8904 12316 8910 12368
rect 11054 12356 11060 12368
rect 9968 12328 11060 12356
rect 5353 12291 5411 12297
rect 5353 12288 5365 12291
rect 4672 12260 5365 12288
rect 4672 12248 4678 12260
rect 5353 12257 5365 12260
rect 5399 12257 5411 12291
rect 5353 12251 5411 12257
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12257 8631 12291
rect 8573 12251 8631 12257
rect 8665 12291 8723 12297
rect 8665 12257 8677 12291
rect 8711 12288 8723 12291
rect 8754 12288 8760 12300
rect 8711 12260 8760 12288
rect 8711 12257 8723 12260
rect 8665 12251 8723 12257
rect 8754 12248 8760 12260
rect 8812 12248 8818 12300
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 8864 12260 9505 12288
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12189 3019 12223
rect 3142 12220 3148 12232
rect 3103 12192 3148 12220
rect 2961 12183 3019 12189
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 3878 12220 3884 12232
rect 3839 12192 3884 12220
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 6914 12220 6920 12232
rect 6875 12192 6920 12220
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 7926 12180 7932 12232
rect 7984 12220 7990 12232
rect 8864 12220 8892 12260
rect 9493 12257 9505 12260
rect 9539 12257 9551 12291
rect 9493 12251 9551 12257
rect 7984 12192 8892 12220
rect 9309 12223 9367 12229
rect 7984 12180 7990 12192
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 9398 12220 9404 12232
rect 9355 12192 9404 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 8849 12155 8907 12161
rect 8849 12121 8861 12155
rect 8895 12152 8907 12155
rect 9968 12152 9996 12328
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 12066 12316 12072 12368
rect 12124 12356 12130 12368
rect 16114 12356 16120 12368
rect 12124 12328 16120 12356
rect 12124 12316 12130 12328
rect 16114 12316 16120 12328
rect 16172 12316 16178 12368
rect 17126 12316 17132 12368
rect 17184 12356 17190 12368
rect 17313 12359 17371 12365
rect 17313 12356 17325 12359
rect 17184 12328 17325 12356
rect 17184 12316 17190 12328
rect 17313 12325 17325 12328
rect 17359 12325 17371 12359
rect 18785 12359 18843 12365
rect 18785 12356 18797 12359
rect 17313 12319 17371 12325
rect 17420 12328 18797 12356
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10226 12288 10232 12300
rect 10091 12260 10232 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10226 12248 10232 12260
rect 10284 12248 10290 12300
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 10502 12288 10508 12300
rect 10367 12260 10508 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 10864 12291 10922 12297
rect 10864 12257 10876 12291
rect 10910 12288 10922 12291
rect 11238 12288 11244 12300
rect 10910 12260 11244 12288
rect 10910 12257 10922 12260
rect 10864 12251 10922 12257
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 12250 12288 12256 12300
rect 12211 12260 12256 12288
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 14734 12288 14740 12300
rect 13228 12260 14740 12288
rect 13228 12248 13234 12260
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 15194 12288 15200 12300
rect 15155 12260 15200 12288
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15470 12288 15476 12300
rect 15431 12260 15476 12288
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 15654 12248 15660 12300
rect 15712 12288 15718 12300
rect 16301 12291 16359 12297
rect 16301 12288 16313 12291
rect 15712 12260 16313 12288
rect 15712 12248 15718 12260
rect 16301 12257 16313 12260
rect 16347 12257 16359 12291
rect 17420 12288 17448 12328
rect 18785 12325 18797 12328
rect 18831 12325 18843 12359
rect 18785 12319 18843 12325
rect 16301 12251 16359 12257
rect 16500 12260 17448 12288
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 10597 12223 10655 12229
rect 10597 12220 10609 12223
rect 10468 12192 10609 12220
rect 10468 12180 10474 12192
rect 10597 12189 10609 12192
rect 10643 12189 10655 12223
rect 14826 12220 14832 12232
rect 14787 12192 14832 12220
rect 10597 12183 10655 12189
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15010 12220 15016 12232
rect 14971 12192 15016 12220
rect 15010 12180 15016 12192
rect 15068 12220 15074 12232
rect 16025 12223 16083 12229
rect 16025 12220 16037 12223
rect 15068 12192 16037 12220
rect 15068 12180 15074 12192
rect 16025 12189 16037 12192
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12220 16267 12223
rect 16390 12220 16396 12232
rect 16255 12192 16396 12220
rect 16255 12189 16267 12192
rect 16209 12183 16267 12189
rect 16390 12180 16396 12192
rect 16448 12180 16454 12232
rect 8895 12124 9996 12152
rect 8895 12121 8907 12124
rect 8849 12115 8907 12121
rect 13906 12112 13912 12164
rect 13964 12152 13970 12164
rect 15102 12152 15108 12164
rect 13964 12124 15108 12152
rect 13964 12112 13970 12124
rect 15102 12112 15108 12124
rect 15160 12112 15166 12164
rect 15381 12155 15439 12161
rect 15381 12121 15393 12155
rect 15427 12152 15439 12155
rect 16500 12152 16528 12260
rect 17586 12248 17592 12300
rect 17644 12288 17650 12300
rect 17957 12291 18015 12297
rect 17957 12288 17969 12291
rect 17644 12260 17969 12288
rect 17644 12248 17650 12260
rect 17957 12257 17969 12260
rect 18003 12257 18015 12291
rect 17957 12251 18015 12257
rect 18506 12248 18512 12300
rect 18564 12288 18570 12300
rect 19245 12291 19303 12297
rect 18564 12260 18828 12288
rect 18564 12248 18570 12260
rect 17218 12220 17224 12232
rect 17179 12192 17224 12220
rect 17218 12180 17224 12192
rect 17276 12180 17282 12232
rect 17402 12220 17408 12232
rect 17363 12192 17408 12220
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 17681 12223 17739 12229
rect 17681 12220 17693 12223
rect 17503 12192 17693 12220
rect 15427 12124 16528 12152
rect 15427 12121 15439 12124
rect 15381 12115 15439 12121
rect 16574 12112 16580 12164
rect 16632 12152 16638 12164
rect 16853 12155 16911 12161
rect 16853 12152 16865 12155
rect 16632 12124 16865 12152
rect 16632 12112 16638 12124
rect 16853 12121 16865 12124
rect 16899 12121 16911 12155
rect 16853 12115 16911 12121
rect 17126 12112 17132 12164
rect 17184 12152 17190 12164
rect 17503 12152 17531 12192
rect 17681 12189 17693 12192
rect 17727 12189 17739 12223
rect 17681 12183 17739 12189
rect 17770 12180 17776 12232
rect 17828 12180 17834 12232
rect 18616 12229 18644 12260
rect 18601 12223 18659 12229
rect 18601 12189 18613 12223
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18693 12223 18751 12229
rect 18693 12189 18705 12223
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 17788 12152 17816 12180
rect 17184 12124 17531 12152
rect 17604 12124 17816 12152
rect 17184 12112 17190 12124
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 8389 12087 8447 12093
rect 8389 12084 8401 12087
rect 8352 12056 8401 12084
rect 8352 12044 8358 12056
rect 8389 12053 8401 12056
rect 8435 12084 8447 12087
rect 8754 12084 8760 12096
rect 8435 12056 8760 12084
rect 8435 12053 8447 12056
rect 8389 12047 8447 12053
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 10505 12087 10563 12093
rect 10505 12053 10517 12087
rect 10551 12084 10563 12087
rect 11882 12084 11888 12096
rect 10551 12056 11888 12084
rect 10551 12053 10563 12056
rect 10505 12047 10563 12053
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 14366 12084 14372 12096
rect 14327 12056 14372 12084
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 15657 12087 15715 12093
rect 15657 12084 15669 12087
rect 15344 12056 15669 12084
rect 15344 12044 15350 12056
rect 15657 12053 15669 12056
rect 15703 12053 15715 12087
rect 15657 12047 15715 12053
rect 15841 12087 15899 12093
rect 15841 12053 15853 12087
rect 15887 12084 15899 12087
rect 16758 12084 16764 12096
rect 15887 12056 16764 12084
rect 15887 12053 15899 12056
rect 15841 12047 15899 12053
rect 16758 12044 16764 12056
rect 16816 12084 16822 12096
rect 17604 12084 17632 12124
rect 17954 12112 17960 12164
rect 18012 12152 18018 12164
rect 18708 12152 18736 12183
rect 18012 12124 18736 12152
rect 18800 12152 18828 12260
rect 19245 12257 19257 12291
rect 19291 12288 19303 12291
rect 19628 12288 19656 12384
rect 21450 12316 21456 12368
rect 21508 12356 21514 12368
rect 21508 12328 21864 12356
rect 21508 12316 21514 12328
rect 19291 12260 19656 12288
rect 19291 12257 19303 12260
rect 19245 12251 19303 12257
rect 20714 12248 20720 12300
rect 20772 12288 20778 12300
rect 21738 12291 21796 12297
rect 21738 12288 21750 12291
rect 20772 12260 21750 12288
rect 20772 12248 20778 12260
rect 21738 12257 21750 12260
rect 21784 12257 21796 12291
rect 21836 12288 21864 12328
rect 21910 12316 21916 12368
rect 21968 12356 21974 12368
rect 21968 12328 22600 12356
rect 21968 12316 21974 12328
rect 22572 12297 22600 12328
rect 22005 12291 22063 12297
rect 22005 12288 22017 12291
rect 21836 12260 22017 12288
rect 21738 12251 21796 12257
rect 22005 12257 22017 12260
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12257 22615 12291
rect 22738 12288 22744 12300
rect 22699 12260 22744 12288
rect 22557 12251 22615 12257
rect 22738 12248 22744 12260
rect 22796 12248 22802 12300
rect 22830 12248 22836 12300
rect 22888 12288 22894 12300
rect 22888 12260 22933 12288
rect 22888 12248 22894 12260
rect 19058 12180 19064 12232
rect 19116 12220 19122 12232
rect 20073 12223 20131 12229
rect 20073 12220 20085 12223
rect 19116 12192 20085 12220
rect 19116 12180 19122 12192
rect 20073 12189 20085 12192
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12189 20223 12223
rect 20165 12183 20223 12189
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12189 22155 12223
rect 22097 12183 22155 12189
rect 20180 12152 20208 12183
rect 18800 12124 20208 12152
rect 18012 12112 18018 12124
rect 16816 12056 17632 12084
rect 16816 12044 16822 12056
rect 17770 12044 17776 12096
rect 17828 12084 17834 12096
rect 18325 12087 18383 12093
rect 18325 12084 18337 12087
rect 17828 12056 18337 12084
rect 17828 12044 17834 12056
rect 18325 12053 18337 12056
rect 18371 12053 18383 12087
rect 18325 12047 18383 12053
rect 19429 12087 19487 12093
rect 19429 12053 19441 12087
rect 19475 12084 19487 12087
rect 19518 12084 19524 12096
rect 19475 12056 19524 12084
rect 19475 12053 19487 12056
rect 19429 12047 19487 12053
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 19978 12044 19984 12096
rect 20036 12084 20042 12096
rect 20438 12084 20444 12096
rect 20036 12056 20444 12084
rect 20036 12044 20042 12056
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 20622 12084 20628 12096
rect 20583 12056 20628 12084
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 21358 12044 21364 12096
rect 21416 12084 21422 12096
rect 21726 12084 21732 12096
rect 21416 12056 21732 12084
rect 21416 12044 21422 12056
rect 21726 12044 21732 12056
rect 21784 12084 21790 12096
rect 22112 12084 22140 12183
rect 21784 12056 22140 12084
rect 21784 12044 21790 12056
rect 1104 11994 23460 12016
rect 1104 11942 4714 11994
rect 4766 11942 4778 11994
rect 4830 11942 4842 11994
rect 4894 11942 4906 11994
rect 4958 11942 12178 11994
rect 12230 11942 12242 11994
rect 12294 11942 12306 11994
rect 12358 11942 12370 11994
rect 12422 11942 19642 11994
rect 19694 11942 19706 11994
rect 19758 11942 19770 11994
rect 19822 11942 19834 11994
rect 19886 11942 23460 11994
rect 1104 11920 23460 11942
rect 3050 11840 3056 11892
rect 3108 11880 3114 11892
rect 3421 11883 3479 11889
rect 3421 11880 3433 11883
rect 3108 11852 3433 11880
rect 3108 11840 3114 11852
rect 3421 11849 3433 11852
rect 3467 11849 3479 11883
rect 3421 11843 3479 11849
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 10502 11880 10508 11892
rect 4120 11852 10508 11880
rect 4120 11840 4126 11852
rect 10502 11840 10508 11852
rect 10560 11840 10566 11892
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 10873 11883 10931 11889
rect 10873 11880 10885 11883
rect 10652 11852 10885 11880
rect 10652 11840 10658 11852
rect 10873 11849 10885 11852
rect 10919 11849 10931 11883
rect 10873 11843 10931 11849
rect 11054 11840 11060 11892
rect 11112 11880 11118 11892
rect 12069 11883 12127 11889
rect 12069 11880 12081 11883
rect 11112 11852 12081 11880
rect 11112 11840 11118 11852
rect 12069 11849 12081 11852
rect 12115 11849 12127 11883
rect 12069 11843 12127 11849
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 15013 11883 15071 11889
rect 15013 11880 15025 11883
rect 14792 11852 15025 11880
rect 14792 11840 14798 11852
rect 15013 11849 15025 11852
rect 15059 11849 15071 11883
rect 15013 11843 15071 11849
rect 15102 11840 15108 11892
rect 15160 11880 15166 11892
rect 16022 11880 16028 11892
rect 15160 11852 16028 11880
rect 15160 11840 15166 11852
rect 16022 11840 16028 11852
rect 16080 11840 16086 11892
rect 16114 11840 16120 11892
rect 16172 11880 16178 11892
rect 17218 11880 17224 11892
rect 16172 11852 17224 11880
rect 16172 11840 16178 11852
rect 17218 11840 17224 11852
rect 17276 11840 17282 11892
rect 17681 11883 17739 11889
rect 17681 11849 17693 11883
rect 17727 11880 17739 11883
rect 17862 11880 17868 11892
rect 17727 11852 17868 11880
rect 17727 11849 17739 11852
rect 17681 11843 17739 11849
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 18046 11880 18052 11892
rect 18007 11852 18052 11880
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 20438 11880 20444 11892
rect 18432 11852 20444 11880
rect 3789 11815 3847 11821
rect 3789 11781 3801 11815
rect 3835 11812 3847 11815
rect 3878 11812 3884 11824
rect 3835 11784 3884 11812
rect 3835 11781 3847 11784
rect 3789 11775 3847 11781
rect 1394 11636 1400 11688
rect 1452 11676 1458 11688
rect 2041 11679 2099 11685
rect 2041 11676 2053 11679
rect 1452 11648 2053 11676
rect 1452 11636 1458 11648
rect 2041 11645 2053 11648
rect 2087 11676 2099 11679
rect 2590 11676 2596 11688
rect 2087 11648 2596 11676
rect 2087 11645 2099 11648
rect 2041 11639 2099 11645
rect 2590 11636 2596 11648
rect 2648 11676 2654 11688
rect 3804 11676 3832 11775
rect 3878 11772 3884 11784
rect 3936 11772 3942 11824
rect 10410 11772 10416 11824
rect 10468 11812 10474 11824
rect 11146 11812 11152 11824
rect 10468 11784 11152 11812
rect 10468 11772 10474 11784
rect 11146 11772 11152 11784
rect 11204 11812 11210 11824
rect 11204 11784 11249 11812
rect 11204 11772 11210 11784
rect 14826 11772 14832 11824
rect 14884 11812 14890 11824
rect 14921 11815 14979 11821
rect 14921 11812 14933 11815
rect 14884 11784 14933 11812
rect 14884 11772 14890 11784
rect 14921 11781 14933 11784
rect 14967 11781 14979 11815
rect 14921 11775 14979 11781
rect 16485 11815 16543 11821
rect 16485 11781 16497 11815
rect 16531 11812 16543 11815
rect 17954 11812 17960 11824
rect 16531 11784 17816 11812
rect 17915 11784 17960 11812
rect 16531 11781 16543 11784
rect 16485 11775 16543 11781
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 9784 11716 10241 11744
rect 2648 11648 3832 11676
rect 3973 11679 4031 11685
rect 2648 11636 2654 11648
rect 3973 11645 3985 11679
rect 4019 11645 4031 11679
rect 3973 11639 4031 11645
rect 2308 11611 2366 11617
rect 2308 11577 2320 11611
rect 2354 11608 2366 11611
rect 3142 11608 3148 11620
rect 2354 11580 3148 11608
rect 2354 11577 2366 11580
rect 2308 11571 2366 11577
rect 3142 11568 3148 11580
rect 3200 11568 3206 11620
rect 3988 11540 4016 11639
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 6972 11648 7021 11676
rect 6972 11636 6978 11648
rect 7009 11645 7021 11648
rect 7055 11676 7067 11679
rect 8202 11676 8208 11688
rect 7055 11648 8208 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 8202 11636 8208 11648
rect 8260 11676 8266 11688
rect 8573 11679 8631 11685
rect 8573 11676 8585 11679
rect 8260 11648 8585 11676
rect 8260 11636 8266 11648
rect 8573 11645 8585 11648
rect 8619 11645 8631 11679
rect 8573 11639 8631 11645
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 9784 11676 9812 11716
rect 10229 11713 10241 11716
rect 10275 11713 10287 11747
rect 13446 11744 13452 11756
rect 13407 11716 13452 11744
rect 10229 11707 10287 11713
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 9456 11648 9812 11676
rect 9456 11636 9462 11648
rect 9858 11636 9864 11688
rect 9916 11676 9922 11688
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 9916 11648 10977 11676
rect 9916 11636 9922 11648
rect 10965 11645 10977 11648
rect 11011 11645 11023 11679
rect 10965 11639 11023 11645
rect 11974 11636 11980 11688
rect 12032 11676 12038 11688
rect 13182 11679 13240 11685
rect 13182 11676 13194 11679
rect 12032 11648 13194 11676
rect 12032 11636 12038 11648
rect 13182 11645 13194 11648
rect 13228 11645 13240 11679
rect 13182 11639 13240 11645
rect 13541 11679 13599 11685
rect 13541 11645 13553 11679
rect 13587 11676 13599 11679
rect 14550 11676 14556 11688
rect 13587 11648 14556 11676
rect 13587 11645 13599 11648
rect 13541 11639 13599 11645
rect 14550 11636 14556 11648
rect 14608 11636 14614 11688
rect 14936 11676 14964 11775
rect 17037 11747 17095 11753
rect 17037 11744 17049 11747
rect 16316 11716 17049 11744
rect 16316 11688 16344 11716
rect 17037 11713 17049 11716
rect 17083 11744 17095 11747
rect 17126 11744 17132 11756
rect 17083 11716 17132 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11744 17279 11747
rect 17678 11744 17684 11756
rect 17267 11716 17684 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 17678 11704 17684 11716
rect 17736 11704 17742 11756
rect 17788 11744 17816 11784
rect 17954 11772 17960 11784
rect 18012 11772 18018 11824
rect 18432 11744 18460 11852
rect 20438 11840 20444 11852
rect 20496 11840 20502 11892
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 20990 11880 20996 11892
rect 20772 11852 20996 11880
rect 20772 11840 20778 11852
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 22002 11880 22008 11892
rect 21963 11852 22008 11880
rect 22002 11840 22008 11852
rect 22060 11840 22066 11892
rect 22186 11880 22192 11892
rect 22147 11852 22192 11880
rect 22186 11840 22192 11852
rect 22244 11840 22250 11892
rect 17788 11716 18460 11744
rect 19352 11716 20300 11744
rect 16126 11679 16184 11685
rect 16126 11676 16138 11679
rect 14936 11648 16138 11676
rect 16126 11645 16138 11648
rect 16172 11645 16184 11679
rect 16126 11639 16184 11645
rect 16298 11636 16304 11688
rect 16356 11636 16362 11688
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11676 16451 11679
rect 16482 11676 16488 11688
rect 16439 11648 16488 11676
rect 16439 11645 16451 11648
rect 16393 11639 16451 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 16758 11676 16764 11688
rect 16719 11648 16764 11676
rect 16758 11636 16764 11648
rect 16816 11636 16822 11688
rect 16942 11636 16948 11688
rect 17000 11676 17006 11688
rect 17313 11679 17371 11685
rect 17313 11676 17325 11679
rect 17000 11648 17325 11676
rect 17000 11636 17006 11648
rect 17313 11645 17325 11648
rect 17359 11645 17371 11679
rect 17770 11676 17776 11688
rect 17731 11648 17776 11676
rect 17313 11639 17371 11645
rect 17770 11636 17776 11648
rect 17828 11636 17834 11688
rect 19150 11676 19156 11688
rect 19208 11685 19214 11688
rect 19208 11679 19231 11685
rect 19083 11648 19156 11676
rect 19150 11636 19156 11648
rect 19219 11676 19231 11679
rect 19352 11676 19380 11716
rect 19219 11648 19380 11676
rect 19219 11645 19231 11648
rect 19208 11639 19231 11645
rect 19208 11636 19214 11639
rect 19426 11636 19432 11688
rect 19484 11676 19490 11688
rect 20162 11676 20168 11688
rect 19484 11648 19529 11676
rect 20123 11648 20168 11676
rect 19484 11636 19490 11648
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 20272 11676 20300 11716
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 20628 11747 20686 11753
rect 20628 11744 20640 11747
rect 20496 11716 20640 11744
rect 20496 11704 20502 11716
rect 20628 11713 20640 11716
rect 20674 11713 20686 11747
rect 20898 11744 20904 11756
rect 20859 11716 20904 11744
rect 20628 11707 20686 11713
rect 20898 11704 20904 11716
rect 20956 11704 20962 11756
rect 22741 11747 22799 11753
rect 22741 11744 22753 11747
rect 22066 11716 22753 11744
rect 22066 11676 22094 11716
rect 22741 11713 22753 11716
rect 22787 11713 22799 11747
rect 22741 11707 22799 11713
rect 22554 11676 22560 11688
rect 20272 11648 22094 11676
rect 22515 11648 22560 11676
rect 22554 11636 22560 11648
rect 22612 11636 22618 11688
rect 6822 11568 6828 11620
rect 6880 11608 6886 11620
rect 7276 11611 7334 11617
rect 7276 11608 7288 11611
rect 6880 11580 7288 11608
rect 6880 11568 6886 11580
rect 7276 11577 7288 11580
rect 7322 11608 7334 11611
rect 7926 11608 7932 11620
rect 7322 11580 7932 11608
rect 7322 11577 7334 11580
rect 7276 11571 7334 11577
rect 7926 11568 7932 11580
rect 7984 11568 7990 11620
rect 8846 11617 8852 11620
rect 8840 11608 8852 11617
rect 8807 11580 8852 11608
rect 8840 11571 8852 11580
rect 8846 11568 8852 11571
rect 8904 11568 8910 11620
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 13630 11608 13636 11620
rect 8996 11580 10732 11608
rect 8996 11568 9002 11580
rect 7374 11540 7380 11552
rect 3988 11512 7380 11540
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 8352 11512 8401 11540
rect 8352 11500 8358 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 9950 11540 9956 11552
rect 9911 11512 9956 11540
rect 8389 11503 8447 11509
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 10410 11540 10416 11552
rect 10371 11512 10416 11540
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 10502 11500 10508 11552
rect 10560 11540 10566 11552
rect 10704 11540 10732 11580
rect 11256 11580 13636 11608
rect 11256 11540 11284 11580
rect 13630 11568 13636 11580
rect 13688 11568 13694 11620
rect 13808 11611 13866 11617
rect 13808 11577 13820 11611
rect 13854 11608 13866 11611
rect 14182 11608 14188 11620
rect 13854 11580 14188 11608
rect 13854 11577 13866 11580
rect 13808 11571 13866 11577
rect 14182 11568 14188 11580
rect 14240 11568 14246 11620
rect 14918 11568 14924 11620
rect 14976 11608 14982 11620
rect 19058 11608 19064 11620
rect 14976 11580 19064 11608
rect 14976 11568 14982 11580
rect 19058 11568 19064 11580
rect 19116 11568 19122 11620
rect 19334 11568 19340 11620
rect 19392 11608 19398 11620
rect 19521 11611 19579 11617
rect 19521 11608 19533 11611
rect 19392 11580 19533 11608
rect 19392 11568 19398 11580
rect 19521 11577 19533 11580
rect 19567 11577 19579 11611
rect 19521 11571 19579 11577
rect 10560 11512 10605 11540
rect 10704 11512 11284 11540
rect 10560 11500 10566 11512
rect 13538 11500 13544 11552
rect 13596 11540 13602 11552
rect 16485 11543 16543 11549
rect 16485 11540 16497 11543
rect 13596 11512 16497 11540
rect 13596 11500 13602 11512
rect 16485 11509 16497 11512
rect 16531 11509 16543 11543
rect 16485 11503 16543 11509
rect 16577 11543 16635 11549
rect 16577 11509 16589 11543
rect 16623 11540 16635 11543
rect 16758 11540 16764 11552
rect 16623 11512 16764 11540
rect 16623 11509 16635 11512
rect 16577 11503 16635 11509
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 17218 11500 17224 11552
rect 17276 11540 17282 11552
rect 19889 11543 19947 11549
rect 19889 11540 19901 11543
rect 17276 11512 19901 11540
rect 17276 11500 17282 11512
rect 19889 11509 19901 11512
rect 19935 11509 19947 11543
rect 19889 11503 19947 11509
rect 19978 11500 19984 11552
rect 20036 11540 20042 11552
rect 20631 11543 20689 11549
rect 20631 11540 20643 11543
rect 20036 11512 20643 11540
rect 20036 11500 20042 11512
rect 20631 11509 20643 11512
rect 20677 11509 20689 11543
rect 22646 11540 22652 11552
rect 22607 11512 22652 11540
rect 20631 11503 20689 11509
rect 22646 11500 22652 11512
rect 22704 11500 22710 11552
rect 1104 11450 23460 11472
rect 1104 11398 8446 11450
rect 8498 11398 8510 11450
rect 8562 11398 8574 11450
rect 8626 11398 8638 11450
rect 8690 11398 15910 11450
rect 15962 11398 15974 11450
rect 16026 11398 16038 11450
rect 16090 11398 16102 11450
rect 16154 11398 23460 11450
rect 1104 11376 23460 11398
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 3142 11336 3148 11348
rect 2823 11308 3148 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 3142 11296 3148 11308
rect 3200 11296 3206 11348
rect 6822 11336 6828 11348
rect 6783 11308 6828 11336
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 8260 11308 8585 11336
rect 8260 11296 8266 11308
rect 8573 11305 8585 11308
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 9769 11339 9827 11345
rect 9769 11305 9781 11339
rect 9815 11336 9827 11339
rect 10502 11336 10508 11348
rect 9815 11308 10508 11336
rect 9815 11305 9827 11308
rect 9769 11299 9827 11305
rect 10502 11296 10508 11308
rect 10560 11296 10566 11348
rect 11238 11336 11244 11348
rect 11199 11308 11244 11336
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 14182 11336 14188 11348
rect 14143 11308 14188 11336
rect 14182 11296 14188 11308
rect 14240 11336 14246 11348
rect 14737 11339 14795 11345
rect 14737 11336 14749 11339
rect 14240 11308 14749 11336
rect 14240 11296 14246 11308
rect 14737 11305 14749 11308
rect 14783 11305 14795 11339
rect 16761 11339 16819 11345
rect 14737 11299 14795 11305
rect 15488 11308 16712 11336
rect 8018 11277 8024 11280
rect 7960 11271 8024 11277
rect 7960 11237 7972 11271
rect 8006 11237 8024 11271
rect 7960 11231 8024 11237
rect 8018 11228 8024 11231
rect 8076 11228 8082 11280
rect 10410 11228 10416 11280
rect 10468 11268 10474 11280
rect 10882 11271 10940 11277
rect 10882 11268 10894 11271
rect 10468 11240 10894 11268
rect 10468 11228 10474 11240
rect 10882 11237 10894 11240
rect 10928 11237 10940 11271
rect 15488 11268 15516 11308
rect 15654 11277 15660 11280
rect 15648 11268 15660 11277
rect 10882 11231 10940 11237
rect 10980 11240 15516 11268
rect 15615 11240 15660 11268
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 1670 11209 1676 11212
rect 1664 11163 1676 11209
rect 1728 11200 1734 11212
rect 1728 11172 1764 11200
rect 1670 11160 1676 11163
rect 1728 11160 1734 11172
rect 7374 11160 7380 11212
rect 7432 11200 7438 11212
rect 8757 11203 8815 11209
rect 8757 11200 8769 11203
rect 7432 11172 8769 11200
rect 7432 11160 7438 11172
rect 8757 11169 8769 11172
rect 8803 11169 8815 11203
rect 8757 11163 8815 11169
rect 9214 11160 9220 11212
rect 9272 11200 9278 11212
rect 10980 11200 11008 11240
rect 15648 11231 15660 11240
rect 15654 11228 15660 11231
rect 15712 11228 15718 11280
rect 16684 11268 16712 11308
rect 16761 11305 16773 11339
rect 16807 11336 16819 11339
rect 16850 11336 16856 11348
rect 16807 11308 16856 11336
rect 16807 11305 16819 11308
rect 16761 11299 16819 11305
rect 16850 11296 16856 11308
rect 16908 11336 16914 11348
rect 17129 11339 17187 11345
rect 17129 11336 17141 11339
rect 16908 11308 17141 11336
rect 16908 11296 16914 11308
rect 17129 11305 17141 11308
rect 17175 11305 17187 11339
rect 17586 11336 17592 11348
rect 17547 11308 17592 11336
rect 17129 11299 17187 11305
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 17957 11339 18015 11345
rect 17957 11305 17969 11339
rect 18003 11336 18015 11339
rect 22646 11336 22652 11348
rect 18003 11308 22652 11336
rect 18003 11305 18015 11308
rect 17957 11299 18015 11305
rect 22646 11296 22652 11308
rect 22704 11296 22710 11348
rect 16684 11240 17724 11268
rect 9272 11172 11008 11200
rect 9272 11160 9278 11172
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12354 11203 12412 11209
rect 12354 11200 12366 11203
rect 12124 11172 12366 11200
rect 12124 11160 12130 11172
rect 12354 11169 12366 11172
rect 12400 11169 12412 11203
rect 12354 11163 12412 11169
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13072 11203 13130 11209
rect 13072 11200 13084 11203
rect 12952 11172 13084 11200
rect 12952 11160 12958 11172
rect 13072 11169 13084 11172
rect 13118 11200 13130 11203
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 13118 11172 14841 11200
rect 13118 11169 13130 11172
rect 13072 11163 13130 11169
rect 14829 11169 14841 11172
rect 14875 11169 14887 11203
rect 14829 11163 14887 11169
rect 15028 11172 16436 11200
rect 15028 11144 15056 11172
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 8570 11132 8576 11144
rect 8251 11104 8576 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 11146 11132 11152 11144
rect 11107 11104 11152 11132
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11132 12679 11135
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12667 11104 12817 11132
rect 12667 11101 12679 11104
rect 12621 11095 12679 11101
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 15010 11132 15016 11144
rect 14971 11104 15016 11132
rect 12805 11095 12863 11101
rect 12820 10996 12848 11095
rect 15010 11092 15016 11104
rect 15068 11092 15074 11144
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11101 15439 11135
rect 16408 11132 16436 11172
rect 16482 11160 16488 11212
rect 16540 11200 16546 11212
rect 17221 11203 17279 11209
rect 17221 11200 17233 11203
rect 16540 11172 17233 11200
rect 16540 11160 16546 11172
rect 17221 11169 17233 11172
rect 17267 11169 17279 11203
rect 17221 11163 17279 11169
rect 16945 11135 17003 11141
rect 16945 11132 16957 11135
rect 16408 11104 16957 11132
rect 15381 11095 15439 11101
rect 16945 11101 16957 11104
rect 16991 11132 17003 11135
rect 17402 11132 17408 11144
rect 16991 11104 17408 11132
rect 16991 11101 17003 11104
rect 16945 11095 17003 11101
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 14369 11067 14427 11073
rect 14369 11064 14381 11067
rect 13872 11036 14381 11064
rect 13872 11024 13878 11036
rect 14369 11033 14381 11036
rect 14415 11033 14427 11067
rect 14369 11027 14427 11033
rect 14550 10996 14556 11008
rect 12820 10968 14556 10996
rect 14550 10956 14556 10968
rect 14608 10996 14614 11008
rect 15396 10996 15424 11095
rect 17402 11092 17408 11104
rect 17460 11092 17466 11144
rect 17696 11064 17724 11240
rect 18046 11228 18052 11280
rect 18104 11268 18110 11280
rect 18294 11271 18352 11277
rect 18294 11268 18306 11271
rect 18104 11240 18306 11268
rect 18104 11228 18110 11240
rect 18294 11237 18306 11240
rect 18340 11237 18352 11271
rect 18294 11231 18352 11237
rect 18690 11228 18696 11280
rect 18748 11268 18754 11280
rect 19150 11268 19156 11280
rect 18748 11240 19156 11268
rect 18748 11228 18754 11240
rect 19150 11228 19156 11240
rect 19208 11268 19214 11280
rect 20162 11268 20168 11280
rect 19208 11240 20168 11268
rect 19208 11228 19214 11240
rect 20162 11228 20168 11240
rect 20220 11228 20226 11280
rect 20622 11228 20628 11280
rect 20680 11268 20686 11280
rect 20910 11271 20968 11277
rect 20910 11268 20922 11271
rect 20680 11240 20922 11268
rect 20680 11228 20686 11240
rect 20910 11237 20922 11240
rect 20956 11237 20968 11271
rect 20910 11231 20968 11237
rect 21450 11228 21456 11280
rect 21508 11277 21514 11280
rect 21508 11271 21572 11277
rect 21508 11237 21526 11271
rect 21560 11237 21572 11271
rect 21508 11231 21572 11237
rect 21508 11228 21514 11231
rect 17773 11203 17831 11209
rect 17773 11169 17785 11203
rect 17819 11200 17831 11203
rect 19242 11200 19248 11212
rect 17819 11172 19248 11200
rect 17819 11169 17831 11172
rect 17773 11163 17831 11169
rect 19242 11160 19248 11172
rect 19300 11160 19306 11212
rect 20530 11160 20536 11212
rect 20588 11200 20594 11212
rect 21177 11203 21235 11209
rect 21177 11200 21189 11203
rect 20588 11172 21189 11200
rect 20588 11160 20594 11172
rect 21177 11169 21189 11172
rect 21223 11200 21235 11203
rect 21269 11203 21327 11209
rect 21269 11200 21281 11203
rect 21223 11172 21281 11200
rect 21223 11169 21235 11172
rect 21177 11163 21235 11169
rect 21269 11169 21281 11172
rect 21315 11169 21327 11203
rect 21269 11163 21327 11169
rect 18046 11132 18052 11144
rect 18007 11104 18052 11132
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 19392 11104 19625 11132
rect 19392 11092 19398 11104
rect 19613 11101 19625 11104
rect 19659 11132 19671 11135
rect 19978 11132 19984 11144
rect 19659 11104 19984 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 19978 11092 19984 11104
rect 20036 11092 20042 11144
rect 22554 11092 22560 11144
rect 22612 11132 22618 11144
rect 22741 11135 22799 11141
rect 22741 11132 22753 11135
rect 22612 11104 22753 11132
rect 22612 11092 22618 11104
rect 22741 11101 22753 11104
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 19797 11067 19855 11073
rect 19797 11064 19809 11067
rect 17696 11036 18092 11064
rect 16574 10996 16580 11008
rect 14608 10968 16580 10996
rect 14608 10956 14614 10968
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 18064 10996 18092 11036
rect 18984 11036 19809 11064
rect 18984 10996 19012 11036
rect 19797 11033 19809 11036
rect 19843 11064 19855 11067
rect 19843 11036 20300 11064
rect 19843 11033 19855 11036
rect 19797 11027 19855 11033
rect 18064 10968 19012 10996
rect 19429 10999 19487 11005
rect 19429 10965 19441 10999
rect 19475 10996 19487 10999
rect 19978 10996 19984 11008
rect 19475 10968 19984 10996
rect 19475 10965 19487 10968
rect 19429 10959 19487 10965
rect 19978 10956 19984 10968
rect 20036 10956 20042 11008
rect 20272 10996 20300 11036
rect 20990 10996 20996 11008
rect 20272 10968 20996 10996
rect 20990 10956 20996 10968
rect 21048 10956 21054 11008
rect 21910 10956 21916 11008
rect 21968 10996 21974 11008
rect 22649 10999 22707 11005
rect 22649 10996 22661 10999
rect 21968 10968 22661 10996
rect 21968 10956 21974 10968
rect 22649 10965 22661 10968
rect 22695 10996 22707 10999
rect 22738 10996 22744 11008
rect 22695 10968 22744 10996
rect 22695 10965 22707 10968
rect 22649 10959 22707 10965
rect 22738 10956 22744 10968
rect 22796 10956 22802 11008
rect 1104 10906 23460 10928
rect 1104 10854 4714 10906
rect 4766 10854 4778 10906
rect 4830 10854 4842 10906
rect 4894 10854 4906 10906
rect 4958 10854 12178 10906
rect 12230 10854 12242 10906
rect 12294 10854 12306 10906
rect 12358 10854 12370 10906
rect 12422 10854 19642 10906
rect 19694 10854 19706 10906
rect 19758 10854 19770 10906
rect 19822 10854 19834 10906
rect 19886 10854 23460 10906
rect 1104 10832 23460 10854
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9858 10792 9864 10804
rect 9171 10764 9864 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9858 10752 9864 10764
rect 9916 10752 9922 10804
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 10468 10764 10609 10792
rect 10468 10752 10474 10764
rect 10597 10761 10609 10764
rect 10643 10761 10655 10795
rect 11698 10792 11704 10804
rect 11659 10764 11704 10792
rect 10597 10755 10655 10761
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 12805 10795 12863 10801
rect 12805 10761 12817 10795
rect 12851 10792 12863 10795
rect 12894 10792 12900 10804
rect 12851 10764 12900 10792
rect 12851 10761 12863 10764
rect 12805 10755 12863 10761
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 15013 10795 15071 10801
rect 15013 10761 15025 10795
rect 15059 10792 15071 10795
rect 15654 10792 15660 10804
rect 15059 10764 15660 10792
rect 15059 10761 15071 10764
rect 15013 10755 15071 10761
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 16485 10795 16543 10801
rect 16485 10761 16497 10795
rect 16531 10792 16543 10795
rect 17494 10792 17500 10804
rect 16531 10764 17500 10792
rect 16531 10761 16543 10764
rect 16485 10755 16543 10761
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 19426 10792 19432 10804
rect 18708 10764 19432 10792
rect 16761 10727 16819 10733
rect 10796 10696 12296 10724
rect 8570 10656 8576 10668
rect 8483 10628 8576 10656
rect 8570 10616 8576 10628
rect 8628 10656 8634 10668
rect 8628 10628 9260 10656
rect 8628 10616 8634 10628
rect 9232 10600 9260 10628
rect 8294 10548 8300 10600
rect 8352 10597 8358 10600
rect 8352 10588 8364 10597
rect 8352 10560 8397 10588
rect 8352 10551 8364 10560
rect 8352 10548 8358 10551
rect 8754 10548 8760 10600
rect 8812 10588 8818 10600
rect 8941 10591 8999 10597
rect 8941 10588 8953 10591
rect 8812 10560 8953 10588
rect 8812 10548 8818 10560
rect 8941 10557 8953 10560
rect 8987 10557 8999 10591
rect 9214 10588 9220 10600
rect 9175 10560 9220 10588
rect 8941 10551 8999 10557
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9484 10591 9542 10597
rect 9484 10557 9496 10591
rect 9530 10588 9542 10591
rect 9950 10588 9956 10600
rect 9530 10560 9956 10588
rect 9530 10557 9542 10560
rect 9484 10551 9542 10557
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 9398 10480 9404 10532
rect 9456 10520 9462 10532
rect 10796 10529 10824 10696
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 12268 10665 12296 10696
rect 16761 10693 16773 10727
rect 16807 10693 16819 10727
rect 16761 10687 16819 10693
rect 12161 10659 12219 10665
rect 12161 10656 12173 10659
rect 12124 10628 12173 10656
rect 12124 10616 12130 10628
rect 12161 10625 12173 10628
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10625 12311 10659
rect 16666 10656 16672 10668
rect 12253 10619 12311 10625
rect 16316 10628 16672 10656
rect 11333 10591 11391 10597
rect 11333 10557 11345 10591
rect 11379 10588 11391 10591
rect 11422 10588 11428 10600
rect 11379 10560 11428 10588
rect 11379 10557 11391 10560
rect 11333 10551 11391 10557
rect 11422 10548 11428 10560
rect 11480 10548 11486 10600
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10588 14243 10591
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 14231 10560 14289 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10588 14611 10591
rect 14642 10588 14648 10600
rect 14599 10560 14648 10588
rect 14599 10557 14611 10560
rect 14553 10551 14611 10557
rect 14642 10548 14648 10560
rect 14700 10548 14706 10600
rect 14737 10591 14795 10597
rect 14737 10557 14749 10591
rect 14783 10588 14795 10591
rect 16316 10588 16344 10628
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 16776 10656 16804 10687
rect 18708 10665 18736 10764
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 22005 10795 22063 10801
rect 22005 10761 22017 10795
rect 22051 10792 22063 10795
rect 22370 10792 22376 10804
rect 22051 10764 22376 10792
rect 22051 10761 22063 10764
rect 22005 10755 22063 10761
rect 22370 10752 22376 10764
rect 22428 10752 22434 10804
rect 22833 10727 22891 10733
rect 22833 10693 22845 10727
rect 22879 10724 22891 10727
rect 23198 10724 23204 10736
rect 22879 10696 23204 10724
rect 22879 10693 22891 10696
rect 22833 10687 22891 10693
rect 23198 10684 23204 10696
rect 23256 10684 23262 10736
rect 18693 10659 18751 10665
rect 16776 10628 17448 10656
rect 14783 10560 16344 10588
rect 16393 10591 16451 10597
rect 14783 10557 14795 10560
rect 14737 10551 14795 10557
rect 16393 10557 16405 10591
rect 16439 10557 16451 10591
rect 16393 10551 16451 10557
rect 16577 10591 16635 10597
rect 16577 10557 16589 10591
rect 16623 10588 16635 10591
rect 17126 10588 17132 10600
rect 16623 10560 17132 10588
rect 16623 10557 16635 10560
rect 16577 10551 16635 10557
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 9456 10492 10793 10520
rect 9456 10480 9462 10492
rect 10781 10489 10793 10492
rect 10827 10489 10839 10523
rect 10781 10483 10839 10489
rect 11238 10480 11244 10532
rect 11296 10520 11302 10532
rect 12069 10523 12127 10529
rect 12069 10520 12081 10523
rect 11296 10492 12081 10520
rect 11296 10480 11302 10492
rect 12069 10489 12081 10492
rect 12115 10489 12127 10523
rect 12069 10483 12127 10489
rect 13940 10523 13998 10529
rect 13940 10489 13952 10523
rect 13986 10520 13998 10523
rect 15746 10520 15752 10532
rect 13986 10492 15752 10520
rect 13986 10489 13998 10492
rect 13940 10483 13998 10489
rect 15746 10480 15752 10492
rect 15804 10480 15810 10532
rect 16148 10523 16206 10529
rect 16148 10489 16160 10523
rect 16194 10520 16206 10523
rect 16298 10520 16304 10532
rect 16194 10492 16304 10520
rect 16194 10489 16206 10492
rect 16148 10483 16206 10489
rect 16298 10480 16304 10492
rect 16356 10480 16362 10532
rect 16408 10520 16436 10551
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 17218 10520 17224 10532
rect 16408 10492 17224 10520
rect 16592 10464 16620 10492
rect 17218 10480 17224 10492
rect 17276 10480 17282 10532
rect 17420 10520 17448 10628
rect 18693 10625 18705 10659
rect 18739 10625 18751 10659
rect 19426 10656 19432 10668
rect 18693 10619 18751 10625
rect 18800 10628 19432 10656
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 18064 10560 18429 10588
rect 18064 10532 18092 10560
rect 18417 10557 18429 10560
rect 18463 10588 18475 10591
rect 18800 10588 18828 10628
rect 19426 10616 19432 10628
rect 19484 10616 19490 10668
rect 19794 10665 19800 10668
rect 19751 10659 19800 10665
rect 19751 10625 19763 10659
rect 19797 10625 19800 10659
rect 19751 10619 19800 10625
rect 19794 10616 19800 10619
rect 19852 10616 19858 10668
rect 21450 10656 21456 10668
rect 21411 10628 21456 10656
rect 21450 10616 21456 10628
rect 21508 10616 21514 10668
rect 22186 10616 22192 10668
rect 22244 10656 22250 10668
rect 22462 10656 22468 10668
rect 22244 10628 22468 10656
rect 22244 10616 22250 10628
rect 22462 10616 22468 10628
rect 22520 10616 22526 10668
rect 18966 10588 18972 10600
rect 18463 10560 18828 10588
rect 18927 10560 18972 10588
rect 18463 10557 18475 10560
rect 18417 10551 18475 10557
rect 18966 10548 18972 10560
rect 19024 10548 19030 10600
rect 19150 10548 19156 10600
rect 19208 10588 19214 10600
rect 19245 10591 19303 10597
rect 19245 10588 19257 10591
rect 19208 10560 19257 10588
rect 19208 10548 19214 10560
rect 19245 10557 19257 10560
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 19978 10548 19984 10600
rect 20036 10588 20042 10600
rect 20036 10560 20081 10588
rect 20036 10548 20042 10560
rect 17420 10492 18000 10520
rect 7193 10455 7251 10461
rect 7193 10421 7205 10455
rect 7239 10452 7251 10455
rect 8754 10452 8760 10464
rect 7239 10424 8760 10452
rect 7239 10421 7251 10424
rect 7193 10415 7251 10421
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 14277 10455 14335 10461
rect 14277 10421 14289 10455
rect 14323 10452 14335 10455
rect 14369 10455 14427 10461
rect 14369 10452 14381 10455
rect 14323 10424 14381 10452
rect 14323 10421 14335 10424
rect 14277 10415 14335 10421
rect 14369 10421 14381 10424
rect 14415 10452 14427 10455
rect 14550 10452 14556 10464
rect 14415 10424 14556 10452
rect 14415 10421 14427 10424
rect 14369 10415 14427 10421
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 14921 10455 14979 10461
rect 14921 10421 14933 10455
rect 14967 10452 14979 10455
rect 16485 10455 16543 10461
rect 16485 10452 16497 10455
rect 14967 10424 16497 10452
rect 14967 10421 14979 10424
rect 14921 10415 14979 10421
rect 16485 10421 16497 10424
rect 16531 10421 16543 10455
rect 16485 10415 16543 10421
rect 16574 10412 16580 10464
rect 16632 10412 16638 10464
rect 17037 10455 17095 10461
rect 17037 10421 17049 10455
rect 17083 10452 17095 10455
rect 17494 10452 17500 10464
rect 17083 10424 17500 10452
rect 17083 10421 17095 10424
rect 17037 10415 17095 10421
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 17972 10452 18000 10492
rect 18046 10480 18052 10532
rect 18104 10480 18110 10532
rect 18172 10523 18230 10529
rect 18172 10489 18184 10523
rect 18218 10520 18230 10523
rect 21637 10523 21695 10529
rect 21637 10520 21649 10523
rect 18218 10492 19334 10520
rect 18218 10489 18230 10492
rect 18172 10483 18230 10489
rect 19306 10464 19334 10492
rect 20640 10492 21649 10520
rect 18506 10452 18512 10464
rect 17972 10424 18512 10452
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 18690 10412 18696 10464
rect 18748 10452 18754 10464
rect 18785 10455 18843 10461
rect 18785 10452 18797 10455
rect 18748 10424 18797 10452
rect 18748 10412 18754 10424
rect 18785 10421 18797 10424
rect 18831 10421 18843 10455
rect 18785 10415 18843 10421
rect 18874 10412 18880 10464
rect 18932 10452 18938 10464
rect 19153 10455 19211 10461
rect 19153 10452 19165 10455
rect 18932 10424 19165 10452
rect 18932 10412 18938 10424
rect 19153 10421 19165 10424
rect 19199 10421 19211 10455
rect 19306 10424 19340 10464
rect 19153 10415 19211 10421
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 19702 10412 19708 10464
rect 19760 10461 19766 10464
rect 19760 10452 19769 10461
rect 19760 10424 19805 10452
rect 19760 10415 19769 10424
rect 19760 10412 19766 10415
rect 19886 10412 19892 10464
rect 19944 10452 19950 10464
rect 20640 10452 20668 10492
rect 21637 10489 21649 10492
rect 21683 10489 21695 10523
rect 21637 10483 21695 10489
rect 22281 10523 22339 10529
rect 22281 10489 22293 10523
rect 22327 10520 22339 10523
rect 22462 10520 22468 10532
rect 22327 10492 22468 10520
rect 22327 10489 22339 10492
rect 22281 10483 22339 10489
rect 22462 10480 22468 10492
rect 22520 10480 22526 10532
rect 22557 10523 22615 10529
rect 22557 10489 22569 10523
rect 22603 10520 22615 10523
rect 22646 10520 22652 10532
rect 22603 10492 22652 10520
rect 22603 10489 22615 10492
rect 22557 10483 22615 10489
rect 22646 10480 22652 10492
rect 22704 10480 22710 10532
rect 19944 10424 20668 10452
rect 19944 10412 19950 10424
rect 20898 10412 20904 10464
rect 20956 10452 20962 10464
rect 21085 10455 21143 10461
rect 21085 10452 21097 10455
rect 20956 10424 21097 10452
rect 20956 10412 20962 10424
rect 21085 10421 21097 10424
rect 21131 10452 21143 10455
rect 21545 10455 21603 10461
rect 21545 10452 21557 10455
rect 21131 10424 21557 10452
rect 21131 10421 21143 10424
rect 21085 10415 21143 10421
rect 21545 10421 21557 10424
rect 21591 10421 21603 10455
rect 22370 10452 22376 10464
rect 22331 10424 22376 10452
rect 21545 10415 21603 10421
rect 22370 10412 22376 10424
rect 22428 10412 22434 10464
rect 1104 10362 23460 10384
rect 1104 10310 8446 10362
rect 8498 10310 8510 10362
rect 8562 10310 8574 10362
rect 8626 10310 8638 10362
rect 8690 10310 15910 10362
rect 15962 10310 15974 10362
rect 16026 10310 16038 10362
rect 16090 10310 16102 10362
rect 16154 10310 23460 10362
rect 1104 10288 23460 10310
rect 7561 10251 7619 10257
rect 7561 10217 7573 10251
rect 7607 10248 7619 10251
rect 8846 10248 8852 10260
rect 7607 10220 8852 10248
rect 7607 10217 7619 10220
rect 7561 10211 7619 10217
rect 8846 10208 8852 10220
rect 8904 10248 8910 10260
rect 9585 10251 9643 10257
rect 9585 10248 9597 10251
rect 8904 10220 9597 10248
rect 8904 10208 8910 10220
rect 9585 10217 9597 10220
rect 9631 10217 9643 10251
rect 9585 10211 9643 10217
rect 9677 10251 9735 10257
rect 9677 10217 9689 10251
rect 9723 10248 9735 10251
rect 9950 10248 9956 10260
rect 9723 10220 9956 10248
rect 9723 10217 9735 10220
rect 9677 10211 9735 10217
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 10045 10251 10103 10257
rect 10045 10217 10057 10251
rect 10091 10248 10103 10251
rect 10686 10248 10692 10260
rect 10091 10220 10692 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 11517 10251 11575 10257
rect 11517 10217 11529 10251
rect 11563 10248 11575 10251
rect 12066 10248 12072 10260
rect 11563 10220 12072 10248
rect 11563 10217 11575 10220
rect 11517 10211 11575 10217
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 15746 10248 15752 10260
rect 15659 10220 15752 10248
rect 15746 10208 15752 10220
rect 15804 10248 15810 10260
rect 16390 10248 16396 10260
rect 15804 10220 16396 10248
rect 15804 10208 15810 10220
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 18782 10248 18788 10260
rect 17144 10220 18788 10248
rect 8754 10189 8760 10192
rect 8696 10183 8760 10189
rect 8696 10149 8708 10183
rect 8742 10149 8760 10183
rect 8696 10143 8760 10149
rect 8754 10140 8760 10143
rect 8812 10140 8818 10192
rect 10404 10183 10462 10189
rect 10404 10149 10416 10183
rect 10450 10180 10462 10183
rect 10502 10180 10508 10192
rect 10450 10152 10508 10180
rect 10450 10149 10462 10152
rect 10404 10143 10462 10149
rect 10502 10140 10508 10152
rect 10560 10140 10566 10192
rect 13817 10183 13875 10189
rect 13817 10149 13829 10183
rect 13863 10180 13875 10183
rect 15286 10180 15292 10192
rect 13863 10152 15292 10180
rect 13863 10149 13875 10152
rect 13817 10143 13875 10149
rect 15286 10140 15292 10152
rect 15344 10140 15350 10192
rect 16850 10140 16856 10192
rect 16908 10189 16914 10192
rect 16908 10180 16920 10189
rect 16908 10152 16953 10180
rect 16908 10143 16920 10152
rect 16908 10140 16914 10143
rect 9214 10072 9220 10124
rect 9272 10112 9278 10124
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 9272 10084 10149 10112
rect 9272 10072 9278 10084
rect 10137 10081 10149 10084
rect 10183 10112 10195 10115
rect 11146 10112 11152 10124
rect 10183 10084 11152 10112
rect 10183 10081 10195 10084
rect 10137 10075 10195 10081
rect 11146 10072 11152 10084
rect 11204 10072 11210 10124
rect 12917 10115 12975 10121
rect 12917 10081 12929 10115
rect 12963 10112 12975 10115
rect 13446 10112 13452 10124
rect 12963 10084 13452 10112
rect 12963 10081 12975 10084
rect 12917 10075 12975 10081
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 13538 10072 13544 10124
rect 13596 10112 13602 10124
rect 14461 10115 14519 10121
rect 14461 10112 14473 10115
rect 13596 10084 14473 10112
rect 13596 10072 13602 10084
rect 14461 10081 14473 10084
rect 14507 10081 14519 10115
rect 14461 10075 14519 10081
rect 15013 10115 15071 10121
rect 15013 10081 15025 10115
rect 15059 10112 15071 10115
rect 17144 10112 17172 10220
rect 18782 10208 18788 10220
rect 18840 10208 18846 10260
rect 19245 10251 19303 10257
rect 19245 10217 19257 10251
rect 19291 10248 19303 10251
rect 19978 10248 19984 10260
rect 19291 10220 19984 10248
rect 19291 10217 19303 10220
rect 19245 10211 19303 10217
rect 19978 10208 19984 10220
rect 20036 10208 20042 10260
rect 21450 10208 21456 10260
rect 21508 10248 21514 10260
rect 22465 10251 22523 10257
rect 22465 10248 22477 10251
rect 21508 10220 22477 10248
rect 21508 10208 21514 10220
rect 22465 10217 22477 10220
rect 22511 10217 22523 10251
rect 22465 10211 22523 10217
rect 19426 10140 19432 10192
rect 19484 10180 19490 10192
rect 19610 10180 19616 10192
rect 19484 10152 19616 10180
rect 19484 10140 19490 10152
rect 19610 10140 19616 10152
rect 19668 10180 19674 10192
rect 19858 10183 19916 10189
rect 19858 10180 19870 10183
rect 19668 10152 19870 10180
rect 19668 10140 19674 10152
rect 19858 10149 19870 10152
rect 19904 10149 19916 10183
rect 19858 10143 19916 10149
rect 17402 10112 17408 10124
rect 15059 10084 17172 10112
rect 17363 10084 17408 10112
rect 15059 10081 15071 10084
rect 15013 10075 15071 10081
rect 17402 10072 17408 10084
rect 17460 10072 17466 10124
rect 20806 10112 20812 10124
rect 18064 10084 20812 10112
rect 8941 10047 8999 10053
rect 8941 10013 8953 10047
rect 8987 10044 8999 10047
rect 9398 10044 9404 10056
rect 8987 10016 9260 10044
rect 9359 10016 9404 10044
rect 8987 10013 8999 10016
rect 8941 10007 8999 10013
rect 9232 9976 9260 10016
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 13170 10044 13176 10056
rect 13131 10016 13176 10044
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10013 13691 10047
rect 13633 10007 13691 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 17129 10047 17187 10053
rect 13771 10016 14412 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 9674 9976 9680 9988
rect 9232 9948 9680 9976
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 13648 9976 13676 10007
rect 14090 9976 14096 9988
rect 13648 9948 14096 9976
rect 14090 9936 14096 9948
rect 14148 9936 14154 9988
rect 14384 9976 14412 10016
rect 17129 10013 17141 10047
rect 17175 10044 17187 10047
rect 17218 10044 17224 10056
rect 17175 10016 17224 10044
rect 17175 10013 17187 10016
rect 17129 10007 17187 10013
rect 17218 10004 17224 10016
rect 17276 10004 17282 10056
rect 17728 10047 17786 10053
rect 17728 10044 17740 10047
rect 17328 10016 17740 10044
rect 15470 9976 15476 9988
rect 14384 9948 15476 9976
rect 15470 9936 15476 9948
rect 15528 9936 15534 9988
rect 17328 9976 17356 10016
rect 17728 10013 17740 10016
rect 17774 10013 17786 10047
rect 17728 10007 17786 10013
rect 17911 10047 17969 10053
rect 17911 10013 17923 10047
rect 17957 10044 17969 10047
rect 18064 10044 18092 10084
rect 20806 10072 20812 10084
rect 20864 10072 20870 10124
rect 20898 10072 20904 10124
rect 20956 10112 20962 10124
rect 21341 10115 21399 10121
rect 21341 10112 21353 10115
rect 20956 10084 21353 10112
rect 20956 10072 20962 10084
rect 21341 10081 21353 10084
rect 21387 10081 21399 10115
rect 21341 10075 21399 10081
rect 23109 10115 23167 10121
rect 23109 10081 23121 10115
rect 23155 10112 23167 10115
rect 23290 10112 23296 10124
rect 23155 10084 23296 10112
rect 23155 10081 23167 10084
rect 23109 10075 23167 10081
rect 23290 10072 23296 10084
rect 23348 10072 23354 10124
rect 17957 10016 18092 10044
rect 18141 10047 18199 10053
rect 17957 10013 17969 10016
rect 17911 10007 17969 10013
rect 18141 10013 18153 10047
rect 18187 10044 18199 10047
rect 18322 10044 18328 10056
rect 18187 10016 18328 10044
rect 18187 10013 18199 10016
rect 18141 10007 18199 10013
rect 18322 10004 18328 10016
rect 18380 10004 18386 10056
rect 18506 10004 18512 10056
rect 18564 10044 18570 10056
rect 18564 10016 19564 10044
rect 18564 10004 18570 10016
rect 17144 9948 17356 9976
rect 11606 9868 11612 9920
rect 11664 9908 11670 9920
rect 11793 9911 11851 9917
rect 11793 9908 11805 9911
rect 11664 9880 11805 9908
rect 11664 9868 11670 9880
rect 11793 9877 11805 9880
rect 11839 9877 11851 9911
rect 11793 9871 11851 9877
rect 12066 9868 12072 9920
rect 12124 9908 12130 9920
rect 13906 9908 13912 9920
rect 12124 9880 13912 9908
rect 12124 9868 12130 9880
rect 13906 9868 13912 9880
rect 13964 9868 13970 9920
rect 14182 9908 14188 9920
rect 14143 9880 14188 9908
rect 14182 9868 14188 9880
rect 14240 9868 14246 9920
rect 15378 9868 15384 9920
rect 15436 9908 15442 9920
rect 15654 9908 15660 9920
rect 15436 9880 15660 9908
rect 15436 9868 15442 9880
rect 15654 9868 15660 9880
rect 15712 9908 15718 9920
rect 17144 9908 17172 9948
rect 15712 9880 17172 9908
rect 15712 9868 15718 9880
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 17313 9911 17371 9917
rect 17313 9908 17325 9911
rect 17276 9880 17325 9908
rect 17276 9868 17282 9880
rect 17313 9877 17325 9880
rect 17359 9908 17371 9911
rect 19242 9908 19248 9920
rect 17359 9880 19248 9908
rect 17359 9877 17371 9880
rect 17313 9871 17371 9877
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 19536 9908 19564 10016
rect 19610 10004 19616 10056
rect 19668 10044 19674 10056
rect 19668 10016 19713 10044
rect 19668 10004 19674 10016
rect 20622 10004 20628 10056
rect 20680 10044 20686 10056
rect 21085 10047 21143 10053
rect 21085 10044 21097 10047
rect 20680 10016 21097 10044
rect 20680 10004 20686 10016
rect 21085 10013 21097 10016
rect 21131 10013 21143 10047
rect 22830 10044 22836 10056
rect 22791 10016 22836 10044
rect 21085 10007 21143 10013
rect 22830 10004 22836 10016
rect 22888 10004 22894 10056
rect 20824 9948 21128 9976
rect 20824 9908 20852 9948
rect 19536 9880 20852 9908
rect 20898 9868 20904 9920
rect 20956 9908 20962 9920
rect 20993 9911 21051 9917
rect 20993 9908 21005 9911
rect 20956 9880 21005 9908
rect 20956 9868 20962 9880
rect 20993 9877 21005 9880
rect 21039 9877 21051 9911
rect 21100 9908 21128 9948
rect 21818 9908 21824 9920
rect 21100 9880 21824 9908
rect 20993 9871 21051 9877
rect 21818 9868 21824 9880
rect 21876 9868 21882 9920
rect 1104 9818 23460 9840
rect 1104 9766 4714 9818
rect 4766 9766 4778 9818
rect 4830 9766 4842 9818
rect 4894 9766 4906 9818
rect 4958 9766 12178 9818
rect 12230 9766 12242 9818
rect 12294 9766 12306 9818
rect 12358 9766 12370 9818
rect 12422 9766 19642 9818
rect 19694 9766 19706 9818
rect 19758 9766 19770 9818
rect 19822 9766 19834 9818
rect 19886 9766 23460 9818
rect 1104 9744 23460 9766
rect 13446 9704 13452 9716
rect 12268 9676 13452 9704
rect 8665 9639 8723 9645
rect 8665 9605 8677 9639
rect 8711 9636 8723 9639
rect 9766 9636 9772 9648
rect 8711 9608 9772 9636
rect 8711 9605 8723 9608
rect 8665 9599 8723 9605
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 11517 9639 11575 9645
rect 11517 9605 11529 9639
rect 11563 9636 11575 9639
rect 11701 9639 11759 9645
rect 11701 9636 11713 9639
rect 11563 9608 11713 9636
rect 11563 9605 11575 9608
rect 11517 9599 11575 9605
rect 11701 9605 11713 9608
rect 11747 9605 11759 9639
rect 11701 9599 11759 9605
rect 11793 9639 11851 9645
rect 11793 9605 11805 9639
rect 11839 9636 11851 9639
rect 12268 9636 12296 9676
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 14550 9704 14556 9716
rect 13556 9676 14556 9704
rect 13556 9636 13584 9676
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 16025 9707 16083 9713
rect 16025 9673 16037 9707
rect 16071 9704 16083 9707
rect 16298 9704 16304 9716
rect 16071 9676 16304 9704
rect 16071 9673 16083 9676
rect 16025 9667 16083 9673
rect 16298 9664 16304 9676
rect 16356 9664 16362 9716
rect 19334 9704 19340 9716
rect 16592 9676 19340 9704
rect 11839 9608 12296 9636
rect 13188 9608 13584 9636
rect 13633 9639 13691 9645
rect 11839 9605 11851 9608
rect 11793 9599 11851 9605
rect 13188 9580 13216 9608
rect 13633 9605 13645 9639
rect 13679 9636 13691 9639
rect 16482 9636 16488 9648
rect 13679 9608 14320 9636
rect 16443 9608 16488 9636
rect 13679 9605 13691 9608
rect 13633 9599 13691 9605
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9568 8263 9571
rect 8294 9568 8300 9580
rect 8251 9540 8300 9568
rect 8251 9537 8263 9540
rect 8205 9531 8263 9537
rect 8128 9500 8156 9531
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9568 11023 9571
rect 12066 9568 12072 9580
rect 11011 9540 12072 9568
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 12066 9528 12072 9540
rect 12124 9528 12130 9580
rect 13170 9568 13176 9580
rect 13131 9540 13176 9568
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 13814 9568 13820 9580
rect 13280 9540 13820 9568
rect 9398 9500 9404 9512
rect 8128 9472 9404 9500
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 9858 9500 9864 9512
rect 9819 9472 9864 9500
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9500 11207 9503
rect 11195 9472 12112 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 8297 9435 8355 9441
rect 8297 9401 8309 9435
rect 8343 9432 8355 9435
rect 8754 9432 8760 9444
rect 8343 9404 8760 9432
rect 8343 9401 8355 9404
rect 8297 9395 8355 9401
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 11701 9435 11759 9441
rect 11701 9401 11713 9435
rect 11747 9432 11759 9435
rect 12084 9432 12112 9472
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 13280 9500 13308 9540
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 13998 9568 14004 9580
rect 13959 9540 14004 9568
rect 13998 9528 14004 9540
rect 14056 9528 14062 9580
rect 14093 9571 14151 9577
rect 14093 9537 14105 9571
rect 14139 9568 14151 9571
rect 14182 9568 14188 9580
rect 14139 9540 14188 9568
rect 14139 9537 14151 9540
rect 14093 9531 14151 9537
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 14292 9568 14320 9608
rect 16482 9596 16488 9608
rect 16540 9596 16546 9648
rect 16209 9571 16267 9577
rect 14292 9540 14780 9568
rect 14366 9500 14372 9512
rect 12216 9472 13308 9500
rect 13372 9472 14372 9500
rect 12216 9460 12222 9472
rect 11747 9404 12020 9432
rect 12084 9404 12848 9432
rect 11747 9401 11759 9404
rect 11701 9395 11759 9401
rect 9674 9324 9680 9376
rect 9732 9364 9738 9376
rect 10045 9367 10103 9373
rect 10045 9364 10057 9367
rect 9732 9336 10057 9364
rect 9732 9324 9738 9336
rect 10045 9333 10057 9336
rect 10091 9333 10103 9367
rect 10045 9327 10103 9333
rect 11057 9367 11115 9373
rect 11057 9333 11069 9367
rect 11103 9364 11115 9367
rect 11882 9364 11888 9376
rect 11103 9336 11888 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 11992 9364 12020 9404
rect 12710 9364 12716 9376
rect 11992 9336 12716 9364
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 12820 9364 12848 9404
rect 12894 9392 12900 9444
rect 12952 9441 12958 9444
rect 12952 9432 12964 9441
rect 13372 9432 13400 9472
rect 14366 9460 14372 9472
rect 14424 9460 14430 9512
rect 14550 9460 14556 9512
rect 14608 9500 14614 9512
rect 14645 9503 14703 9509
rect 14645 9500 14657 9503
rect 14608 9472 14657 9500
rect 14608 9460 14614 9472
rect 14645 9469 14657 9472
rect 14691 9469 14703 9503
rect 14752 9500 14780 9540
rect 16209 9537 16221 9571
rect 16255 9568 16267 9571
rect 16592 9568 16620 9676
rect 19334 9664 19340 9676
rect 19392 9664 19398 9716
rect 22189 9707 22247 9713
rect 22189 9673 22201 9707
rect 22235 9704 22247 9707
rect 22370 9704 22376 9716
rect 22235 9676 22376 9704
rect 22235 9673 22247 9676
rect 22189 9667 22247 9673
rect 22370 9664 22376 9676
rect 22428 9664 22434 9716
rect 16761 9639 16819 9645
rect 16761 9605 16773 9639
rect 16807 9636 16819 9639
rect 16850 9636 16856 9648
rect 16807 9608 16856 9636
rect 16807 9605 16819 9608
rect 16761 9599 16819 9605
rect 16850 9596 16856 9608
rect 16908 9596 16914 9648
rect 18598 9636 18604 9648
rect 18559 9608 18604 9636
rect 18598 9596 18604 9608
rect 18656 9596 18662 9648
rect 19058 9636 19064 9648
rect 18708 9608 19064 9636
rect 16255 9540 16620 9568
rect 16255 9537 16267 9540
rect 16209 9531 16267 9537
rect 16298 9500 16304 9512
rect 14752 9472 16160 9500
rect 16259 9472 16304 9500
rect 14645 9463 14703 9469
rect 12952 9404 12997 9432
rect 13188 9404 13400 9432
rect 13449 9435 13507 9441
rect 12952 9395 12964 9404
rect 12952 9392 12958 9395
rect 13188 9364 13216 9404
rect 13449 9401 13461 9435
rect 13495 9432 13507 9435
rect 13633 9435 13691 9441
rect 13633 9432 13645 9435
rect 13495 9404 13645 9432
rect 13495 9401 13507 9404
rect 13449 9395 13507 9401
rect 13633 9401 13645 9404
rect 13679 9401 13691 9435
rect 13633 9395 13691 9401
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 14890 9435 14948 9441
rect 14890 9432 14902 9435
rect 14056 9404 14902 9432
rect 14056 9392 14062 9404
rect 14890 9401 14902 9404
rect 14936 9401 14948 9435
rect 16132 9432 16160 9472
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 16592 9509 16620 9540
rect 18414 9528 18420 9580
rect 18472 9568 18478 9580
rect 18708 9568 18736 9608
rect 19058 9596 19064 9608
rect 19116 9596 19122 9648
rect 21634 9596 21640 9648
rect 21692 9636 21698 9648
rect 22005 9639 22063 9645
rect 22005 9636 22017 9639
rect 21692 9608 22017 9636
rect 21692 9596 21698 9608
rect 22005 9605 22017 9608
rect 22051 9636 22063 9639
rect 23382 9636 23388 9648
rect 22051 9608 23388 9636
rect 22051 9605 22063 9608
rect 22005 9599 22063 9605
rect 23382 9596 23388 9608
rect 23440 9596 23446 9648
rect 18472 9540 18736 9568
rect 18472 9528 18478 9540
rect 18782 9528 18788 9580
rect 18840 9568 18846 9580
rect 19245 9571 19303 9577
rect 19245 9568 19257 9571
rect 18840 9540 19257 9568
rect 18840 9528 18846 9540
rect 19245 9537 19257 9540
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 19426 9528 19432 9580
rect 19484 9568 19490 9580
rect 19613 9571 19671 9577
rect 19613 9568 19625 9571
rect 19484 9540 19625 9568
rect 19484 9528 19490 9540
rect 19613 9537 19625 9540
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 19797 9571 19855 9577
rect 19797 9537 19809 9571
rect 19843 9568 19855 9571
rect 19978 9568 19984 9580
rect 19843 9540 19984 9568
rect 19843 9537 19855 9540
rect 19797 9531 19855 9537
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 22738 9568 22744 9580
rect 22699 9540 22744 9568
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 16577 9503 16635 9509
rect 16577 9469 16589 9503
rect 16623 9469 16635 9503
rect 16577 9463 16635 9469
rect 17034 9460 17040 9512
rect 17092 9500 17098 9512
rect 17129 9503 17187 9509
rect 17129 9500 17141 9503
rect 17092 9472 17141 9500
rect 17092 9460 17098 9472
rect 17129 9469 17141 9472
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 17221 9503 17279 9509
rect 17221 9469 17233 9503
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9500 19947 9503
rect 20070 9500 20076 9512
rect 19935 9472 20076 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 17227 9432 17255 9463
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 20622 9500 20628 9512
rect 20583 9472 20628 9500
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 22094 9500 22100 9512
rect 20824 9472 22100 9500
rect 17310 9432 17316 9444
rect 16132 9404 17080 9432
rect 17227 9404 17316 9432
rect 14890 9395 14948 9401
rect 12820 9336 13216 9364
rect 13357 9367 13415 9373
rect 13357 9333 13369 9367
rect 13403 9364 13415 9367
rect 13722 9364 13728 9376
rect 13403 9336 13728 9364
rect 13403 9333 13415 9336
rect 13357 9327 13415 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 14182 9364 14188 9376
rect 14143 9336 14188 9364
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 14553 9367 14611 9373
rect 14553 9333 14565 9367
rect 14599 9364 14611 9367
rect 15010 9364 15016 9376
rect 14599 9336 15016 9364
rect 14599 9333 14611 9336
rect 14553 9327 14611 9333
rect 15010 9324 15016 9336
rect 15068 9324 15074 9376
rect 16942 9364 16948 9376
rect 16903 9336 16948 9364
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 17052 9364 17080 9404
rect 17310 9392 17316 9404
rect 17368 9392 17374 9444
rect 17494 9441 17500 9444
rect 17488 9432 17500 9441
rect 17455 9404 17500 9432
rect 17488 9395 17500 9404
rect 17494 9392 17500 9395
rect 17552 9392 17558 9444
rect 17586 9392 17592 9444
rect 17644 9432 17650 9444
rect 18138 9432 18144 9444
rect 17644 9404 18144 9432
rect 17644 9392 17650 9404
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 19334 9392 19340 9444
rect 19392 9432 19398 9444
rect 20533 9435 20591 9441
rect 19392 9404 20392 9432
rect 19392 9392 19398 9404
rect 18414 9364 18420 9376
rect 17052 9336 18420 9364
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 18690 9364 18696 9376
rect 18651 9336 18696 9364
rect 18690 9324 18696 9336
rect 18748 9324 18754 9376
rect 19058 9364 19064 9376
rect 19019 9336 19064 9364
rect 19058 9324 19064 9336
rect 19116 9324 19122 9376
rect 19153 9367 19211 9373
rect 19153 9333 19165 9367
rect 19199 9364 19211 9367
rect 19426 9364 19432 9376
rect 19199 9336 19432 9364
rect 19199 9333 19211 9336
rect 19153 9327 19211 9333
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 20254 9364 20260 9376
rect 20215 9336 20260 9364
rect 20254 9324 20260 9336
rect 20312 9324 20318 9376
rect 20364 9364 20392 9404
rect 20533 9401 20545 9435
rect 20579 9432 20591 9435
rect 20824 9432 20852 9472
rect 22094 9460 22100 9472
rect 22152 9460 22158 9512
rect 20579 9404 20852 9432
rect 20892 9435 20950 9441
rect 20579 9401 20591 9404
rect 20533 9395 20591 9401
rect 20892 9401 20904 9435
rect 20938 9432 20950 9435
rect 20990 9432 20996 9444
rect 20938 9404 20996 9432
rect 20938 9401 20950 9404
rect 20892 9395 20950 9401
rect 20990 9392 20996 9404
rect 21048 9392 21054 9444
rect 21634 9392 21640 9444
rect 21692 9432 21698 9444
rect 22557 9435 22615 9441
rect 22557 9432 22569 9435
rect 21692 9404 22569 9432
rect 21692 9392 21698 9404
rect 22557 9401 22569 9404
rect 22603 9401 22615 9435
rect 22557 9395 22615 9401
rect 21542 9364 21548 9376
rect 20364 9336 21548 9364
rect 21542 9324 21548 9336
rect 21600 9324 21606 9376
rect 22094 9324 22100 9376
rect 22152 9364 22158 9376
rect 22649 9367 22707 9373
rect 22649 9364 22661 9367
rect 22152 9336 22661 9364
rect 22152 9324 22158 9336
rect 22649 9333 22661 9336
rect 22695 9333 22707 9367
rect 22649 9327 22707 9333
rect 23109 9367 23167 9373
rect 23109 9333 23121 9367
rect 23155 9364 23167 9367
rect 23290 9364 23296 9376
rect 23155 9336 23296 9364
rect 23155 9333 23167 9336
rect 23109 9327 23167 9333
rect 23290 9324 23296 9336
rect 23348 9324 23354 9376
rect 1104 9274 23460 9296
rect 1104 9222 8446 9274
rect 8498 9222 8510 9274
rect 8562 9222 8574 9274
rect 8626 9222 8638 9274
rect 8690 9222 15910 9274
rect 15962 9222 15974 9274
rect 16026 9222 16038 9274
rect 16090 9222 16102 9274
rect 16154 9222 23460 9274
rect 1104 9200 23460 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 1670 9160 1676 9172
rect 1627 9132 1676 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 13081 9163 13139 9169
rect 13081 9160 13093 9163
rect 12860 9132 13093 9160
rect 12860 9120 12866 9132
rect 13081 9129 13093 9132
rect 13127 9129 13139 9163
rect 13446 9160 13452 9172
rect 13407 9132 13452 9160
rect 13081 9123 13139 9129
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 13998 9120 14004 9172
rect 14056 9160 14062 9172
rect 14369 9163 14427 9169
rect 14369 9160 14381 9163
rect 14056 9132 14381 9160
rect 14056 9120 14062 9132
rect 14369 9129 14381 9132
rect 14415 9129 14427 9163
rect 14369 9123 14427 9129
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 19889 9163 19947 9169
rect 17552 9132 19748 9160
rect 17552 9120 17558 9132
rect 9674 9092 9680 9104
rect 9140 9064 9680 9092
rect 1394 9024 1400 9036
rect 1355 8996 1400 9024
rect 1394 8984 1400 8996
rect 1452 9024 1458 9036
rect 9140 9033 9168 9064
rect 9674 9052 9680 9064
rect 9732 9092 9738 9104
rect 9732 9064 11468 9092
rect 9732 9052 9738 9064
rect 1673 9027 1731 9033
rect 1673 9024 1685 9027
rect 1452 8996 1685 9024
rect 1452 8984 1458 8996
rect 1673 8993 1685 8996
rect 1719 8993 1731 9027
rect 1673 8987 1731 8993
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 9214 8984 9220 9036
rect 9272 9024 9278 9036
rect 9381 9027 9439 9033
rect 9381 9024 9393 9027
rect 9272 8996 9393 9024
rect 9272 8984 9278 8996
rect 9381 8993 9393 8996
rect 9427 8993 9439 9027
rect 9381 8987 9439 8993
rect 10965 9027 11023 9033
rect 10965 8993 10977 9027
rect 11011 9024 11023 9027
rect 11330 9024 11336 9036
rect 11011 8996 11336 9024
rect 11011 8993 11023 8996
rect 10965 8987 11023 8993
rect 11330 8984 11336 8996
rect 11388 8984 11394 9036
rect 11440 9024 11468 9064
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 13541 9095 13599 9101
rect 13541 9092 13553 9095
rect 11664 9064 13553 9092
rect 11664 9052 11670 9064
rect 13541 9061 13553 9064
rect 13587 9061 13599 9095
rect 13541 9055 13599 9061
rect 14090 9052 14096 9104
rect 14148 9092 14154 9104
rect 15482 9095 15540 9101
rect 15482 9092 15494 9095
rect 14148 9064 15494 9092
rect 14148 9052 14154 9064
rect 15482 9061 15494 9064
rect 15528 9061 15540 9095
rect 17712 9095 17770 9101
rect 15482 9055 15540 9061
rect 15764 9064 17080 9092
rect 15764 9036 15792 9064
rect 11701 9027 11759 9033
rect 11701 9024 11713 9027
rect 11440 8996 11713 9024
rect 11701 8993 11713 8996
rect 11747 8993 11759 9027
rect 11701 8987 11759 8993
rect 11968 9027 12026 9033
rect 11968 8993 11980 9027
rect 12014 9024 12026 9027
rect 12526 9024 12532 9036
rect 12014 8996 12532 9024
rect 12014 8993 12026 8996
rect 11968 8987 12026 8993
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 12710 8984 12716 9036
rect 12768 9024 12774 9036
rect 15194 9024 15200 9036
rect 12768 8996 15200 9024
rect 12768 8984 12774 8996
rect 15194 8984 15200 8996
rect 15252 8984 15258 9036
rect 15746 9024 15752 9036
rect 15659 8996 15752 9024
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 16025 9027 16083 9033
rect 16025 8993 16037 9027
rect 16071 9024 16083 9027
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 16071 8996 16497 9024
rect 16071 8993 16083 8996
rect 16025 8987 16083 8993
rect 16485 8993 16497 8996
rect 16531 9024 16543 9027
rect 16942 9024 16948 9036
rect 16531 8996 16948 9024
rect 16531 8993 16543 8996
rect 16485 8987 16543 8993
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17052 9024 17080 9064
rect 17712 9061 17724 9095
rect 17758 9092 17770 9095
rect 17954 9092 17960 9104
rect 17758 9064 17960 9092
rect 17758 9061 17770 9064
rect 17712 9055 17770 9061
rect 17954 9052 17960 9064
rect 18012 9052 18018 9104
rect 19334 9092 19340 9104
rect 18055 9064 19340 9092
rect 17052 8996 18000 9024
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8956 10931 8959
rect 11054 8956 11060 8968
rect 10919 8928 11060 8956
rect 10919 8925 10931 8928
rect 10873 8919 10931 8925
rect 10796 8888 10824 8919
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 12894 8916 12900 8968
rect 12952 8956 12958 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 12952 8928 13369 8956
rect 12952 8916 12958 8928
rect 13357 8925 13369 8928
rect 13403 8956 13415 8959
rect 13538 8956 13544 8968
rect 13403 8928 13544 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 17972 8965 18000 8996
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 13722 8888 13728 8900
rect 10796 8860 11560 8888
rect 10502 8820 10508 8832
rect 10463 8792 10508 8820
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 11333 8823 11391 8829
rect 11333 8789 11345 8823
rect 11379 8820 11391 8823
rect 11422 8820 11428 8832
rect 11379 8792 11428 8820
rect 11379 8789 11391 8792
rect 11333 8783 11391 8789
rect 11422 8780 11428 8792
rect 11480 8780 11486 8832
rect 11532 8820 11560 8860
rect 12912 8860 13728 8888
rect 12618 8820 12624 8832
rect 11532 8792 12624 8820
rect 12618 8780 12624 8792
rect 12676 8820 12682 8832
rect 12912 8820 12940 8860
rect 13722 8848 13728 8860
rect 13780 8848 13786 8900
rect 18055 8888 18083 9064
rect 19334 9052 19340 9064
rect 19392 9052 19398 9104
rect 18874 8984 18880 9036
rect 18932 9024 18938 9036
rect 19162 9027 19220 9033
rect 19162 9024 19174 9027
rect 18932 8996 19174 9024
rect 18932 8984 18938 8996
rect 19162 8993 19174 8996
rect 19208 8993 19220 9027
rect 19162 8987 19220 8993
rect 19720 8965 19748 9132
rect 19889 9129 19901 9163
rect 19935 9160 19947 9163
rect 20070 9160 20076 9172
rect 19935 9132 20076 9160
rect 19935 9129 19947 9132
rect 19889 9123 19947 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 20349 9163 20407 9169
rect 20349 9129 20361 9163
rect 20395 9160 20407 9163
rect 22186 9160 22192 9172
rect 20395 9132 22192 9160
rect 20395 9129 20407 9132
rect 20349 9123 20407 9129
rect 22186 9120 22192 9132
rect 22244 9120 22250 9172
rect 22462 9120 22468 9172
rect 22520 9160 22526 9172
rect 22925 9163 22983 9169
rect 22925 9160 22937 9163
rect 22520 9132 22937 9160
rect 22520 9120 22526 9132
rect 22925 9129 22937 9132
rect 22971 9129 22983 9163
rect 22925 9123 22983 9129
rect 20254 9052 20260 9104
rect 20312 9092 20318 9104
rect 20312 9064 21128 9092
rect 20312 9052 20318 9064
rect 19981 9027 20039 9033
rect 19981 8993 19993 9027
rect 20027 8993 20039 9027
rect 20898 9024 20904 9036
rect 20859 8996 20904 9024
rect 19981 8987 20039 8993
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8925 19763 8959
rect 19705 8919 19763 8925
rect 19444 8888 19472 8919
rect 19518 8888 19524 8900
rect 17972 8860 18083 8888
rect 19431 8860 19524 8888
rect 12676 8792 12940 8820
rect 12676 8780 12682 8792
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 13909 8823 13967 8829
rect 13909 8820 13921 8823
rect 13596 8792 13921 8820
rect 13596 8780 13602 8792
rect 13909 8789 13921 8792
rect 13955 8789 13967 8823
rect 13909 8783 13967 8789
rect 14642 8780 14648 8832
rect 14700 8820 14706 8832
rect 15841 8823 15899 8829
rect 15841 8820 15853 8823
rect 14700 8792 15853 8820
rect 14700 8780 14706 8792
rect 15841 8789 15853 8792
rect 15887 8789 15899 8823
rect 16298 8820 16304 8832
rect 16259 8792 16304 8820
rect 15841 8783 15899 8789
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 16574 8820 16580 8832
rect 16535 8792 16580 8820
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 17972 8820 18000 8860
rect 19518 8848 19524 8860
rect 19576 8888 19582 8900
rect 19886 8888 19892 8900
rect 19576 8860 19892 8888
rect 19576 8848 19582 8860
rect 19886 8848 19892 8860
rect 19944 8848 19950 8900
rect 16724 8792 18000 8820
rect 16724 8780 16730 8792
rect 18046 8780 18052 8832
rect 18104 8820 18110 8832
rect 18104 8792 18149 8820
rect 18104 8780 18110 8792
rect 18322 8780 18328 8832
rect 18380 8820 18386 8832
rect 19996 8820 20024 8987
rect 20898 8984 20904 8996
rect 20956 8984 20962 9036
rect 21100 9033 21128 9064
rect 21192 9064 21956 9092
rect 21192 9033 21220 9064
rect 21085 9027 21143 9033
rect 21085 8993 21097 9027
rect 21131 8993 21143 9027
rect 21085 8987 21143 8993
rect 21177 9027 21235 9033
rect 21177 8993 21189 9027
rect 21223 8993 21235 9027
rect 21809 9024 21815 9036
rect 21770 8996 21815 9024
rect 21177 8987 21235 8993
rect 21809 8984 21815 8996
rect 21867 8984 21873 9036
rect 21928 9024 21956 9064
rect 22554 9024 22560 9036
rect 21928 8996 22560 9024
rect 22554 8984 22560 8996
rect 22612 8984 22618 9036
rect 20441 8959 20499 8965
rect 20441 8925 20453 8959
rect 20487 8925 20499 8959
rect 20441 8919 20499 8925
rect 20254 8848 20260 8900
rect 20312 8888 20318 8900
rect 20456 8888 20484 8919
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 21545 8959 21603 8965
rect 21545 8956 21557 8959
rect 20680 8928 21557 8956
rect 20680 8916 20686 8928
rect 21545 8925 21557 8928
rect 21591 8925 21603 8959
rect 21545 8919 21603 8925
rect 21174 8888 21180 8900
rect 20312 8860 21180 8888
rect 20312 8848 20318 8860
rect 21174 8848 21180 8860
rect 21232 8848 21238 8900
rect 18380 8792 20024 8820
rect 18380 8780 18386 8792
rect 20530 8780 20536 8832
rect 20588 8820 20594 8832
rect 22462 8820 22468 8832
rect 20588 8792 22468 8820
rect 20588 8780 20594 8792
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 1104 8730 23460 8752
rect 1104 8678 4714 8730
rect 4766 8678 4778 8730
rect 4830 8678 4842 8730
rect 4894 8678 4906 8730
rect 4958 8678 12178 8730
rect 12230 8678 12242 8730
rect 12294 8678 12306 8730
rect 12358 8678 12370 8730
rect 12422 8678 19642 8730
rect 19694 8678 19706 8730
rect 19758 8678 19770 8730
rect 19822 8678 19834 8730
rect 19886 8678 23460 8730
rect 1104 8656 23460 8678
rect 1578 8576 1584 8628
rect 1636 8616 1642 8628
rect 1765 8619 1823 8625
rect 1765 8616 1777 8619
rect 1636 8588 1777 8616
rect 1636 8576 1642 8588
rect 1765 8585 1777 8588
rect 1811 8585 1823 8619
rect 1765 8579 1823 8585
rect 8849 8619 8907 8625
rect 8849 8585 8861 8619
rect 8895 8616 8907 8619
rect 9214 8616 9220 8628
rect 8895 8588 9220 8616
rect 8895 8585 8907 8588
rect 8849 8579 8907 8585
rect 9214 8576 9220 8588
rect 9272 8616 9278 8628
rect 11054 8616 11060 8628
rect 9272 8588 10640 8616
rect 11015 8588 11060 8616
rect 9272 8576 9278 8588
rect 10410 8480 10416 8492
rect 10371 8452 10416 8480
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10612 8489 10640 8588
rect 11054 8576 11060 8588
rect 11112 8576 11118 8628
rect 11517 8619 11575 8625
rect 11517 8585 11529 8619
rect 11563 8616 11575 8619
rect 13262 8616 13268 8628
rect 11563 8588 13268 8616
rect 11563 8585 11575 8588
rect 11517 8579 11575 8585
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 14090 8616 14096 8628
rect 14051 8588 14096 8616
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 18046 8616 18052 8628
rect 14568 8588 18052 8616
rect 14568 8548 14596 8588
rect 18046 8576 18052 8588
rect 18104 8616 18110 8628
rect 18782 8616 18788 8628
rect 18104 8588 18788 8616
rect 18104 8576 18110 8588
rect 18782 8576 18788 8588
rect 18840 8576 18846 8628
rect 21542 8576 21548 8628
rect 21600 8576 21606 8628
rect 21726 8576 21732 8628
rect 21784 8616 21790 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21784 8588 22017 8616
rect 21784 8576 21790 8588
rect 22005 8585 22017 8588
rect 22051 8616 22063 8619
rect 22738 8616 22744 8628
rect 22051 8588 22744 8616
rect 22051 8585 22063 8588
rect 22005 8579 22063 8585
rect 22738 8576 22744 8588
rect 22796 8576 22802 8628
rect 16574 8548 16580 8560
rect 14108 8520 14596 8548
rect 16132 8520 16580 8548
rect 10597 8483 10655 8489
rect 10597 8449 10609 8483
rect 10643 8449 10655 8483
rect 13722 8480 13728 8492
rect 13683 8452 13728 8480
rect 10597 8443 10655 8449
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8412 2007 8415
rect 2133 8415 2191 8421
rect 2133 8412 2145 8415
rect 1995 8384 2145 8412
rect 1995 8381 2007 8384
rect 1949 8375 2007 8381
rect 2133 8381 2145 8384
rect 2179 8412 2191 8415
rect 7374 8412 7380 8424
rect 2179 8384 7380 8412
rect 2179 8381 2191 8384
rect 2133 8375 2191 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 10229 8415 10287 8421
rect 10229 8412 10241 8415
rect 9732 8384 10241 8412
rect 9732 8372 9738 8384
rect 9876 8276 9904 8384
rect 10229 8381 10241 8384
rect 10275 8381 10287 8415
rect 10229 8375 10287 8381
rect 10502 8372 10508 8424
rect 10560 8412 10566 8424
rect 10689 8415 10747 8421
rect 10689 8412 10701 8415
rect 10560 8384 10701 8412
rect 10560 8372 10566 8384
rect 10689 8381 10701 8384
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 11333 8415 11391 8421
rect 11333 8381 11345 8415
rect 11379 8412 11391 8415
rect 13078 8412 13084 8424
rect 11379 8384 12572 8412
rect 13039 8384 13084 8412
rect 11379 8381 11391 8384
rect 11333 8375 11391 8381
rect 9984 8347 10042 8353
rect 9984 8313 9996 8347
rect 10030 8344 10042 8347
rect 11606 8344 11612 8356
rect 10030 8316 11612 8344
rect 10030 8313 10042 8316
rect 9984 8307 10042 8313
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 12434 8344 12440 8356
rect 11716 8316 12440 8344
rect 10778 8276 10784 8288
rect 9876 8248 10784 8276
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 11716 8285 11744 8316
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 11701 8279 11759 8285
rect 11701 8245 11713 8279
rect 11747 8245 11759 8279
rect 12544 8276 12572 8384
rect 13078 8372 13084 8384
rect 13136 8372 13142 8424
rect 13538 8412 13544 8424
rect 13499 8384 13544 8412
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 12836 8347 12894 8353
rect 12836 8313 12848 8347
rect 12882 8344 12894 8347
rect 14108 8344 14136 8520
rect 16132 8489 16160 8520
rect 16574 8508 16580 8520
rect 16632 8508 16638 8560
rect 16666 8508 16672 8560
rect 16724 8548 16730 8560
rect 16942 8548 16948 8560
rect 16724 8520 16769 8548
rect 16903 8520 16948 8548
rect 16724 8508 16730 8520
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 17221 8551 17279 8557
rect 17221 8517 17233 8551
rect 17267 8517 17279 8551
rect 17586 8548 17592 8560
rect 17221 8511 17279 8517
rect 17328 8520 17592 8548
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 15396 8452 16129 8480
rect 15217 8415 15275 8421
rect 15217 8381 15229 8415
rect 15263 8412 15275 8415
rect 15396 8412 15424 8452
rect 16117 8449 16129 8452
rect 16163 8449 16175 8483
rect 17236 8480 17264 8511
rect 16117 8443 16175 8449
rect 16224 8452 17264 8480
rect 15263 8384 15424 8412
rect 15473 8415 15531 8421
rect 15263 8381 15275 8384
rect 15217 8375 15275 8381
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 15746 8412 15752 8424
rect 15519 8384 15752 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 15746 8372 15752 8384
rect 15804 8372 15810 8424
rect 12882 8316 14136 8344
rect 12882 8313 12894 8316
rect 12836 8307 12894 8313
rect 14182 8304 14188 8356
rect 14240 8344 14246 8356
rect 16224 8353 16252 8452
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8412 17187 8415
rect 17328 8412 17356 8520
rect 17586 8508 17592 8520
rect 17644 8508 17650 8560
rect 18322 8548 18328 8560
rect 17696 8520 18328 8548
rect 17696 8489 17724 8520
rect 18322 8508 18328 8520
rect 18380 8508 18386 8560
rect 21560 8548 21588 8576
rect 21560 8520 22094 8548
rect 17681 8483 17739 8489
rect 17175 8384 17356 8412
rect 17420 8452 17632 8480
rect 17175 8381 17187 8384
rect 17129 8375 17187 8381
rect 15565 8347 15623 8353
rect 15565 8344 15577 8347
rect 14240 8316 15577 8344
rect 14240 8304 14246 8316
rect 15565 8313 15577 8316
rect 15611 8313 15623 8347
rect 15565 8307 15623 8313
rect 16209 8347 16267 8353
rect 16209 8313 16221 8347
rect 16255 8313 16267 8347
rect 16209 8307 16267 8313
rect 16393 8347 16451 8353
rect 16393 8313 16405 8347
rect 16439 8344 16451 8347
rect 17420 8344 17448 8452
rect 17604 8412 17632 8452
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8480 17923 8483
rect 17954 8480 17960 8492
rect 17911 8452 17960 8480
rect 17911 8449 17923 8452
rect 17865 8443 17923 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18288 8452 18644 8480
rect 18288 8440 18294 8452
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17604 8384 18061 8412
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 18138 8372 18144 8424
rect 18196 8412 18202 8424
rect 18325 8415 18383 8421
rect 18325 8412 18337 8415
rect 18196 8384 18337 8412
rect 18196 8372 18202 8384
rect 18325 8381 18337 8384
rect 18371 8381 18383 8415
rect 18616 8412 18644 8452
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 18788 8483 18846 8489
rect 18788 8480 18800 8483
rect 18748 8452 18800 8480
rect 18748 8440 18754 8452
rect 18788 8449 18800 8452
rect 18834 8449 18846 8483
rect 22066 8480 22094 8520
rect 22741 8483 22799 8489
rect 22741 8480 22753 8483
rect 22066 8452 22753 8480
rect 18788 8443 18846 8449
rect 22741 8449 22753 8452
rect 22787 8449 22799 8483
rect 22741 8443 22799 8449
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 18616 8384 19073 8412
rect 18325 8375 18383 8381
rect 19061 8381 19073 8384
rect 19107 8412 19119 8415
rect 19150 8412 19156 8424
rect 19107 8384 19156 8412
rect 19107 8381 19119 8384
rect 19061 8375 19119 8381
rect 19150 8372 19156 8384
rect 19208 8372 19214 8424
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 20622 8412 20628 8424
rect 20036 8384 20628 8412
rect 20036 8372 20042 8384
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 22370 8412 22376 8424
rect 20824 8384 22376 8412
rect 17586 8344 17592 8356
rect 16439 8316 17448 8344
rect 17547 8316 17592 8344
rect 16439 8313 16451 8316
rect 16393 8307 16451 8313
rect 17586 8304 17592 8316
rect 17644 8304 17650 8356
rect 20533 8347 20591 8353
rect 20533 8313 20545 8347
rect 20579 8344 20591 8347
rect 20824 8344 20852 8384
rect 22370 8372 22376 8384
rect 22428 8372 22434 8424
rect 20898 8353 20904 8356
rect 20579 8316 20852 8344
rect 20579 8313 20591 8316
rect 20533 8307 20591 8313
rect 20892 8307 20904 8353
rect 20956 8344 20962 8356
rect 22649 8347 22707 8353
rect 22649 8344 22661 8347
rect 20956 8316 20992 8344
rect 21100 8316 22661 8344
rect 20898 8304 20904 8307
rect 20956 8304 20962 8316
rect 13173 8279 13231 8285
rect 13173 8276 13185 8279
rect 12544 8248 13185 8276
rect 11701 8239 11759 8245
rect 13173 8245 13185 8248
rect 13219 8245 13231 8279
rect 13630 8276 13636 8288
rect 13591 8248 13636 8276
rect 13173 8239 13231 8245
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 15194 8236 15200 8288
rect 15252 8276 15258 8288
rect 15654 8276 15660 8288
rect 15252 8248 15660 8276
rect 15252 8236 15258 8248
rect 15654 8236 15660 8248
rect 15712 8276 15718 8288
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 15712 8248 15853 8276
rect 15712 8236 15718 8248
rect 15841 8245 15853 8248
rect 15887 8276 15899 8279
rect 16850 8276 16856 8288
rect 15887 8248 16856 8276
rect 15887 8245 15899 8248
rect 15841 8239 15899 8245
rect 16850 8236 16856 8248
rect 16908 8276 16914 8288
rect 18598 8276 18604 8288
rect 16908 8248 18604 8276
rect 16908 8236 16914 8248
rect 18598 8236 18604 8248
rect 18656 8276 18662 8288
rect 18791 8279 18849 8285
rect 18791 8276 18803 8279
rect 18656 8248 18803 8276
rect 18656 8236 18662 8248
rect 18791 8245 18803 8248
rect 18837 8245 18849 8279
rect 18791 8239 18849 8245
rect 20165 8279 20223 8285
rect 20165 8245 20177 8279
rect 20211 8276 20223 8279
rect 20622 8276 20628 8288
rect 20211 8248 20628 8276
rect 20211 8245 20223 8248
rect 20165 8239 20223 8245
rect 20622 8236 20628 8248
rect 20680 8276 20686 8288
rect 21100 8276 21128 8316
rect 22649 8313 22661 8316
rect 22695 8313 22707 8347
rect 22649 8307 22707 8313
rect 20680 8248 21128 8276
rect 20680 8236 20686 8248
rect 21266 8236 21272 8288
rect 21324 8276 21330 8288
rect 22094 8276 22100 8288
rect 21324 8248 22100 8276
rect 21324 8236 21330 8248
rect 22094 8236 22100 8248
rect 22152 8236 22158 8288
rect 22189 8279 22247 8285
rect 22189 8245 22201 8279
rect 22235 8276 22247 8279
rect 22462 8276 22468 8288
rect 22235 8248 22468 8276
rect 22235 8245 22247 8248
rect 22189 8239 22247 8245
rect 22462 8236 22468 8248
rect 22520 8236 22526 8288
rect 22554 8236 22560 8288
rect 22612 8276 22618 8288
rect 22612 8248 22657 8276
rect 22612 8236 22618 8248
rect 1104 8186 23460 8208
rect 1104 8134 8446 8186
rect 8498 8134 8510 8186
rect 8562 8134 8574 8186
rect 8626 8134 8638 8186
rect 8690 8134 15910 8186
rect 15962 8134 15974 8186
rect 16026 8134 16038 8186
rect 16090 8134 16102 8186
rect 16154 8134 23460 8186
rect 1104 8112 23460 8134
rect 9125 8075 9183 8081
rect 9125 8041 9137 8075
rect 9171 8072 9183 8075
rect 9398 8072 9404 8084
rect 9171 8044 9404 8072
rect 9171 8041 9183 8044
rect 9125 8035 9183 8041
rect 9398 8032 9404 8044
rect 9456 8072 9462 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 9456 8044 10885 8072
rect 9456 8032 9462 8044
rect 10873 8041 10885 8044
rect 10919 8041 10931 8075
rect 11330 8072 11336 8084
rect 11291 8044 11336 8072
rect 10873 8035 10931 8041
rect 11330 8032 11336 8044
rect 11388 8032 11394 8084
rect 11609 8075 11667 8081
rect 11609 8041 11621 8075
rect 11655 8041 11667 8075
rect 11609 8035 11667 8041
rect 10260 8007 10318 8013
rect 10260 7973 10272 8007
rect 10306 8004 10318 8007
rect 10502 8004 10508 8016
rect 10306 7976 10508 8004
rect 10306 7973 10318 7976
rect 10260 7967 10318 7973
rect 10502 7964 10508 7976
rect 10560 7964 10566 8016
rect 11624 8004 11652 8035
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 13262 8072 13268 8084
rect 12492 8044 12537 8072
rect 13223 8044 13268 8072
rect 12492 8032 12498 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 13725 8075 13783 8081
rect 13725 8041 13737 8075
rect 13771 8072 13783 8075
rect 14366 8072 14372 8084
rect 13771 8044 14372 8072
rect 13771 8041 13783 8044
rect 13725 8035 13783 8041
rect 14366 8032 14372 8044
rect 14424 8032 14430 8084
rect 16393 8075 16451 8081
rect 16393 8041 16405 8075
rect 16439 8072 16451 8075
rect 16439 8044 16620 8072
rect 16439 8041 16451 8044
rect 16393 8035 16451 8041
rect 13357 8007 13415 8013
rect 13357 8004 13369 8007
rect 11624 7976 13369 8004
rect 13357 7973 13369 7976
rect 13403 7973 13415 8007
rect 13357 7967 13415 7973
rect 13909 8007 13967 8013
rect 13909 7973 13921 8007
rect 13955 8004 13967 8007
rect 14461 8007 14519 8013
rect 14461 8004 14473 8007
rect 13955 7976 14473 8004
rect 13955 7973 13967 7976
rect 13909 7967 13967 7973
rect 14461 7973 14473 7976
rect 14507 7973 14519 8007
rect 14461 7967 14519 7973
rect 7374 7936 7380 7948
rect 7335 7908 7380 7936
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 8205 7939 8263 7945
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 8251 7908 10916 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 7392 7868 7420 7896
rect 8481 7871 8539 7877
rect 8481 7868 8493 7871
rect 7392 7840 8493 7868
rect 8481 7837 8493 7840
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 8496 7732 8524 7831
rect 10520 7800 10548 7831
rect 10594 7828 10600 7880
rect 10652 7868 10658 7880
rect 10689 7871 10747 7877
rect 10689 7868 10701 7871
rect 10652 7840 10701 7868
rect 10652 7828 10658 7840
rect 10689 7837 10701 7840
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 10778 7800 10784 7812
rect 10520 7772 10784 7800
rect 10778 7760 10784 7772
rect 10836 7760 10842 7812
rect 10888 7800 10916 7908
rect 10962 7896 10968 7948
rect 11020 7936 11026 7948
rect 11422 7936 11428 7948
rect 11020 7908 11065 7936
rect 11383 7908 11428 7936
rect 11020 7896 11026 7908
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7936 11943 7939
rect 11974 7936 11980 7948
rect 11931 7908 11980 7936
rect 11931 7905 11943 7908
rect 11885 7899 11943 7905
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7936 12587 7939
rect 12710 7936 12716 7948
rect 12575 7908 12716 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 12894 7896 12900 7948
rect 12952 7896 12958 7948
rect 13998 7936 14004 7948
rect 13959 7908 14004 7936
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 14476 7936 14504 7967
rect 14876 7939 14934 7945
rect 14876 7936 14888 7939
rect 14476 7908 14888 7936
rect 14876 7905 14888 7908
rect 14922 7936 14934 7939
rect 15194 7936 15200 7948
rect 14922 7908 15200 7936
rect 14922 7905 14934 7908
rect 14876 7899 14934 7905
rect 15194 7896 15200 7908
rect 15252 7896 15258 7948
rect 15286 7896 15292 7948
rect 15344 7936 15350 7948
rect 16592 7936 16620 8044
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 16951 8075 17009 8081
rect 16951 8072 16963 8075
rect 16908 8044 16963 8072
rect 16908 8032 16914 8044
rect 16951 8041 16963 8044
rect 16997 8041 17009 8075
rect 18322 8072 18328 8084
rect 18283 8044 18328 8072
rect 16951 8035 17009 8041
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 18601 8075 18659 8081
rect 18601 8041 18613 8075
rect 18647 8072 18659 8075
rect 19058 8072 19064 8084
rect 18647 8044 19064 8072
rect 18647 8041 18659 8044
rect 18601 8035 18659 8041
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 19426 8072 19432 8084
rect 19387 8044 19432 8072
rect 19426 8032 19432 8044
rect 19484 8032 19490 8084
rect 22554 8072 22560 8084
rect 19996 8044 22560 8072
rect 18969 8007 19027 8013
rect 18969 7973 18981 8007
rect 19015 8004 19027 8007
rect 19996 8004 20024 8044
rect 22554 8032 22560 8044
rect 22612 8032 22618 8084
rect 19015 7976 20024 8004
rect 19015 7973 19027 7976
rect 18969 7967 19027 7973
rect 21726 7964 21732 8016
rect 21784 8004 21790 8016
rect 21784 7976 22692 8004
rect 21784 7964 21790 7976
rect 17218 7936 17224 7948
rect 15344 7908 15389 7936
rect 16592 7908 17224 7936
rect 15344 7896 15350 7908
rect 17218 7896 17224 7908
rect 17276 7896 17282 7948
rect 17310 7896 17316 7948
rect 17368 7936 17374 7948
rect 19061 7939 19119 7945
rect 17368 7908 19012 7936
rect 17368 7896 17374 7908
rect 12345 7871 12403 7877
rect 12345 7837 12357 7871
rect 12391 7868 12403 7871
rect 12912 7868 12940 7896
rect 12391 7840 12940 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 12986 7828 12992 7880
rect 13044 7868 13050 7880
rect 13173 7871 13231 7877
rect 13173 7868 13185 7871
rect 13044 7840 13185 7868
rect 13044 7828 13050 7840
rect 13173 7837 13185 7840
rect 13219 7868 13231 7871
rect 14550 7868 14556 7880
rect 13219 7840 14320 7868
rect 14511 7840 14556 7868
rect 13219 7837 13231 7840
rect 13173 7831 13231 7837
rect 12897 7803 12955 7809
rect 10888 7772 12848 7800
rect 11882 7732 11888 7744
rect 8496 7704 11888 7732
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 12066 7732 12072 7744
rect 12027 7704 12072 7732
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 12820 7732 12848 7772
rect 12897 7769 12909 7803
rect 12943 7800 12955 7803
rect 13630 7800 13636 7812
rect 12943 7772 13636 7800
rect 12943 7769 12955 7772
rect 12897 7763 12955 7769
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 13909 7735 13967 7741
rect 13909 7732 13921 7735
rect 12820 7704 13921 7732
rect 13909 7701 13921 7704
rect 13955 7701 13967 7735
rect 14182 7732 14188 7744
rect 14143 7704 14188 7732
rect 13909 7695 13967 7701
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 14292 7732 14320 7840
rect 14550 7828 14556 7840
rect 14608 7828 14614 7880
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15068 7840 15113 7868
rect 15068 7828 15074 7840
rect 16482 7828 16488 7880
rect 16540 7868 16546 7880
rect 16991 7871 17049 7877
rect 16540 7840 16585 7868
rect 16540 7828 16546 7840
rect 16991 7837 17003 7871
rect 17037 7868 17049 7871
rect 17586 7868 17592 7880
rect 17037 7840 17592 7868
rect 17037 7837 17049 7840
rect 16991 7831 17049 7837
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 18874 7868 18880 7880
rect 18835 7840 18880 7868
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 18984 7868 19012 7908
rect 19061 7905 19073 7939
rect 19107 7936 19119 7939
rect 19150 7936 19156 7948
rect 19107 7908 19156 7936
rect 19107 7905 19119 7908
rect 19061 7899 19119 7905
rect 19150 7896 19156 7908
rect 19208 7896 19214 7948
rect 19797 7939 19855 7945
rect 19797 7905 19809 7939
rect 19843 7936 19855 7939
rect 19843 7908 21404 7936
rect 19843 7905 19855 7908
rect 19797 7899 19855 7905
rect 19702 7868 19708 7880
rect 18984 7840 19708 7868
rect 19702 7828 19708 7840
rect 19760 7828 19766 7880
rect 19889 7871 19947 7877
rect 19889 7837 19901 7871
rect 19935 7837 19947 7871
rect 19889 7831 19947 7837
rect 18138 7760 18144 7812
rect 18196 7800 18202 7812
rect 19242 7800 19248 7812
rect 18196 7772 19248 7800
rect 18196 7760 18202 7772
rect 19242 7760 19248 7772
rect 19300 7800 19306 7812
rect 19904 7800 19932 7831
rect 20070 7828 20076 7880
rect 20128 7868 20134 7880
rect 20438 7877 20444 7880
rect 20212 7871 20270 7877
rect 20212 7868 20224 7871
rect 20128 7840 20224 7868
rect 20128 7828 20134 7840
rect 20212 7837 20224 7840
rect 20258 7837 20270 7871
rect 20212 7831 20270 7837
rect 20395 7871 20444 7877
rect 20395 7837 20407 7871
rect 20441 7837 20444 7871
rect 20395 7831 20444 7837
rect 20438 7828 20444 7831
rect 20496 7828 20502 7880
rect 20622 7868 20628 7880
rect 20583 7840 20628 7868
rect 20622 7828 20628 7840
rect 20680 7828 20686 7880
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 21266 7868 21272 7880
rect 20864 7840 21272 7868
rect 20864 7828 20870 7840
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 21376 7868 21404 7908
rect 21818 7896 21824 7948
rect 21876 7936 21882 7948
rect 22462 7936 22468 7948
rect 21876 7908 21921 7936
rect 22423 7908 22468 7936
rect 21876 7896 21882 7908
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 22664 7945 22692 7976
rect 22649 7939 22707 7945
rect 22649 7905 22661 7939
rect 22695 7905 22707 7939
rect 22649 7899 22707 7905
rect 22370 7868 22376 7880
rect 21376 7840 22140 7868
rect 22331 7840 22376 7868
rect 19300 7772 19932 7800
rect 21284 7800 21312 7828
rect 21729 7803 21787 7809
rect 21729 7800 21741 7803
rect 21284 7772 21741 7800
rect 19300 7760 19306 7772
rect 21729 7769 21741 7772
rect 21775 7769 21787 7803
rect 22112 7800 22140 7840
rect 22370 7828 22376 7840
rect 22428 7828 22434 7880
rect 22922 7828 22928 7880
rect 22980 7868 22986 7880
rect 23109 7871 23167 7877
rect 23109 7868 23121 7871
rect 22980 7840 23121 7868
rect 22980 7828 22986 7840
rect 23109 7837 23121 7840
rect 23155 7837 23167 7871
rect 23109 7831 23167 7837
rect 22646 7800 22652 7812
rect 22112 7772 22652 7800
rect 21729 7763 21787 7769
rect 22646 7760 22652 7772
rect 22704 7760 22710 7812
rect 16942 7732 16948 7744
rect 14292 7704 16948 7732
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 18598 7692 18604 7744
rect 18656 7732 18662 7744
rect 19150 7732 19156 7744
rect 18656 7704 19156 7732
rect 18656 7692 18662 7704
rect 19150 7692 19156 7704
rect 19208 7732 19214 7744
rect 20070 7732 20076 7744
rect 19208 7704 20076 7732
rect 19208 7692 19214 7704
rect 20070 7692 20076 7704
rect 20128 7692 20134 7744
rect 20438 7692 20444 7744
rect 20496 7732 20502 7744
rect 21634 7732 21640 7744
rect 20496 7704 21640 7732
rect 20496 7692 20502 7704
rect 21634 7692 21640 7704
rect 21692 7732 21698 7744
rect 22005 7735 22063 7741
rect 22005 7732 22017 7735
rect 21692 7704 22017 7732
rect 21692 7692 21698 7704
rect 22005 7701 22017 7704
rect 22051 7701 22063 7735
rect 22005 7695 22063 7701
rect 1104 7642 23460 7664
rect 1104 7590 4714 7642
rect 4766 7590 4778 7642
rect 4830 7590 4842 7642
rect 4894 7590 4906 7642
rect 4958 7590 12178 7642
rect 12230 7590 12242 7642
rect 12294 7590 12306 7642
rect 12358 7590 12370 7642
rect 12422 7590 19642 7642
rect 19694 7590 19706 7642
rect 19758 7590 19770 7642
rect 19822 7590 19834 7642
rect 19886 7590 23460 7642
rect 1104 7568 23460 7590
rect 10502 7528 10508 7540
rect 10415 7500 10508 7528
rect 10502 7488 10508 7500
rect 10560 7528 10566 7540
rect 10962 7528 10968 7540
rect 10560 7500 10968 7528
rect 10560 7488 10566 7500
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11974 7528 11980 7540
rect 11935 7500 11980 7528
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 13998 7528 14004 7540
rect 13679 7500 14004 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 17586 7488 17592 7540
rect 17644 7528 17650 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 17644 7500 18061 7528
rect 17644 7488 17650 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 18049 7491 18107 7497
rect 18325 7531 18383 7537
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 18782 7528 18788 7540
rect 18371 7500 18788 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 20530 7528 20536 7540
rect 20364 7500 20536 7528
rect 11885 7463 11943 7469
rect 11885 7429 11897 7463
rect 11931 7460 11943 7463
rect 11931 7432 13124 7460
rect 11931 7429 11943 7432
rect 11885 7423 11943 7429
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7392 10839 7395
rect 12618 7392 12624 7404
rect 10827 7364 12624 7392
rect 10827 7361 10839 7364
rect 10781 7355 10839 7361
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 12986 7392 12992 7404
rect 12947 7364 12992 7392
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 13096 7401 13124 7432
rect 15488 7432 18276 7460
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7361 13139 7395
rect 14182 7392 14188 7404
rect 14143 7364 14188 7392
rect 13081 7355 13139 7361
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 14366 7392 14372 7404
rect 14327 7364 14372 7392
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7392 15163 7395
rect 15378 7392 15384 7404
rect 15151 7364 15384 7392
rect 15151 7361 15163 7364
rect 15105 7355 15163 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 9398 7333 9404 7336
rect 9125 7327 9183 7333
rect 9125 7293 9137 7327
rect 9171 7293 9183 7327
rect 9392 7324 9404 7333
rect 9359 7296 9404 7324
rect 9125 7287 9183 7293
rect 9392 7287 9404 7296
rect 9140 7256 9168 7287
rect 9398 7284 9404 7287
rect 9456 7284 9462 7336
rect 11701 7327 11759 7333
rect 11701 7324 11713 7327
rect 11348 7296 11713 7324
rect 9674 7256 9680 7268
rect 9140 7228 9680 7256
rect 9674 7216 9680 7228
rect 9732 7216 9738 7268
rect 10873 7259 10931 7265
rect 10873 7225 10885 7259
rect 10919 7256 10931 7259
rect 11146 7256 11152 7268
rect 10919 7228 11152 7256
rect 10919 7225 10931 7228
rect 10873 7219 10931 7225
rect 11146 7216 11152 7228
rect 11204 7216 11210 7268
rect 10965 7191 11023 7197
rect 10965 7157 10977 7191
rect 11011 7188 11023 7191
rect 11238 7188 11244 7200
rect 11011 7160 11244 7188
rect 11011 7157 11023 7160
rect 10965 7151 11023 7157
rect 11238 7148 11244 7160
rect 11296 7148 11302 7200
rect 11348 7197 11376 7296
rect 11701 7293 11713 7296
rect 11747 7293 11759 7327
rect 11701 7287 11759 7293
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 13173 7327 13231 7333
rect 13173 7324 13185 7327
rect 12124 7296 13185 7324
rect 12124 7284 12130 7296
rect 13173 7293 13185 7296
rect 13219 7293 13231 7327
rect 14461 7327 14519 7333
rect 14461 7324 14473 7327
rect 13173 7287 13231 7293
rect 13924 7296 14473 7324
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 12437 7259 12495 7265
rect 12437 7256 12449 7259
rect 12308 7228 12449 7256
rect 12308 7216 12314 7228
rect 12437 7225 12449 7228
rect 12483 7225 12495 7259
rect 13814 7256 13820 7268
rect 13775 7228 13820 7256
rect 12437 7219 12495 7225
rect 13814 7216 13820 7228
rect 13872 7216 13878 7268
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7157 11391 7191
rect 11333 7151 11391 7157
rect 12345 7191 12403 7197
rect 12345 7157 12357 7191
rect 12391 7188 12403 7191
rect 12986 7188 12992 7200
rect 12391 7160 12992 7188
rect 12391 7157 12403 7160
rect 12345 7151 12403 7157
rect 12986 7148 12992 7160
rect 13044 7148 13050 7200
rect 13541 7191 13599 7197
rect 13541 7157 13553 7191
rect 13587 7188 13599 7191
rect 13924 7188 13952 7296
rect 14461 7293 14473 7296
rect 14507 7324 14519 7327
rect 15488 7324 15516 7432
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 15838 7392 15844 7404
rect 15795 7364 15844 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 15838 7352 15844 7364
rect 15896 7352 15902 7404
rect 17126 7392 17132 7404
rect 16224 7364 17132 7392
rect 16224 7333 16252 7364
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 17218 7352 17224 7404
rect 17276 7392 17282 7404
rect 17405 7395 17463 7401
rect 17405 7392 17417 7395
rect 17276 7364 17417 7392
rect 17276 7352 17282 7364
rect 17405 7361 17417 7364
rect 17451 7361 17463 7395
rect 17586 7392 17592 7404
rect 17547 7364 17592 7392
rect 17405 7355 17463 7361
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 18248 7333 18276 7432
rect 20364 7392 20392 7500
rect 20530 7488 20536 7500
rect 20588 7488 20594 7540
rect 20990 7488 20996 7540
rect 21048 7528 21054 7540
rect 21726 7528 21732 7540
rect 21048 7500 21732 7528
rect 21048 7488 21054 7500
rect 21726 7488 21732 7500
rect 21784 7488 21790 7540
rect 22554 7488 22560 7540
rect 22612 7528 22618 7540
rect 22833 7531 22891 7537
rect 22833 7528 22845 7531
rect 22612 7500 22845 7528
rect 22612 7488 22618 7500
rect 22833 7497 22845 7500
rect 22879 7497 22891 7531
rect 22833 7491 22891 7497
rect 21634 7420 21640 7472
rect 21692 7460 21698 7472
rect 21821 7463 21879 7469
rect 21821 7460 21833 7463
rect 21692 7432 21833 7460
rect 21692 7420 21698 7432
rect 21821 7429 21833 7432
rect 21867 7429 21879 7463
rect 21821 7423 21879 7429
rect 22370 7392 22376 7404
rect 19628 7364 20392 7392
rect 22331 7364 22376 7392
rect 14507 7296 15516 7324
rect 16209 7327 16267 7333
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 16209 7293 16221 7327
rect 16255 7293 16267 7327
rect 16209 7287 16267 7293
rect 16393 7327 16451 7333
rect 16393 7293 16405 7327
rect 16439 7293 16451 7327
rect 16393 7287 16451 7293
rect 16485 7327 16543 7333
rect 16485 7293 16497 7327
rect 16531 7324 16543 7327
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 16531 7296 17785 7324
rect 16531 7293 16543 7296
rect 16485 7287 16543 7293
rect 17773 7293 17785 7296
rect 17819 7293 17831 7327
rect 17773 7287 17831 7293
rect 18233 7327 18291 7333
rect 18233 7293 18245 7327
rect 18279 7293 18291 7327
rect 18233 7287 18291 7293
rect 19449 7327 19507 7333
rect 19449 7293 19461 7327
rect 19495 7324 19507 7327
rect 19628 7324 19656 7364
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 19495 7296 19656 7324
rect 19705 7327 19763 7333
rect 19495 7293 19507 7296
rect 19449 7287 19507 7293
rect 19705 7293 19717 7327
rect 19751 7324 19763 7327
rect 19978 7324 19984 7336
rect 19751 7296 19984 7324
rect 19751 7293 19763 7296
rect 19705 7287 19763 7293
rect 14001 7259 14059 7265
rect 14001 7225 14013 7259
rect 14047 7256 14059 7259
rect 16408 7256 16436 7287
rect 14047 7228 15792 7256
rect 16408 7228 16988 7256
rect 14047 7225 14059 7228
rect 14001 7219 14059 7225
rect 13587 7160 13952 7188
rect 13587 7157 13599 7160
rect 13541 7151 13599 7157
rect 14550 7148 14556 7200
rect 14608 7188 14614 7200
rect 14829 7191 14887 7197
rect 14829 7188 14841 7191
rect 14608 7160 14841 7188
rect 14608 7148 14614 7160
rect 14829 7157 14841 7160
rect 14875 7157 14887 7191
rect 15194 7188 15200 7200
rect 15155 7160 15200 7188
rect 14829 7151 14887 7157
rect 15194 7148 15200 7160
rect 15252 7148 15258 7200
rect 15286 7148 15292 7200
rect 15344 7188 15350 7200
rect 15654 7188 15660 7200
rect 15344 7160 15389 7188
rect 15615 7160 15660 7188
rect 15344 7148 15350 7160
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 15764 7188 15792 7228
rect 16758 7188 16764 7200
rect 15764 7160 16764 7188
rect 16758 7148 16764 7160
rect 16816 7148 16822 7200
rect 16960 7197 16988 7228
rect 19610 7216 19616 7268
rect 19668 7256 19674 7268
rect 19720 7256 19748 7287
rect 19978 7284 19984 7296
rect 20036 7324 20042 7336
rect 20349 7327 20407 7333
rect 20349 7324 20361 7327
rect 20036 7296 20361 7324
rect 20036 7284 20042 7296
rect 20349 7293 20361 7296
rect 20395 7293 20407 7327
rect 20349 7287 20407 7293
rect 22005 7327 22063 7333
rect 22005 7293 22017 7327
rect 22051 7324 22063 7327
rect 22094 7324 22100 7336
rect 22051 7296 22100 7324
rect 22051 7293 22063 7296
rect 22005 7287 22063 7293
rect 22094 7284 22100 7296
rect 22152 7324 22158 7336
rect 23017 7327 23075 7333
rect 23017 7324 23029 7327
rect 22152 7296 23029 7324
rect 22152 7284 22158 7296
rect 23017 7293 23029 7296
rect 23063 7293 23075 7327
rect 23017 7287 23075 7293
rect 19668 7228 19748 7256
rect 19889 7259 19947 7265
rect 19668 7216 19674 7228
rect 19889 7225 19901 7259
rect 19935 7256 19947 7259
rect 20070 7256 20076 7268
rect 19935 7228 20076 7256
rect 19935 7225 19947 7228
rect 19889 7219 19947 7225
rect 20070 7216 20076 7228
rect 20128 7216 20134 7268
rect 20257 7259 20315 7265
rect 20257 7225 20269 7259
rect 20303 7256 20315 7259
rect 20438 7256 20444 7268
rect 20303 7228 20444 7256
rect 20303 7225 20315 7228
rect 20257 7219 20315 7225
rect 16945 7191 17003 7197
rect 16945 7157 16957 7191
rect 16991 7157 17003 7191
rect 17310 7188 17316 7200
rect 17271 7160 17316 7188
rect 16945 7151 17003 7157
rect 17310 7148 17316 7160
rect 17368 7148 17374 7200
rect 17402 7148 17408 7200
rect 17460 7188 17466 7200
rect 20272 7188 20300 7219
rect 20438 7216 20444 7228
rect 20496 7216 20502 7268
rect 20616 7259 20674 7265
rect 20616 7225 20628 7259
rect 20662 7225 20674 7259
rect 20616 7219 20674 7225
rect 17460 7160 20300 7188
rect 20640 7188 20668 7219
rect 20714 7216 20720 7268
rect 20772 7256 20778 7268
rect 20772 7228 21680 7256
rect 20772 7216 20778 7228
rect 20990 7188 20996 7200
rect 20640 7160 20996 7188
rect 17460 7148 17466 7160
rect 20990 7148 20996 7160
rect 21048 7188 21054 7200
rect 21542 7188 21548 7200
rect 21048 7160 21548 7188
rect 21048 7148 21054 7160
rect 21542 7148 21548 7160
rect 21600 7148 21606 7200
rect 21652 7188 21680 7228
rect 22186 7216 22192 7268
rect 22244 7256 22250 7268
rect 22281 7259 22339 7265
rect 22281 7256 22293 7259
rect 22244 7228 22293 7256
rect 22244 7216 22250 7228
rect 22281 7225 22293 7228
rect 22327 7225 22339 7259
rect 22281 7219 22339 7225
rect 22373 7191 22431 7197
rect 22373 7188 22385 7191
rect 21652 7160 22385 7188
rect 22373 7157 22385 7160
rect 22419 7157 22431 7191
rect 22373 7151 22431 7157
rect 1104 7098 23460 7120
rect 1104 7046 8446 7098
rect 8498 7046 8510 7098
rect 8562 7046 8574 7098
rect 8626 7046 8638 7098
rect 8690 7046 15910 7098
rect 15962 7046 15974 7098
rect 16026 7046 16038 7098
rect 16090 7046 16102 7098
rect 16154 7046 23460 7098
rect 1104 7024 23460 7046
rect 10042 6944 10048 6996
rect 10100 6984 10106 6996
rect 10965 6987 11023 6993
rect 10965 6984 10977 6987
rect 10100 6956 10977 6984
rect 10100 6944 10106 6956
rect 10965 6953 10977 6956
rect 11011 6953 11023 6987
rect 10965 6947 11023 6953
rect 11238 6944 11244 6996
rect 11296 6984 11302 6996
rect 11425 6987 11483 6993
rect 11425 6984 11437 6987
rect 11296 6956 11437 6984
rect 11296 6944 11302 6956
rect 11425 6953 11437 6956
rect 11471 6953 11483 6987
rect 12250 6984 12256 6996
rect 12211 6956 12256 6984
rect 11425 6947 11483 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 13081 6987 13139 6993
rect 13081 6984 13093 6987
rect 13044 6956 13093 6984
rect 13044 6944 13050 6956
rect 13081 6953 13093 6956
rect 13127 6953 13139 6987
rect 13081 6947 13139 6953
rect 17221 6987 17279 6993
rect 17221 6953 17233 6987
rect 17267 6953 17279 6987
rect 17221 6947 17279 6953
rect 20441 6987 20499 6993
rect 20441 6953 20453 6987
rect 20487 6984 20499 6987
rect 20898 6984 20904 6996
rect 20487 6956 20904 6984
rect 20487 6953 20499 6956
rect 20441 6947 20499 6953
rect 10260 6919 10318 6925
rect 10260 6885 10272 6919
rect 10306 6916 10318 6919
rect 10502 6916 10508 6928
rect 10306 6888 10508 6916
rect 10306 6885 10318 6888
rect 10260 6879 10318 6885
rect 10502 6876 10508 6888
rect 10560 6876 10566 6928
rect 14366 6916 14372 6928
rect 14016 6888 14372 6916
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 9732 6820 10456 6848
rect 9732 6808 9738 6820
rect 10428 6780 10456 6820
rect 11514 6808 11520 6860
rect 11572 6848 11578 6860
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11572 6820 11805 6848
rect 11572 6808 11578 6820
rect 11793 6817 11805 6820
rect 11839 6817 11851 6851
rect 12618 6848 12624 6860
rect 12579 6820 12624 6848
rect 11793 6811 11851 6817
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 14016 6857 14044 6888
rect 14366 6876 14372 6888
rect 14424 6876 14430 6928
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 13412 6820 13461 6848
rect 13412 6808 13418 6820
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 14001 6851 14059 6857
rect 14001 6817 14013 6851
rect 14047 6817 14059 6851
rect 14001 6811 14059 6817
rect 14636 6851 14694 6857
rect 14636 6817 14648 6851
rect 14682 6848 14694 6851
rect 15378 6848 15384 6860
rect 14682 6820 15384 6848
rect 14682 6817 14694 6820
rect 14636 6811 14694 6817
rect 15378 6808 15384 6820
rect 15436 6808 15442 6860
rect 16097 6851 16155 6857
rect 16097 6848 16109 6851
rect 15672 6820 16109 6848
rect 10505 6783 10563 6789
rect 10505 6780 10517 6783
rect 10428 6752 10517 6780
rect 10505 6749 10517 6752
rect 10551 6749 10563 6783
rect 10505 6743 10563 6749
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 10689 6783 10747 6789
rect 10689 6780 10701 6783
rect 10652 6752 10701 6780
rect 10652 6740 10658 6752
rect 10689 6749 10701 6752
rect 10735 6780 10747 6783
rect 10778 6780 10784 6792
rect 10735 6752 10784 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 8938 6604 8944 6656
rect 8996 6644 9002 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 8996 6616 9137 6644
rect 8996 6604 9002 6616
rect 9125 6613 9137 6616
rect 9171 6644 9183 6647
rect 10888 6644 10916 6743
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 11112 6752 11897 6780
rect 11112 6740 11118 6752
rect 11885 6749 11897 6752
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 11146 6672 11152 6724
rect 11204 6712 11210 6724
rect 11333 6715 11391 6721
rect 11333 6712 11345 6715
rect 11204 6684 11345 6712
rect 11204 6672 11210 6684
rect 11333 6681 11345 6684
rect 11379 6681 11391 6715
rect 11992 6712 12020 6743
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 12584 6752 12725 6780
rect 12584 6740 12590 6752
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 12894 6780 12900 6792
rect 12855 6752 12900 6780
rect 12713 6743 12771 6749
rect 12894 6740 12900 6752
rect 12952 6740 12958 6792
rect 13538 6780 13544 6792
rect 13499 6752 13544 6780
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 13633 6783 13691 6789
rect 13633 6749 13645 6783
rect 13679 6749 13691 6783
rect 14366 6780 14372 6792
rect 14327 6752 14372 6780
rect 13633 6743 13691 6749
rect 12912 6712 12940 6740
rect 13648 6712 13676 6743
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 11333 6675 11391 6681
rect 11900 6684 13676 6712
rect 15672 6712 15700 6820
rect 16097 6817 16109 6820
rect 16143 6817 16155 6851
rect 17236 6848 17264 6947
rect 20898 6944 20904 6956
rect 20956 6984 20962 6996
rect 21726 6984 21732 6996
rect 20956 6956 21732 6984
rect 20956 6944 20962 6956
rect 21726 6944 21732 6956
rect 21784 6944 21790 6996
rect 19150 6876 19156 6928
rect 19208 6916 19214 6928
rect 20622 6916 20628 6928
rect 19208 6888 20628 6916
rect 19208 6876 19214 6888
rect 20622 6876 20628 6888
rect 20680 6876 20686 6928
rect 21634 6916 21640 6928
rect 20824 6888 21640 6916
rect 17586 6848 17592 6860
rect 17236 6820 17592 6848
rect 16097 6811 16155 6817
rect 17586 6808 17592 6820
rect 17644 6848 17650 6860
rect 18426 6851 18484 6857
rect 18426 6848 18438 6851
rect 17644 6820 18438 6848
rect 17644 6808 17650 6820
rect 18426 6817 18438 6820
rect 18472 6817 18484 6851
rect 18782 6848 18788 6860
rect 18743 6820 18788 6848
rect 18426 6811 18484 6817
rect 18782 6808 18788 6820
rect 18840 6848 18846 6860
rect 19334 6848 19340 6860
rect 18840 6820 19340 6848
rect 18840 6808 18846 6820
rect 19334 6808 19340 6820
rect 19392 6808 19398 6860
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 20824 6848 20852 6888
rect 21634 6876 21640 6888
rect 21692 6876 21698 6928
rect 19843 6820 20852 6848
rect 20901 6851 20959 6857
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 20901 6817 20913 6851
rect 20947 6848 20959 6851
rect 20947 6820 21496 6848
rect 20947 6817 20959 6820
rect 20901 6811 20959 6817
rect 15746 6740 15752 6792
rect 15804 6780 15810 6792
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15804 6752 15853 6780
rect 15804 6740 15810 6752
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6780 19119 6783
rect 20257 6783 20315 6789
rect 19107 6752 20116 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 15672 6684 15792 6712
rect 9171 6616 10916 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11900 6644 11928 6684
rect 15764 6656 15792 6684
rect 11020 6616 11928 6644
rect 14185 6647 14243 6653
rect 11020 6604 11026 6616
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 15286 6644 15292 6656
rect 14231 6616 15292 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 15746 6644 15752 6656
rect 15707 6616 15752 6644
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 15856 6644 15884 6743
rect 17126 6672 17132 6724
rect 17184 6712 17190 6724
rect 17313 6715 17371 6721
rect 17313 6712 17325 6715
rect 17184 6684 17325 6712
rect 17184 6672 17190 6684
rect 17313 6681 17325 6684
rect 17359 6681 17371 6715
rect 17313 6675 17371 6681
rect 16206 6644 16212 6656
rect 15856 6616 16212 6644
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 18708 6644 18736 6743
rect 19978 6712 19984 6724
rect 19939 6684 19984 6712
rect 19978 6672 19984 6684
rect 20036 6672 20042 6724
rect 17000 6616 18736 6644
rect 20088 6644 20116 6752
rect 20257 6749 20269 6783
rect 20303 6749 20315 6783
rect 20257 6743 20315 6749
rect 20272 6712 20300 6743
rect 20346 6740 20352 6792
rect 20404 6780 20410 6792
rect 20806 6780 20812 6792
rect 20404 6752 20449 6780
rect 20548 6752 20812 6780
rect 20404 6740 20410 6752
rect 20438 6712 20444 6724
rect 20272 6684 20444 6712
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 20548 6644 20576 6752
rect 20806 6740 20812 6752
rect 20864 6740 20870 6792
rect 21174 6780 21180 6792
rect 21100 6752 21180 6780
rect 20622 6672 20628 6724
rect 20680 6712 20686 6724
rect 21100 6721 21128 6752
rect 21174 6740 21180 6752
rect 21232 6740 21238 6792
rect 21085 6715 21143 6721
rect 20680 6684 20935 6712
rect 20680 6672 20686 6684
rect 20806 6644 20812 6656
rect 20088 6616 20576 6644
rect 20767 6616 20812 6644
rect 17000 6604 17006 6616
rect 20806 6604 20812 6616
rect 20864 6604 20870 6656
rect 20907 6644 20935 6684
rect 21085 6681 21097 6715
rect 21131 6681 21143 6715
rect 21468 6712 21496 6820
rect 21542 6808 21548 6860
rect 21600 6848 21606 6860
rect 22750 6851 22808 6857
rect 22750 6848 22762 6851
rect 21600 6820 22762 6848
rect 21600 6808 21606 6820
rect 22750 6817 22762 6820
rect 22796 6817 22808 6851
rect 22750 6811 22808 6817
rect 23017 6783 23075 6789
rect 23017 6749 23029 6783
rect 23063 6749 23075 6783
rect 23017 6743 23075 6749
rect 21468 6684 22094 6712
rect 21085 6675 21143 6681
rect 21177 6647 21235 6653
rect 21177 6644 21189 6647
rect 20907 6616 21189 6644
rect 21177 6613 21189 6616
rect 21223 6613 21235 6647
rect 21634 6644 21640 6656
rect 21595 6616 21640 6644
rect 21177 6607 21235 6613
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 22066 6644 22094 6684
rect 22738 6644 22744 6656
rect 22066 6616 22744 6644
rect 22738 6604 22744 6616
rect 22796 6604 22802 6656
rect 22830 6604 22836 6656
rect 22888 6644 22894 6656
rect 23032 6644 23060 6743
rect 22888 6616 23060 6644
rect 22888 6604 22894 6616
rect 1104 6554 23460 6576
rect 1104 6502 4714 6554
rect 4766 6502 4778 6554
rect 4830 6502 4842 6554
rect 4894 6502 4906 6554
rect 4958 6502 12178 6554
rect 12230 6502 12242 6554
rect 12294 6502 12306 6554
rect 12358 6502 12370 6554
rect 12422 6502 19642 6554
rect 19694 6502 19706 6554
rect 19758 6502 19770 6554
rect 19822 6502 19834 6554
rect 19886 6502 23460 6554
rect 1104 6480 23460 6502
rect 10042 6440 10048 6452
rect 10003 6412 10048 6440
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 11514 6440 11520 6452
rect 11475 6412 11520 6440
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 13081 6443 13139 6449
rect 13081 6440 13093 6443
rect 12676 6412 13093 6440
rect 12676 6400 12682 6412
rect 13081 6409 13093 6412
rect 13127 6409 13139 6443
rect 13081 6403 13139 6409
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 13872 6412 14565 6440
rect 13872 6400 13878 6412
rect 14553 6409 14565 6412
rect 14599 6409 14611 6443
rect 14553 6403 14611 6409
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 10137 6307 10195 6313
rect 10137 6304 10149 6307
rect 9732 6276 10149 6304
rect 9732 6264 9738 6276
rect 10137 6273 10149 6276
rect 10183 6273 10195 6307
rect 14568 6304 14596 6403
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 15436 6412 16037 6440
rect 15436 6400 15442 6412
rect 16025 6409 16037 6412
rect 16071 6409 16083 6443
rect 16025 6403 16083 6409
rect 16577 6443 16635 6449
rect 16577 6409 16589 6443
rect 16623 6440 16635 6443
rect 17310 6440 17316 6452
rect 16623 6412 17316 6440
rect 16623 6409 16635 6412
rect 16577 6403 16635 6409
rect 17310 6400 17316 6412
rect 17368 6400 17374 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 18325 6443 18383 6449
rect 18325 6440 18337 6443
rect 18012 6412 18337 6440
rect 18012 6400 18018 6412
rect 18325 6409 18337 6412
rect 18371 6409 18383 6443
rect 18325 6403 18383 6409
rect 18509 6443 18567 6449
rect 18509 6409 18521 6443
rect 18555 6440 18567 6443
rect 19150 6440 19156 6452
rect 18555 6412 19156 6440
rect 18555 6409 18567 6412
rect 18509 6403 18567 6409
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 19337 6443 19395 6449
rect 19337 6409 19349 6443
rect 19383 6440 19395 6443
rect 19383 6412 20392 6440
rect 19383 6409 19395 6412
rect 19337 6403 19395 6409
rect 18874 6332 18880 6384
rect 18932 6372 18938 6384
rect 20364 6372 20392 6412
rect 20438 6400 20444 6452
rect 20496 6440 20502 6452
rect 22646 6440 22652 6452
rect 20496 6412 22652 6440
rect 20496 6400 20502 6412
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 20714 6372 20720 6384
rect 18932 6344 19472 6372
rect 20364 6344 20720 6372
rect 18932 6332 18938 6344
rect 18785 6307 18843 6313
rect 14568 6276 14780 6304
rect 10137 6267 10195 6273
rect 8938 6245 8944 6248
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6205 8723 6239
rect 8932 6236 8944 6245
rect 8899 6208 8944 6236
rect 8665 6199 8723 6205
rect 8932 6199 8944 6208
rect 8680 6168 8708 6199
rect 8938 6196 8944 6199
rect 8996 6196 9002 6248
rect 9692 6168 9720 6264
rect 10152 6236 10180 6267
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 10152 6208 11713 6236
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 13078 6196 13084 6248
rect 13136 6236 13142 6248
rect 13173 6239 13231 6245
rect 13173 6236 13185 6239
rect 13136 6208 13185 6236
rect 13136 6196 13142 6208
rect 13173 6205 13185 6208
rect 13219 6236 13231 6239
rect 14366 6236 14372 6248
rect 13219 6208 14372 6236
rect 13219 6205 13231 6208
rect 13173 6199 13231 6205
rect 14366 6196 14372 6208
rect 14424 6236 14430 6248
rect 14645 6239 14703 6245
rect 14645 6236 14657 6239
rect 14424 6208 14657 6236
rect 14424 6196 14430 6208
rect 14645 6205 14657 6208
rect 14691 6205 14703 6239
rect 14752 6236 14780 6276
rect 18785 6273 18797 6307
rect 18831 6304 18843 6307
rect 19150 6304 19156 6316
rect 18831 6276 19156 6304
rect 18831 6273 18843 6276
rect 18785 6267 18843 6273
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 19444 6304 19472 6344
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 20806 6332 20812 6384
rect 20864 6372 20870 6384
rect 23106 6372 23112 6384
rect 20864 6344 23112 6372
rect 20864 6332 20870 6344
rect 23106 6332 23112 6344
rect 23164 6332 23170 6384
rect 21453 6307 21511 6313
rect 21453 6304 21465 6307
rect 19444 6276 19564 6304
rect 14901 6239 14959 6245
rect 14901 6236 14913 6239
rect 14752 6208 14913 6236
rect 14645 6199 14703 6205
rect 14901 6205 14913 6208
rect 14947 6205 14959 6239
rect 14901 6199 14959 6205
rect 8680 6140 9720 6168
rect 10404 6171 10462 6177
rect 10404 6137 10416 6171
rect 10450 6168 10462 6171
rect 11054 6168 11060 6180
rect 10450 6140 11060 6168
rect 10450 6137 10462 6140
rect 10404 6131 10462 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 11968 6171 12026 6177
rect 11968 6137 11980 6171
rect 12014 6168 12026 6171
rect 12526 6168 12532 6180
rect 12014 6140 12532 6168
rect 12014 6137 12026 6140
rect 11968 6131 12026 6137
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 13354 6128 13360 6180
rect 13412 6177 13418 6180
rect 13412 6171 13476 6177
rect 13412 6137 13430 6171
rect 13464 6137 13476 6171
rect 14660 6168 14688 6199
rect 15470 6196 15476 6248
rect 15528 6236 15534 6248
rect 16117 6239 16175 6245
rect 16117 6236 16129 6239
rect 15528 6208 16129 6236
rect 15528 6196 15534 6208
rect 16117 6205 16129 6208
rect 16163 6205 16175 6239
rect 16942 6236 16948 6248
rect 16903 6208 16948 6236
rect 16117 6199 16175 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 19426 6236 19432 6248
rect 19387 6208 19432 6236
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 19536 6236 19564 6276
rect 20456 6276 21465 6304
rect 20456 6236 20484 6276
rect 21453 6273 21465 6276
rect 21499 6273 21511 6307
rect 21453 6267 21511 6273
rect 19536 6208 20484 6236
rect 21269 6239 21327 6245
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 22278 6236 22284 6248
rect 21315 6208 22094 6236
rect 22239 6208 22284 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 14734 6168 14740 6180
rect 14660 6140 14740 6168
rect 13412 6131 13476 6137
rect 13412 6128 13418 6131
rect 14734 6128 14740 6140
rect 14792 6128 14798 6180
rect 17126 6128 17132 6180
rect 17184 6177 17190 6180
rect 17184 6171 17248 6177
rect 17184 6137 17202 6171
rect 17236 6137 17248 6171
rect 17184 6131 17248 6137
rect 17184 6128 17190 6131
rect 18230 6128 18236 6180
rect 18288 6168 18294 6180
rect 18782 6168 18788 6180
rect 18288 6140 18788 6168
rect 18288 6128 18294 6140
rect 18782 6128 18788 6140
rect 18840 6128 18846 6180
rect 18877 6171 18935 6177
rect 18877 6137 18889 6171
rect 18923 6168 18935 6171
rect 19696 6171 19754 6177
rect 18923 6140 19656 6168
rect 18923 6137 18935 6140
rect 18877 6131 18935 6137
rect 18966 6100 18972 6112
rect 18927 6072 18972 6100
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 19628 6100 19656 6140
rect 19696 6137 19708 6171
rect 19742 6168 19754 6171
rect 20714 6168 20720 6180
rect 19742 6140 20720 6168
rect 19742 6137 19754 6140
rect 19696 6131 19754 6137
rect 20714 6128 20720 6140
rect 20772 6128 20778 6180
rect 21726 6168 21732 6180
rect 21687 6140 21732 6168
rect 21726 6128 21732 6140
rect 21784 6128 21790 6180
rect 21910 6168 21916 6180
rect 21871 6140 21916 6168
rect 21910 6128 21916 6140
rect 21968 6128 21974 6180
rect 20622 6100 20628 6112
rect 19628 6072 20628 6100
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 20806 6100 20812 6112
rect 20767 6072 20812 6100
rect 20806 6060 20812 6072
rect 20864 6060 20870 6112
rect 20898 6060 20904 6112
rect 20956 6100 20962 6112
rect 20956 6072 21001 6100
rect 20956 6060 20962 6072
rect 21266 6060 21272 6112
rect 21324 6100 21330 6112
rect 21361 6103 21419 6109
rect 21361 6100 21373 6103
rect 21324 6072 21373 6100
rect 21324 6060 21330 6072
rect 21361 6069 21373 6072
rect 21407 6069 21419 6103
rect 22066 6100 22094 6208
rect 22278 6196 22284 6208
rect 22336 6196 22342 6248
rect 22738 6168 22744 6180
rect 22699 6140 22744 6168
rect 22738 6128 22744 6140
rect 22796 6128 22802 6180
rect 23014 6100 23020 6112
rect 22066 6072 23020 6100
rect 21361 6063 21419 6069
rect 23014 6060 23020 6072
rect 23072 6060 23078 6112
rect 1104 6010 23460 6032
rect 1104 5958 8446 6010
rect 8498 5958 8510 6010
rect 8562 5958 8574 6010
rect 8626 5958 8638 6010
rect 8690 5958 15910 6010
rect 15962 5958 15974 6010
rect 16026 5958 16038 6010
rect 16090 5958 16102 6010
rect 16154 5958 23460 6010
rect 1104 5936 23460 5958
rect 11054 5896 11060 5908
rect 11015 5868 11060 5896
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 12526 5896 12532 5908
rect 12487 5868 12532 5896
rect 12526 5856 12532 5868
rect 12584 5856 12590 5908
rect 13538 5856 13544 5908
rect 13596 5896 13602 5908
rect 14001 5899 14059 5905
rect 14001 5896 14013 5899
rect 13596 5868 14013 5896
rect 13596 5856 13602 5868
rect 14001 5865 14013 5868
rect 14047 5865 14059 5899
rect 14001 5859 14059 5865
rect 14553 5899 14611 5905
rect 14553 5865 14565 5899
rect 14599 5896 14611 5899
rect 15194 5896 15200 5908
rect 14599 5868 15200 5896
rect 14599 5865 14611 5868
rect 14553 5859 14611 5865
rect 15194 5856 15200 5868
rect 15252 5856 15258 5908
rect 15289 5899 15347 5905
rect 15289 5865 15301 5899
rect 15335 5896 15347 5899
rect 15654 5896 15660 5908
rect 15335 5868 15660 5896
rect 15335 5865 15347 5868
rect 15289 5859 15347 5865
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 17218 5856 17224 5908
rect 17276 5896 17282 5908
rect 17313 5899 17371 5905
rect 17313 5896 17325 5899
rect 17276 5868 17325 5896
rect 17276 5856 17282 5868
rect 17313 5865 17325 5868
rect 17359 5896 17371 5899
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17359 5868 17693 5896
rect 17359 5865 17371 5868
rect 17313 5859 17371 5865
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 18325 5899 18383 5905
rect 18325 5865 18337 5899
rect 18371 5896 18383 5899
rect 18506 5896 18512 5908
rect 18371 5868 18512 5896
rect 18371 5865 18383 5868
rect 18325 5859 18383 5865
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 18601 5899 18659 5905
rect 18601 5865 18613 5899
rect 18647 5896 18659 5899
rect 18966 5896 18972 5908
rect 18647 5868 18972 5896
rect 18647 5865 18659 5868
rect 18601 5859 18659 5865
rect 18966 5856 18972 5868
rect 19024 5856 19030 5908
rect 19429 5899 19487 5905
rect 19429 5865 19441 5899
rect 19475 5896 19487 5899
rect 20346 5896 20352 5908
rect 19475 5868 20352 5896
rect 19475 5865 19487 5868
rect 19429 5859 19487 5865
rect 9944 5831 10002 5837
rect 9944 5797 9956 5831
rect 9990 5828 10002 5831
rect 10042 5828 10048 5840
rect 9990 5800 10048 5828
rect 9990 5797 10002 5800
rect 9944 5791 10002 5797
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 11416 5831 11474 5837
rect 11416 5797 11428 5831
rect 11462 5828 11474 5831
rect 11514 5828 11520 5840
rect 11462 5800 11520 5828
rect 11462 5797 11474 5800
rect 11416 5791 11474 5797
rect 11514 5788 11520 5800
rect 11572 5788 11578 5840
rect 12618 5788 12624 5840
rect 12676 5828 12682 5840
rect 12866 5831 12924 5837
rect 12866 5828 12878 5831
rect 12676 5800 12878 5828
rect 12676 5788 12682 5800
rect 12866 5797 12878 5800
rect 12912 5797 12924 5831
rect 12866 5791 12924 5797
rect 13078 5788 13084 5840
rect 13136 5788 13142 5840
rect 15562 5788 15568 5840
rect 15620 5828 15626 5840
rect 16178 5831 16236 5837
rect 16178 5828 16190 5831
rect 15620 5800 16190 5828
rect 15620 5788 15626 5800
rect 16178 5797 16190 5800
rect 16224 5797 16236 5831
rect 18046 5828 18052 5840
rect 16178 5791 16236 5797
rect 17604 5800 18052 5828
rect 9674 5760 9680 5772
rect 9635 5732 9680 5760
rect 9674 5720 9680 5732
rect 9732 5760 9738 5772
rect 11149 5763 11207 5769
rect 11149 5760 11161 5763
rect 9732 5732 11161 5760
rect 9732 5720 9738 5732
rect 11149 5729 11161 5732
rect 11195 5729 11207 5763
rect 13096 5760 13124 5788
rect 11149 5723 11207 5729
rect 12636 5732 13124 5760
rect 14369 5763 14427 5769
rect 12636 5701 12664 5732
rect 14369 5729 14381 5763
rect 14415 5760 14427 5763
rect 14550 5760 14556 5772
rect 14415 5732 14556 5760
rect 14415 5729 14427 5732
rect 14369 5723 14427 5729
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 14642 5720 14648 5772
rect 14700 5760 14706 5772
rect 15378 5760 15384 5772
rect 14700 5732 14745 5760
rect 15339 5732 15384 5760
rect 14700 5720 14706 5732
rect 15378 5720 15384 5732
rect 15436 5720 15442 5772
rect 15933 5763 15991 5769
rect 15933 5729 15945 5763
rect 15979 5760 15991 5763
rect 16022 5760 16028 5772
rect 15979 5732 16028 5760
rect 15979 5729 15991 5732
rect 15933 5723 15991 5729
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5692 15255 5695
rect 15746 5692 15752 5704
rect 15243 5664 15752 5692
rect 15243 5661 15255 5664
rect 15197 5655 15255 5661
rect 15746 5652 15752 5664
rect 15804 5652 15810 5704
rect 14734 5584 14740 5636
rect 14792 5624 14798 5636
rect 14829 5627 14887 5633
rect 14829 5624 14841 5627
rect 14792 5596 14841 5624
rect 14792 5584 14798 5596
rect 14829 5593 14841 5596
rect 14875 5624 14887 5627
rect 15948 5624 15976 5723
rect 16022 5720 16028 5732
rect 16080 5720 16086 5772
rect 17604 5701 17632 5800
rect 18046 5788 18052 5800
rect 18104 5788 18110 5840
rect 19444 5828 19472 5859
rect 20346 5856 20352 5868
rect 20404 5856 20410 5908
rect 21542 5896 21548 5908
rect 21284 5868 21548 5896
rect 21082 5828 21088 5840
rect 18432 5800 19472 5828
rect 21043 5800 21088 5828
rect 17773 5763 17831 5769
rect 17773 5729 17785 5763
rect 17819 5760 17831 5763
rect 17862 5760 17868 5772
rect 17819 5732 17868 5760
rect 17819 5729 17831 5732
rect 17773 5723 17831 5729
rect 17862 5720 17868 5732
rect 17920 5720 17926 5772
rect 18432 5769 18460 5800
rect 21082 5788 21088 5800
rect 21140 5788 21146 5840
rect 21284 5837 21312 5868
rect 21542 5856 21548 5868
rect 21600 5856 21606 5908
rect 21269 5831 21327 5837
rect 21269 5797 21281 5831
rect 21315 5797 21327 5831
rect 21269 5791 21327 5797
rect 22462 5788 22468 5840
rect 22520 5828 22526 5840
rect 22658 5831 22716 5837
rect 22658 5828 22670 5831
rect 22520 5800 22670 5828
rect 22520 5788 22526 5800
rect 22658 5797 22670 5800
rect 22704 5797 22716 5831
rect 22658 5791 22716 5797
rect 18417 5763 18475 5769
rect 18417 5729 18429 5763
rect 18463 5729 18475 5763
rect 19061 5763 19119 5769
rect 19061 5760 19073 5763
rect 18417 5723 18475 5729
rect 18524 5732 19073 5760
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5661 17647 5695
rect 17589 5655 17647 5661
rect 17678 5652 17684 5704
rect 17736 5692 17742 5704
rect 18524 5692 18552 5732
rect 19061 5729 19073 5732
rect 19107 5729 19119 5763
rect 19061 5723 19119 5729
rect 19150 5720 19156 5772
rect 19208 5760 19214 5772
rect 19880 5763 19938 5769
rect 19880 5760 19892 5763
rect 19208 5732 19892 5760
rect 19208 5720 19214 5732
rect 19880 5729 19892 5732
rect 19926 5760 19938 5763
rect 21634 5760 21640 5772
rect 19926 5732 21640 5760
rect 19926 5729 19938 5732
rect 19880 5723 19938 5729
rect 21634 5720 21640 5732
rect 21692 5720 21698 5772
rect 22830 5720 22836 5772
rect 22888 5760 22894 5772
rect 22925 5763 22983 5769
rect 22925 5760 22937 5763
rect 22888 5732 22937 5760
rect 22888 5720 22894 5732
rect 22925 5729 22937 5732
rect 22971 5729 22983 5763
rect 22925 5723 22983 5729
rect 18874 5692 18880 5704
rect 17736 5664 18552 5692
rect 18835 5664 18880 5692
rect 17736 5652 17742 5664
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 18969 5695 19027 5701
rect 18969 5661 18981 5695
rect 19015 5661 19027 5695
rect 18969 5655 19027 5661
rect 14875 5596 15976 5624
rect 14875 5593 14887 5596
rect 14829 5587 14887 5593
rect 17954 5584 17960 5636
rect 18012 5624 18018 5636
rect 18984 5624 19012 5655
rect 19518 5652 19524 5704
rect 19576 5692 19582 5704
rect 19613 5695 19671 5701
rect 19613 5692 19625 5695
rect 19576 5664 19625 5692
rect 19576 5652 19582 5664
rect 19613 5661 19625 5664
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 18012 5596 19012 5624
rect 18012 5584 18018 5596
rect 20714 5584 20720 5636
rect 20772 5624 20778 5636
rect 20993 5627 21051 5633
rect 20993 5624 21005 5627
rect 20772 5596 21005 5624
rect 20772 5584 20778 5596
rect 20993 5593 21005 5596
rect 21039 5624 21051 5627
rect 21039 5596 21588 5624
rect 21039 5593 21051 5596
rect 20993 5587 21051 5593
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 15749 5559 15807 5565
rect 15749 5556 15761 5559
rect 15528 5528 15761 5556
rect 15528 5516 15534 5528
rect 15749 5525 15761 5528
rect 15795 5525 15807 5559
rect 18138 5556 18144 5568
rect 18099 5528 18144 5556
rect 15749 5519 15807 5525
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 18506 5516 18512 5568
rect 18564 5556 18570 5568
rect 20346 5556 20352 5568
rect 18564 5528 20352 5556
rect 18564 5516 18570 5528
rect 20346 5516 20352 5528
rect 20404 5516 20410 5568
rect 21450 5556 21456 5568
rect 21411 5528 21456 5556
rect 21450 5516 21456 5528
rect 21508 5516 21514 5568
rect 21560 5556 21588 5596
rect 22186 5556 22192 5568
rect 21560 5528 22192 5556
rect 22186 5516 22192 5528
rect 22244 5516 22250 5568
rect 1104 5466 23460 5488
rect 1104 5414 4714 5466
rect 4766 5414 4778 5466
rect 4830 5414 4842 5466
rect 4894 5414 4906 5466
rect 4958 5414 12178 5466
rect 12230 5414 12242 5466
rect 12294 5414 12306 5466
rect 12358 5414 12370 5466
rect 12422 5414 19642 5466
rect 19694 5414 19706 5466
rect 19758 5414 19770 5466
rect 19822 5414 19834 5466
rect 19886 5414 23460 5466
rect 1104 5392 23460 5414
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 13354 5352 13360 5364
rect 12299 5324 13360 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 17862 5312 17868 5364
rect 17920 5352 17926 5364
rect 18325 5355 18383 5361
rect 18325 5352 18337 5355
rect 17920 5324 18337 5352
rect 17920 5312 17926 5324
rect 18325 5321 18337 5324
rect 18371 5321 18383 5355
rect 18325 5315 18383 5321
rect 16025 5287 16083 5293
rect 16025 5253 16037 5287
rect 16071 5284 16083 5287
rect 22370 5284 22376 5296
rect 16071 5256 16988 5284
rect 16071 5253 16083 5256
rect 16025 5247 16083 5253
rect 16960 5228 16988 5256
rect 19444 5256 22376 5284
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 14734 5216 14740 5228
rect 13679 5188 14740 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 15378 5176 15384 5228
rect 15436 5216 15442 5228
rect 16117 5219 16175 5225
rect 16117 5216 16129 5219
rect 15436 5188 16129 5216
rect 15436 5176 15442 5188
rect 16117 5185 16129 5188
rect 16163 5185 16175 5219
rect 16942 5216 16948 5228
rect 16903 5188 16948 5216
rect 16117 5179 16175 5185
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 19444 5225 19472 5256
rect 22370 5244 22376 5256
rect 22428 5244 22434 5296
rect 18877 5219 18935 5225
rect 18877 5216 18889 5219
rect 18196 5188 18889 5216
rect 18196 5176 18202 5188
rect 18877 5185 18889 5188
rect 18923 5185 18935 5219
rect 18877 5179 18935 5185
rect 18969 5219 19027 5225
rect 18969 5185 18981 5219
rect 19015 5185 19027 5219
rect 18969 5179 19027 5185
rect 19429 5219 19487 5225
rect 19429 5185 19441 5219
rect 19475 5185 19487 5219
rect 19429 5179 19487 5185
rect 19613 5219 19671 5225
rect 19613 5185 19625 5219
rect 19659 5216 19671 5219
rect 19659 5188 20944 5216
rect 19659 5185 19671 5188
rect 19613 5179 19671 5185
rect 13377 5151 13435 5157
rect 13377 5117 13389 5151
rect 13423 5148 13435 5151
rect 13538 5148 13544 5160
rect 13423 5120 13544 5148
rect 13423 5117 13435 5120
rect 13377 5111 13435 5117
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 16298 5148 16304 5160
rect 15887 5120 16304 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 16298 5108 16304 5120
rect 16356 5108 16362 5160
rect 17218 5157 17224 5160
rect 16577 5151 16635 5157
rect 16577 5117 16589 5151
rect 16623 5117 16635 5151
rect 17212 5148 17224 5157
rect 17179 5120 17224 5148
rect 16577 5111 16635 5117
rect 17212 5111 17224 5120
rect 16592 5080 16620 5111
rect 17218 5108 17224 5111
rect 17276 5108 17282 5160
rect 18782 5108 18788 5160
rect 18840 5148 18846 5160
rect 18984 5148 19012 5179
rect 19628 5148 19656 5179
rect 18840 5120 19656 5148
rect 19797 5151 19855 5157
rect 18840 5108 18846 5120
rect 19797 5117 19809 5151
rect 19843 5148 19855 5151
rect 20806 5148 20812 5160
rect 19843 5120 20812 5148
rect 19843 5117 19855 5120
rect 19797 5111 19855 5117
rect 20806 5108 20812 5120
rect 20864 5108 20870 5160
rect 20916 5148 20944 5188
rect 20990 5176 20996 5228
rect 21048 5216 21054 5228
rect 21269 5219 21327 5225
rect 21048 5188 21093 5216
rect 21048 5176 21054 5188
rect 21269 5185 21281 5219
rect 21315 5185 21327 5219
rect 21269 5179 21327 5185
rect 21284 5148 21312 5179
rect 21542 5176 21548 5228
rect 21600 5216 21606 5228
rect 22649 5219 22707 5225
rect 22649 5216 22661 5219
rect 21600 5188 22661 5216
rect 21600 5176 21606 5188
rect 22649 5185 22661 5188
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 22738 5176 22744 5228
rect 22796 5216 22802 5228
rect 22796 5188 22889 5216
rect 22796 5176 22802 5188
rect 20916 5120 21312 5148
rect 19889 5083 19947 5089
rect 16592 5052 18460 5080
rect 16761 5015 16819 5021
rect 16761 4981 16773 5015
rect 16807 5012 16819 5015
rect 17954 5012 17960 5024
rect 16807 4984 17960 5012
rect 16807 4981 16819 4984
rect 16761 4975 16819 4981
rect 17954 4972 17960 4984
rect 18012 4972 18018 5024
rect 18432 5021 18460 5052
rect 19889 5049 19901 5083
rect 19935 5080 19947 5083
rect 19935 5052 20392 5080
rect 19935 5049 19947 5052
rect 19889 5043 19947 5049
rect 18417 5015 18475 5021
rect 18417 4981 18429 5015
rect 18463 4981 18475 5015
rect 18417 4975 18475 4981
rect 18598 4972 18604 5024
rect 18656 5012 18662 5024
rect 18785 5015 18843 5021
rect 18785 5012 18797 5015
rect 18656 4984 18797 5012
rect 18656 4972 18662 4984
rect 18785 4981 18797 4984
rect 18831 4981 18843 5015
rect 18785 4975 18843 4981
rect 19978 4972 19984 5024
rect 20036 5012 20042 5024
rect 20364 5021 20392 5052
rect 20257 5015 20315 5021
rect 20257 5012 20269 5015
rect 20036 4984 20269 5012
rect 20036 4972 20042 4984
rect 20257 4981 20269 4984
rect 20303 4981 20315 5015
rect 20257 4975 20315 4981
rect 20349 5015 20407 5021
rect 20349 4981 20361 5015
rect 20395 4981 20407 5015
rect 20714 5012 20720 5024
rect 20675 4984 20720 5012
rect 20349 4975 20407 4981
rect 20714 4972 20720 4984
rect 20772 4972 20778 5024
rect 20809 5015 20867 5021
rect 20809 4981 20821 5015
rect 20855 5012 20867 5015
rect 21082 5012 21088 5024
rect 20855 4984 21088 5012
rect 20855 4981 20867 4984
rect 20809 4975 20867 4981
rect 21082 4972 21088 4984
rect 21140 4972 21146 5024
rect 21284 5012 21312 5120
rect 21453 5151 21511 5157
rect 21453 5117 21465 5151
rect 21499 5148 21511 5151
rect 22186 5148 22192 5160
rect 21499 5120 22192 5148
rect 21499 5117 21511 5120
rect 21453 5111 21511 5117
rect 22186 5108 22192 5120
rect 22244 5108 22250 5160
rect 22278 5108 22284 5160
rect 22336 5148 22342 5160
rect 22756 5148 22784 5176
rect 22336 5120 22784 5148
rect 22336 5108 22342 5120
rect 21545 5083 21603 5089
rect 21545 5049 21557 5083
rect 21591 5080 21603 5083
rect 21591 5052 22232 5080
rect 21591 5049 21603 5052
rect 21545 5043 21603 5049
rect 21726 5012 21732 5024
rect 21284 4984 21732 5012
rect 21726 4972 21732 4984
rect 21784 4972 21790 5024
rect 21913 5015 21971 5021
rect 21913 4981 21925 5015
rect 21959 5012 21971 5015
rect 22094 5012 22100 5024
rect 21959 4984 22100 5012
rect 21959 4981 21971 4984
rect 21913 4975 21971 4981
rect 22094 4972 22100 4984
rect 22152 4972 22158 5024
rect 22204 5021 22232 5052
rect 22370 5040 22376 5092
rect 22428 5080 22434 5092
rect 23017 5083 23075 5089
rect 23017 5080 23029 5083
rect 22428 5052 23029 5080
rect 22428 5040 22434 5052
rect 23017 5049 23029 5052
rect 23063 5080 23075 5083
rect 23382 5080 23388 5092
rect 23063 5052 23388 5080
rect 23063 5049 23075 5052
rect 23017 5043 23075 5049
rect 23382 5040 23388 5052
rect 23440 5040 23446 5092
rect 22189 5015 22247 5021
rect 22189 4981 22201 5015
rect 22235 4981 22247 5015
rect 22189 4975 22247 4981
rect 22462 4972 22468 5024
rect 22520 5012 22526 5024
rect 22557 5015 22615 5021
rect 22557 5012 22569 5015
rect 22520 4984 22569 5012
rect 22520 4972 22526 4984
rect 22557 4981 22569 4984
rect 22603 4981 22615 5015
rect 22557 4975 22615 4981
rect 1104 4922 23460 4944
rect 1104 4870 8446 4922
rect 8498 4870 8510 4922
rect 8562 4870 8574 4922
rect 8626 4870 8638 4922
rect 8690 4870 15910 4922
rect 15962 4870 15974 4922
rect 16026 4870 16038 4922
rect 16090 4870 16102 4922
rect 16154 4870 23460 4922
rect 1104 4848 23460 4870
rect 16301 4811 16359 4817
rect 16301 4777 16313 4811
rect 16347 4808 16359 4811
rect 17678 4808 17684 4820
rect 16347 4780 17684 4808
rect 16347 4777 16359 4780
rect 16301 4771 16359 4777
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 18598 4808 18604 4820
rect 18559 4780 18604 4808
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 17528 4743 17586 4749
rect 17528 4709 17540 4743
rect 17574 4740 17586 4743
rect 17862 4740 17868 4752
rect 17574 4712 17868 4740
rect 17574 4709 17586 4712
rect 17528 4703 17586 4709
rect 17862 4700 17868 4712
rect 17920 4700 17926 4752
rect 19880 4743 19938 4749
rect 19880 4709 19892 4743
rect 19926 4740 19938 4743
rect 20070 4740 20076 4752
rect 19926 4712 20076 4740
rect 19926 4709 19938 4712
rect 19880 4703 19938 4709
rect 20070 4700 20076 4712
rect 20128 4700 20134 4752
rect 21358 4740 21364 4752
rect 21319 4712 21364 4740
rect 21358 4700 21364 4712
rect 21416 4700 21422 4752
rect 22370 4700 22376 4752
rect 22428 4700 22434 4752
rect 16114 4672 16120 4684
rect 16075 4644 16120 4672
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 17218 4672 17224 4684
rect 16408 4644 17224 4672
rect 16408 4545 16436 4644
rect 17218 4632 17224 4644
rect 17276 4672 17282 4684
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 17276 4644 18153 4672
rect 17276 4632 17282 4644
rect 18141 4641 18153 4644
rect 18187 4641 18199 4675
rect 18141 4635 18199 4641
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4672 18291 4675
rect 18322 4672 18328 4684
rect 18279 4644 18328 4672
rect 18279 4641 18291 4644
rect 18233 4635 18291 4641
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 18690 4632 18696 4684
rect 18748 4672 18754 4684
rect 19061 4675 19119 4681
rect 19061 4672 19073 4675
rect 18748 4644 19073 4672
rect 18748 4632 18754 4644
rect 19061 4641 19073 4644
rect 19107 4641 19119 4675
rect 19061 4635 19119 4641
rect 21177 4675 21235 4681
rect 21177 4641 21189 4675
rect 21223 4672 21235 4675
rect 22388 4672 22416 4700
rect 22554 4672 22560 4684
rect 22612 4681 22618 4684
rect 21223 4644 22416 4672
rect 22524 4644 22560 4672
rect 21223 4641 21235 4644
rect 21177 4635 21235 4641
rect 22554 4632 22560 4644
rect 22612 4635 22624 4681
rect 22830 4672 22836 4684
rect 22791 4644 22836 4672
rect 22612 4632 22618 4635
rect 22830 4632 22836 4644
rect 22888 4632 22894 4684
rect 23106 4672 23112 4684
rect 23067 4644 23112 4672
rect 23106 4632 23112 4644
rect 23164 4632 23170 4684
rect 17770 4604 17776 4616
rect 17731 4576 17776 4604
rect 17770 4564 17776 4576
rect 17828 4564 17834 4616
rect 18046 4604 18052 4616
rect 18007 4576 18052 4604
rect 18046 4564 18052 4576
rect 18104 4564 18110 4616
rect 19150 4604 19156 4616
rect 19111 4576 19156 4604
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4573 19303 4607
rect 19245 4567 19303 4573
rect 16393 4539 16451 4545
rect 16393 4505 16405 4539
rect 16439 4505 16451 4539
rect 18064 4536 18092 4564
rect 19058 4536 19064 4548
rect 18064 4508 19064 4536
rect 16393 4499 16451 4505
rect 19058 4496 19064 4508
rect 19116 4536 19122 4548
rect 19260 4536 19288 4567
rect 19518 4564 19524 4616
rect 19576 4604 19582 4616
rect 19613 4607 19671 4613
rect 19613 4604 19625 4607
rect 19576 4576 19625 4604
rect 19576 4564 19582 4576
rect 19613 4573 19625 4576
rect 19659 4573 19671 4607
rect 19613 4567 19671 4573
rect 20990 4564 20996 4616
rect 21048 4604 21054 4616
rect 21358 4604 21364 4616
rect 21048 4576 21364 4604
rect 21048 4564 21054 4576
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 19116 4508 19288 4536
rect 19116 4496 19122 4508
rect 20622 4496 20628 4548
rect 20680 4536 20686 4548
rect 21453 4539 21511 4545
rect 20680 4508 21128 4536
rect 20680 4496 20686 4508
rect 16666 4428 16672 4480
rect 16724 4468 16730 4480
rect 18693 4471 18751 4477
rect 18693 4468 18705 4471
rect 16724 4440 18705 4468
rect 16724 4428 16730 4440
rect 18693 4437 18705 4440
rect 18739 4437 18751 4471
rect 20990 4468 20996 4480
rect 20951 4440 20996 4468
rect 18693 4431 18751 4437
rect 20990 4428 20996 4440
rect 21048 4428 21054 4480
rect 21100 4468 21128 4508
rect 21453 4505 21465 4539
rect 21499 4536 21511 4539
rect 21542 4536 21548 4548
rect 21499 4508 21548 4536
rect 21499 4505 21511 4508
rect 21453 4499 21511 4505
rect 21542 4496 21548 4508
rect 21600 4496 21606 4548
rect 22925 4471 22983 4477
rect 22925 4468 22937 4471
rect 21100 4440 22937 4468
rect 22925 4437 22937 4440
rect 22971 4437 22983 4471
rect 22925 4431 22983 4437
rect 1104 4378 23460 4400
rect 1104 4326 4714 4378
rect 4766 4326 4778 4378
rect 4830 4326 4842 4378
rect 4894 4326 4906 4378
rect 4958 4326 12178 4378
rect 12230 4326 12242 4378
rect 12294 4326 12306 4378
rect 12358 4326 12370 4378
rect 12422 4326 19642 4378
rect 19694 4326 19706 4378
rect 19758 4326 19770 4378
rect 19822 4326 19834 4378
rect 19886 4326 23460 4378
rect 1104 4304 23460 4326
rect 16025 4267 16083 4273
rect 16025 4233 16037 4267
rect 16071 4264 16083 4267
rect 16114 4264 16120 4276
rect 16071 4236 16120 4264
rect 16071 4233 16083 4236
rect 16025 4227 16083 4233
rect 16114 4224 16120 4236
rect 16172 4224 16178 4276
rect 18782 4264 18788 4276
rect 16592 4236 18788 4264
rect 16592 4137 16620 4236
rect 18782 4224 18788 4236
rect 18840 4224 18846 4276
rect 21358 4224 21364 4276
rect 21416 4264 21422 4276
rect 22186 4264 22192 4276
rect 21416 4236 21680 4264
rect 22147 4236 22192 4264
rect 21416 4224 21422 4236
rect 18322 4196 18328 4208
rect 18283 4168 18328 4196
rect 18322 4156 18328 4168
rect 18380 4156 18386 4208
rect 20438 4196 20444 4208
rect 19996 4168 20444 4196
rect 16577 4131 16635 4137
rect 16577 4097 16589 4131
rect 16623 4097 16635 4131
rect 16942 4128 16948 4140
rect 16903 4100 16948 4128
rect 16577 4091 16635 4097
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 19426 4088 19432 4140
rect 19484 4128 19490 4140
rect 19996 4128 20024 4168
rect 20438 4156 20444 4168
rect 20496 4156 20502 4208
rect 20162 4128 20168 4140
rect 19484 4100 20024 4128
rect 20123 4100 20168 4128
rect 19484 4088 19490 4100
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20530 4128 20536 4140
rect 20491 4100 20536 4128
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 21652 4128 21680 4236
rect 22186 4224 22192 4236
rect 22244 4224 22250 4276
rect 22005 4199 22063 4205
rect 22005 4165 22017 4199
rect 22051 4196 22063 4199
rect 22462 4196 22468 4208
rect 22051 4168 22468 4196
rect 22051 4165 22063 4168
rect 22005 4159 22063 4165
rect 22462 4156 22468 4168
rect 22520 4156 22526 4208
rect 22278 4128 22284 4140
rect 21652 4100 22284 4128
rect 22278 4088 22284 4100
rect 22336 4128 22342 4140
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 22336 4100 22753 4128
rect 22336 4088 22342 4100
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 16393 4063 16451 4069
rect 16393 4029 16405 4063
rect 16439 4060 16451 4063
rect 16666 4060 16672 4072
rect 16439 4032 16672 4060
rect 16439 4029 16451 4032
rect 16393 4023 16451 4029
rect 16666 4020 16672 4032
rect 16724 4020 16730 4072
rect 15933 3995 15991 4001
rect 15933 3961 15945 3995
rect 15979 3992 15991 3995
rect 16960 3992 16988 4088
rect 17218 4069 17224 4072
rect 17212 4060 17224 4069
rect 17179 4032 17224 4060
rect 17212 4023 17224 4032
rect 17218 4020 17224 4023
rect 17276 4020 17282 4072
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4060 18475 4063
rect 19518 4060 19524 4072
rect 18463 4032 19524 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 17770 3992 17776 4004
rect 15979 3964 16896 3992
rect 16960 3964 17776 3992
rect 15979 3961 15991 3964
rect 15933 3955 15991 3961
rect 16482 3924 16488 3936
rect 16443 3896 16488 3924
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 16868 3924 16896 3964
rect 17770 3952 17776 3964
rect 17828 3992 17834 4004
rect 18432 3992 18460 4023
rect 19518 4020 19524 4032
rect 19576 4020 19582 4072
rect 20346 4060 20352 4072
rect 20307 4032 20352 4060
rect 20346 4020 20352 4032
rect 20404 4020 20410 4072
rect 20622 4060 20628 4072
rect 20583 4032 20628 4060
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 21634 4060 21640 4072
rect 20824 4032 21640 4060
rect 18690 4001 18696 4004
rect 18684 3992 18696 4001
rect 17828 3964 18460 3992
rect 18651 3964 18696 3992
rect 17828 3952 17834 3964
rect 18684 3955 18696 3964
rect 18690 3952 18696 3955
rect 18748 3952 18754 4004
rect 19981 3995 20039 4001
rect 19981 3992 19993 3995
rect 19720 3964 19993 3992
rect 19720 3924 19748 3964
rect 19981 3961 19993 3964
rect 20027 3992 20039 3995
rect 20824 3992 20852 4032
rect 21634 4020 21640 4032
rect 21692 4020 21698 4072
rect 22554 4060 22560 4072
rect 22515 4032 22560 4060
rect 22554 4020 22560 4032
rect 22612 4020 22618 4072
rect 20027 3964 20852 3992
rect 20892 3995 20950 4001
rect 20027 3961 20039 3964
rect 19981 3955 20039 3961
rect 20892 3961 20904 3995
rect 20938 3992 20950 3995
rect 21542 3992 21548 4004
rect 20938 3964 21548 3992
rect 20938 3961 20950 3964
rect 20892 3955 20950 3961
rect 21542 3952 21548 3964
rect 21600 3952 21606 4004
rect 22649 3995 22707 4001
rect 22649 3992 22661 3995
rect 22066 3964 22661 3992
rect 16868 3896 19748 3924
rect 19797 3927 19855 3933
rect 19797 3893 19809 3927
rect 19843 3924 19855 3927
rect 20070 3924 20076 3936
rect 19843 3896 20076 3924
rect 19843 3893 19855 3896
rect 19797 3887 19855 3893
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20806 3884 20812 3936
rect 20864 3924 20870 3936
rect 21174 3924 21180 3936
rect 20864 3896 21180 3924
rect 20864 3884 20870 3896
rect 21174 3884 21180 3896
rect 21232 3884 21238 3936
rect 21726 3884 21732 3936
rect 21784 3924 21790 3936
rect 22066 3924 22094 3964
rect 22649 3961 22661 3964
rect 22695 3961 22707 3995
rect 22649 3955 22707 3961
rect 21784 3896 22094 3924
rect 23109 3927 23167 3933
rect 21784 3884 21790 3896
rect 23109 3893 23121 3927
rect 23155 3924 23167 3927
rect 23290 3924 23296 3936
rect 23155 3896 23296 3924
rect 23155 3893 23167 3896
rect 23109 3887 23167 3893
rect 23290 3884 23296 3896
rect 23348 3924 23354 3936
rect 23569 3927 23627 3933
rect 23569 3924 23581 3927
rect 23348 3896 23581 3924
rect 23348 3884 23354 3896
rect 23569 3893 23581 3896
rect 23615 3893 23627 3927
rect 23569 3887 23627 3893
rect 1104 3834 23460 3856
rect 1104 3782 8446 3834
rect 8498 3782 8510 3834
rect 8562 3782 8574 3834
rect 8626 3782 8638 3834
rect 8690 3782 15910 3834
rect 15962 3782 15974 3834
rect 16026 3782 16038 3834
rect 16090 3782 16102 3834
rect 16154 3782 23460 3834
rect 1104 3760 23460 3782
rect 16393 3723 16451 3729
rect 16393 3689 16405 3723
rect 16439 3720 16451 3723
rect 16439 3692 18644 3720
rect 16439 3689 16451 3692
rect 16393 3683 16451 3689
rect 3329 3655 3387 3661
rect 3329 3621 3341 3655
rect 3375 3652 3387 3655
rect 4062 3652 4068 3664
rect 3375 3624 4068 3652
rect 3375 3621 3387 3624
rect 3329 3615 3387 3621
rect 4062 3612 4068 3624
rect 4120 3612 4126 3664
rect 17620 3655 17678 3661
rect 17620 3621 17632 3655
rect 17666 3652 17678 3655
rect 18322 3652 18328 3664
rect 17666 3624 18328 3652
rect 17666 3621 17678 3624
rect 17620 3615 17678 3621
rect 18322 3612 18328 3624
rect 18380 3612 18386 3664
rect 18616 3652 18644 3692
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 19337 3723 19395 3729
rect 19337 3720 19349 3723
rect 18748 3692 19349 3720
rect 18748 3680 18754 3692
rect 19337 3689 19349 3692
rect 19383 3689 19395 3723
rect 20346 3720 20352 3732
rect 19337 3683 19395 3689
rect 19720 3692 20352 3720
rect 19720 3661 19748 3692
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 20714 3680 20720 3732
rect 20772 3720 20778 3732
rect 20898 3720 20904 3732
rect 20772 3692 20904 3720
rect 20772 3680 20778 3692
rect 20898 3680 20904 3692
rect 20956 3720 20962 3732
rect 21361 3723 21419 3729
rect 21361 3720 21373 3723
rect 20956 3692 21373 3720
rect 20956 3680 20962 3692
rect 21361 3689 21373 3692
rect 21407 3689 21419 3723
rect 21361 3683 21419 3689
rect 22554 3680 22560 3732
rect 22612 3720 22618 3732
rect 22833 3723 22891 3729
rect 22833 3720 22845 3723
rect 22612 3692 22845 3720
rect 22612 3680 22618 3692
rect 22833 3689 22845 3692
rect 22879 3689 22891 3723
rect 22833 3683 22891 3689
rect 22925 3723 22983 3729
rect 22925 3689 22937 3723
rect 22971 3720 22983 3723
rect 23014 3720 23020 3732
rect 22971 3692 23020 3720
rect 22971 3689 22983 3692
rect 22925 3683 22983 3689
rect 23014 3680 23020 3692
rect 23072 3680 23078 3732
rect 19705 3655 19763 3661
rect 19705 3652 19717 3655
rect 18616 3624 19717 3652
rect 19705 3621 19717 3624
rect 19751 3621 19763 3655
rect 19886 3652 19892 3664
rect 19847 3624 19892 3652
rect 19705 3615 19763 3621
rect 19886 3612 19892 3624
rect 19944 3612 19950 3664
rect 20254 3661 20260 3664
rect 20248 3615 20260 3661
rect 20312 3652 20318 3664
rect 21082 3652 21088 3664
rect 20312 3624 21088 3652
rect 20254 3612 20260 3615
rect 20312 3612 20318 3624
rect 21082 3612 21088 3624
rect 21140 3612 21146 3664
rect 22738 3652 22744 3664
rect 21468 3624 22744 3652
rect 2685 3587 2743 3593
rect 2685 3553 2697 3587
rect 2731 3584 2743 3587
rect 2731 3556 3740 3584
rect 2731 3553 2743 3556
rect 2685 3547 2743 3553
rect 3712 3392 3740 3556
rect 17770 3544 17776 3596
rect 17828 3584 17834 3596
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 17828 3556 17877 3584
rect 17828 3544 17834 3556
rect 17865 3553 17877 3556
rect 17911 3584 17923 3587
rect 17957 3587 18015 3593
rect 17957 3584 17969 3587
rect 17911 3556 17969 3584
rect 17911 3553 17923 3556
rect 17865 3547 17923 3553
rect 17957 3553 17969 3556
rect 18003 3553 18015 3587
rect 17957 3547 18015 3553
rect 18224 3587 18282 3593
rect 18224 3553 18236 3587
rect 18270 3584 18282 3587
rect 18506 3584 18512 3596
rect 18270 3556 18512 3584
rect 18270 3553 18282 3556
rect 18224 3547 18282 3553
rect 18506 3544 18512 3556
rect 18564 3584 18570 3596
rect 19150 3584 19156 3596
rect 18564 3556 19156 3584
rect 18564 3544 18570 3556
rect 19150 3544 19156 3556
rect 19208 3544 19214 3596
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 19981 3587 20039 3593
rect 19981 3584 19993 3587
rect 19576 3556 19993 3584
rect 19576 3544 19582 3556
rect 19981 3553 19993 3556
rect 20027 3584 20039 3587
rect 20622 3584 20628 3596
rect 20027 3556 20628 3584
rect 20027 3553 20039 3556
rect 19981 3547 20039 3553
rect 20622 3544 20628 3556
rect 20680 3584 20686 3596
rect 20806 3584 20812 3596
rect 20680 3556 20812 3584
rect 20680 3544 20686 3556
rect 20806 3544 20812 3556
rect 20864 3584 20870 3596
rect 21468 3593 21496 3624
rect 22738 3612 22744 3624
rect 22796 3612 22802 3664
rect 21726 3593 21732 3596
rect 21453 3587 21511 3593
rect 21453 3584 21465 3587
rect 20864 3556 21465 3584
rect 20864 3544 20870 3556
rect 21453 3553 21465 3556
rect 21499 3553 21511 3587
rect 21720 3584 21732 3593
rect 21687 3556 21732 3584
rect 21453 3547 21511 3553
rect 21720 3547 21732 3556
rect 21726 3544 21732 3547
rect 21784 3544 21790 3596
rect 22094 3544 22100 3596
rect 22152 3584 22158 3596
rect 23109 3587 23167 3593
rect 23109 3584 23121 3587
rect 22152 3556 23121 3584
rect 22152 3544 22158 3556
rect 23109 3553 23121 3556
rect 23155 3553 23167 3587
rect 23109 3547 23167 3553
rect 3694 3380 3700 3392
rect 3655 3352 3700 3380
rect 3694 3340 3700 3352
rect 3752 3340 3758 3392
rect 16485 3383 16543 3389
rect 16485 3349 16497 3383
rect 16531 3380 16543 3383
rect 17218 3380 17224 3392
rect 16531 3352 17224 3380
rect 16531 3349 16543 3352
rect 16485 3343 16543 3349
rect 17218 3340 17224 3352
rect 17276 3340 17282 3392
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 22830 3380 22836 3392
rect 19392 3352 22836 3380
rect 19392 3340 19398 3352
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 1104 3290 23460 3312
rect 1104 3238 4714 3290
rect 4766 3238 4778 3290
rect 4830 3238 4842 3290
rect 4894 3238 4906 3290
rect 4958 3238 12178 3290
rect 12230 3238 12242 3290
rect 12294 3238 12306 3290
rect 12358 3238 12370 3290
rect 12422 3238 19642 3290
rect 19694 3238 19706 3290
rect 19758 3238 19770 3290
rect 19822 3238 19834 3290
rect 19886 3238 23460 3290
rect 1104 3216 23460 3238
rect 2409 3179 2467 3185
rect 2409 3145 2421 3179
rect 2455 3176 2467 3179
rect 3694 3176 3700 3188
rect 2455 3148 3700 3176
rect 2455 3145 2467 3148
rect 2409 3139 2467 3145
rect 1394 3108 1400 3120
rect 1355 3080 1400 3108
rect 1394 3068 1400 3080
rect 1452 3068 1458 3120
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2972 1639 2975
rect 1949 2975 2007 2981
rect 1949 2972 1961 2975
rect 1627 2944 1961 2972
rect 1627 2941 1639 2944
rect 1581 2935 1639 2941
rect 1949 2941 1961 2944
rect 1995 2941 2007 2975
rect 1949 2935 2007 2941
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2424 2972 2452 3139
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 16482 3136 16488 3188
rect 16540 3176 16546 3188
rect 18417 3179 18475 3185
rect 18417 3176 18429 3179
rect 16540 3148 18429 3176
rect 16540 3136 16546 3148
rect 18417 3145 18429 3148
rect 18463 3145 18475 3179
rect 19334 3176 19340 3188
rect 19295 3148 19340 3176
rect 18417 3139 18475 3145
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19429 3179 19487 3185
rect 19429 3145 19441 3179
rect 19475 3176 19487 3179
rect 20162 3176 20168 3188
rect 19475 3148 20168 3176
rect 19475 3145 19487 3148
rect 19429 3139 19487 3145
rect 20162 3136 20168 3148
rect 20220 3136 20226 3188
rect 20438 3136 20444 3188
rect 20496 3176 20502 3188
rect 20901 3179 20959 3185
rect 20496 3148 20852 3176
rect 20496 3136 20502 3148
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 20824 3108 20852 3148
rect 20901 3145 20913 3179
rect 20947 3176 20959 3179
rect 21174 3176 21180 3188
rect 20947 3148 21180 3176
rect 20947 3145 20959 3148
rect 20901 3139 20959 3145
rect 21174 3136 21180 3148
rect 21232 3136 21238 3188
rect 18012 3080 19472 3108
rect 20824 3080 21588 3108
rect 18012 3068 18018 3080
rect 19444 3052 19472 3080
rect 19058 3040 19064 3052
rect 19019 3012 19064 3040
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 19426 3000 19432 3052
rect 19484 3000 19490 3052
rect 21358 3000 21364 3052
rect 21416 3040 21422 3052
rect 21453 3043 21511 3049
rect 21453 3040 21465 3043
rect 21416 3012 21465 3040
rect 21416 3000 21422 3012
rect 21453 3009 21465 3012
rect 21499 3009 21511 3043
rect 21453 3003 21511 3009
rect 2271 2944 2452 2972
rect 2685 2975 2743 2981
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2685 2941 2697 2975
rect 2731 2972 2743 2975
rect 6086 2972 6092 2984
rect 2731 2944 2912 2972
rect 6047 2944 6092 2972
rect 2731 2941 2743 2944
rect 2685 2935 2743 2941
rect 2498 2836 2504 2848
rect 2459 2808 2504 2836
rect 2498 2796 2504 2808
rect 2556 2796 2562 2848
rect 2884 2845 2912 2944
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 16942 2972 16948 2984
rect 16903 2944 16948 2972
rect 16942 2932 16948 2944
rect 17000 2932 17006 2984
rect 17218 2981 17224 2984
rect 17212 2972 17224 2981
rect 17179 2944 17224 2972
rect 17212 2935 17224 2944
rect 17276 2972 17282 2984
rect 18877 2975 18935 2981
rect 18877 2972 18889 2975
rect 17276 2944 18889 2972
rect 17218 2932 17224 2935
rect 17276 2932 17282 2944
rect 18877 2941 18889 2944
rect 18923 2941 18935 2975
rect 19076 2972 19104 3000
rect 20254 2972 20260 2984
rect 19076 2944 20260 2972
rect 18877 2935 18935 2941
rect 20254 2932 20260 2944
rect 20312 2932 20318 2984
rect 20806 2972 20812 2984
rect 20767 2944 20812 2972
rect 20806 2932 20812 2944
rect 20864 2932 20870 2984
rect 20990 2932 20996 2984
rect 21048 2972 21054 2984
rect 21269 2975 21327 2981
rect 21269 2972 21281 2975
rect 21048 2944 21281 2972
rect 21048 2932 21054 2944
rect 21269 2941 21281 2944
rect 21315 2941 21327 2975
rect 21560 2972 21588 3080
rect 23569 3043 23627 3049
rect 23569 3040 23581 3043
rect 22664 3012 23581 3040
rect 22664 2981 22692 3012
rect 23569 3009 23581 3012
rect 23615 3009 23627 3043
rect 23569 3003 23627 3009
rect 21821 2975 21879 2981
rect 21821 2972 21833 2975
rect 21560 2944 21833 2972
rect 21269 2935 21327 2941
rect 21821 2941 21833 2944
rect 21867 2941 21879 2975
rect 21821 2935 21879 2941
rect 22649 2975 22707 2981
rect 22649 2941 22661 2975
rect 22695 2941 22707 2975
rect 22649 2935 22707 2941
rect 22830 2932 22836 2984
rect 22888 2972 22894 2984
rect 22925 2975 22983 2981
rect 22925 2972 22937 2975
rect 22888 2944 22937 2972
rect 22888 2932 22894 2944
rect 22925 2941 22937 2944
rect 22971 2941 22983 2975
rect 22925 2935 22983 2941
rect 3694 2864 3700 2916
rect 3752 2904 3758 2916
rect 18230 2904 18236 2916
rect 3752 2876 18236 2904
rect 3752 2864 3758 2876
rect 18230 2864 18236 2876
rect 18288 2864 18294 2916
rect 18785 2907 18843 2913
rect 18785 2904 18797 2907
rect 18340 2876 18797 2904
rect 18340 2848 18368 2876
rect 18785 2873 18797 2876
rect 18831 2873 18843 2907
rect 18785 2867 18843 2873
rect 19242 2864 19248 2916
rect 19300 2904 19306 2916
rect 20438 2904 20444 2916
rect 19300 2876 20444 2904
rect 19300 2864 19306 2876
rect 20438 2864 20444 2876
rect 20496 2864 20502 2916
rect 20564 2907 20622 2913
rect 20564 2873 20576 2907
rect 20610 2904 20622 2907
rect 21008 2904 21036 2932
rect 20610 2876 21036 2904
rect 20610 2873 20622 2876
rect 20564 2867 20622 2873
rect 22002 2864 22008 2916
rect 22060 2904 22066 2916
rect 22373 2907 22431 2913
rect 22373 2904 22385 2907
rect 22060 2876 22385 2904
rect 22060 2864 22066 2876
rect 22373 2873 22385 2876
rect 22419 2873 22431 2907
rect 22373 2867 22431 2873
rect 2869 2839 2927 2845
rect 2869 2805 2881 2839
rect 2915 2836 2927 2839
rect 10686 2836 10692 2848
rect 2915 2808 10692 2836
rect 2915 2805 2927 2808
rect 2869 2799 2927 2805
rect 10686 2796 10692 2808
rect 10744 2836 10750 2848
rect 17954 2836 17960 2848
rect 10744 2808 17960 2836
rect 10744 2796 10750 2808
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 18322 2836 18328 2848
rect 18235 2808 18328 2836
rect 18322 2796 18328 2808
rect 18380 2796 18386 2848
rect 20070 2796 20076 2848
rect 20128 2836 20134 2848
rect 21361 2839 21419 2845
rect 21361 2836 21373 2839
rect 20128 2808 21373 2836
rect 20128 2796 20134 2808
rect 21361 2805 21373 2808
rect 21407 2805 21419 2839
rect 21910 2836 21916 2848
rect 21871 2808 21916 2836
rect 21361 2799 21419 2805
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 23014 2836 23020 2848
rect 22975 2808 23020 2836
rect 23014 2796 23020 2808
rect 23072 2796 23078 2848
rect 1104 2746 23460 2768
rect 1104 2694 8446 2746
rect 8498 2694 8510 2746
rect 8562 2694 8574 2746
rect 8626 2694 8638 2746
rect 8690 2694 15910 2746
rect 15962 2694 15974 2746
rect 16026 2694 16038 2746
rect 16090 2694 16102 2746
rect 16154 2694 23460 2746
rect 1104 2672 23460 2694
rect 10686 2632 10692 2644
rect 10647 2604 10692 2632
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 18506 2592 18512 2644
rect 18564 2632 18570 2644
rect 18601 2635 18659 2641
rect 18601 2632 18613 2635
rect 18564 2604 18613 2632
rect 18564 2592 18570 2604
rect 18601 2601 18613 2604
rect 18647 2601 18659 2635
rect 19150 2632 19156 2644
rect 19111 2604 19156 2632
rect 18601 2595 18659 2601
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 22462 2632 22468 2644
rect 19751 2604 22468 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 22557 2635 22615 2641
rect 22557 2601 22569 2635
rect 22603 2632 22615 2635
rect 22646 2632 22652 2644
rect 22603 2604 22652 2632
rect 22603 2601 22615 2604
rect 22557 2595 22615 2601
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 2225 2567 2283 2573
rect 2225 2533 2237 2567
rect 2271 2564 2283 2567
rect 2498 2564 2504 2576
rect 2271 2536 2504 2564
rect 2271 2533 2283 2536
rect 2225 2527 2283 2533
rect 2498 2524 2504 2536
rect 2556 2524 2562 2576
rect 6086 2524 6092 2576
rect 6144 2564 6150 2576
rect 6273 2567 6331 2573
rect 6273 2564 6285 2567
rect 6144 2536 6285 2564
rect 6144 2524 6150 2536
rect 6273 2533 6285 2536
rect 6319 2533 6331 2567
rect 6273 2527 6331 2533
rect 10413 2567 10471 2573
rect 10413 2533 10425 2567
rect 10459 2564 10471 2567
rect 10704 2564 10732 2592
rect 10459 2536 10732 2564
rect 17488 2567 17546 2573
rect 10459 2533 10471 2536
rect 10413 2527 10471 2533
rect 17488 2533 17500 2567
rect 17534 2564 17546 2567
rect 18322 2564 18328 2576
rect 17534 2536 18328 2564
rect 17534 2533 17546 2536
rect 17488 2527 17546 2533
rect 18322 2524 18328 2536
rect 18380 2524 18386 2576
rect 22002 2564 22008 2576
rect 19536 2536 22008 2564
rect 14737 2499 14795 2505
rect 14737 2465 14749 2499
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 2038 2360 2044 2372
rect 1999 2332 2044 2360
rect 2038 2320 2044 2332
rect 2096 2320 2102 2372
rect 6086 2360 6092 2372
rect 6047 2332 6092 2360
rect 6086 2320 6092 2332
rect 6144 2320 6150 2372
rect 10226 2360 10232 2372
rect 10187 2332 10232 2360
rect 10226 2320 10232 2332
rect 10284 2320 10290 2372
rect 14274 2252 14280 2304
rect 14332 2292 14338 2304
rect 14752 2292 14780 2459
rect 16942 2456 16948 2508
rect 17000 2496 17006 2508
rect 17221 2499 17279 2505
rect 17221 2496 17233 2499
rect 17000 2468 17233 2496
rect 17000 2456 17006 2468
rect 17221 2465 17233 2468
rect 17267 2496 17279 2499
rect 17770 2496 17776 2508
rect 17267 2468 17776 2496
rect 17267 2465 17279 2468
rect 17221 2459 17279 2465
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 19536 2505 19564 2536
rect 22002 2524 22008 2536
rect 22060 2524 22066 2576
rect 22925 2567 22983 2573
rect 22112 2536 22784 2564
rect 18877 2499 18935 2505
rect 18877 2465 18889 2499
rect 18923 2465 18935 2499
rect 18877 2459 18935 2465
rect 19521 2499 19579 2505
rect 19521 2465 19533 2499
rect 19567 2465 19579 2499
rect 19978 2496 19984 2508
rect 19939 2468 19984 2496
rect 19521 2459 19579 2465
rect 18414 2320 18420 2372
rect 18472 2360 18478 2372
rect 18892 2360 18920 2459
rect 19978 2456 19984 2468
rect 20036 2456 20042 2508
rect 20346 2496 20352 2508
rect 20307 2468 20352 2496
rect 20346 2456 20352 2468
rect 20404 2456 20410 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 20714 2496 20720 2508
rect 20671 2468 20720 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 20714 2456 20720 2468
rect 20772 2456 20778 2508
rect 20898 2505 20904 2508
rect 20892 2496 20904 2505
rect 20859 2468 20904 2496
rect 20892 2459 20904 2468
rect 20898 2456 20904 2459
rect 20956 2456 20962 2508
rect 21450 2456 21456 2508
rect 21508 2496 21514 2508
rect 22112 2496 22140 2536
rect 21508 2468 22140 2496
rect 21508 2456 21514 2468
rect 22186 2456 22192 2508
rect 22244 2496 22250 2508
rect 22756 2505 22784 2536
rect 22925 2533 22937 2567
rect 22971 2564 22983 2567
rect 23198 2564 23204 2576
rect 22971 2536 23204 2564
rect 22971 2533 22983 2536
rect 22925 2527 22983 2533
rect 23198 2524 23204 2536
rect 23256 2524 23262 2576
rect 22741 2499 22799 2505
rect 22244 2468 22508 2496
rect 22244 2456 22250 2468
rect 20530 2428 20536 2440
rect 20491 2400 20536 2428
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 22002 2388 22008 2440
rect 22060 2428 22066 2440
rect 22373 2431 22431 2437
rect 22373 2428 22385 2431
rect 22060 2400 22385 2428
rect 22060 2388 22066 2400
rect 22373 2397 22385 2400
rect 22419 2397 22431 2431
rect 22480 2428 22508 2468
rect 22741 2465 22753 2499
rect 22787 2465 22799 2499
rect 22741 2459 22799 2465
rect 22830 2428 22836 2440
rect 22480 2400 22836 2428
rect 22373 2391 22431 2397
rect 22830 2388 22836 2400
rect 22888 2388 22894 2440
rect 18969 2363 19027 2369
rect 18969 2360 18981 2363
rect 18472 2332 18981 2360
rect 18472 2320 18478 2332
rect 18969 2329 18981 2332
rect 19015 2329 19027 2363
rect 20346 2360 20352 2372
rect 18969 2323 19027 2329
rect 19260 2332 20352 2360
rect 14829 2295 14887 2301
rect 14829 2292 14841 2295
rect 14332 2264 14841 2292
rect 14332 2252 14338 2264
rect 14829 2261 14841 2264
rect 14875 2261 14887 2295
rect 14829 2255 14887 2261
rect 17037 2295 17095 2301
rect 17037 2261 17049 2295
rect 17083 2292 17095 2295
rect 19260 2292 19288 2332
rect 20346 2320 20352 2332
rect 20404 2320 20410 2372
rect 23109 2363 23167 2369
rect 23109 2329 23121 2363
rect 23155 2360 23167 2363
rect 23569 2363 23627 2369
rect 23569 2360 23581 2363
rect 23155 2332 23581 2360
rect 23155 2329 23167 2332
rect 23109 2323 23167 2329
rect 23569 2329 23581 2332
rect 23615 2329 23627 2363
rect 23569 2323 23627 2329
rect 19426 2292 19432 2304
rect 17083 2264 19288 2292
rect 19387 2264 19432 2292
rect 17083 2261 17095 2264
rect 17037 2255 17095 2261
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 20165 2295 20223 2301
rect 20165 2261 20177 2295
rect 20211 2292 20223 2295
rect 21266 2292 21272 2304
rect 20211 2264 21272 2292
rect 20211 2261 20223 2264
rect 20165 2255 20223 2261
rect 21266 2252 21272 2264
rect 21324 2252 21330 2304
rect 21726 2252 21732 2304
rect 21784 2292 21790 2304
rect 22005 2295 22063 2301
rect 22005 2292 22017 2295
rect 21784 2264 22017 2292
rect 21784 2252 21790 2264
rect 22005 2261 22017 2264
rect 22051 2261 22063 2295
rect 22005 2255 22063 2261
rect 1104 2202 23460 2224
rect 1104 2150 4714 2202
rect 4766 2150 4778 2202
rect 4830 2150 4842 2202
rect 4894 2150 4906 2202
rect 4958 2150 12178 2202
rect 12230 2150 12242 2202
rect 12294 2150 12306 2202
rect 12358 2150 12370 2202
rect 12422 2150 19642 2202
rect 19694 2150 19706 2202
rect 19758 2150 19770 2202
rect 19822 2150 19834 2202
rect 19886 2150 23460 2202
rect 1104 2128 23460 2150
rect 19426 2048 19432 2100
rect 19484 2088 19490 2100
rect 22186 2088 22192 2100
rect 19484 2060 22192 2088
rect 19484 2048 19490 2060
rect 22186 2048 22192 2060
rect 22244 2048 22250 2100
rect 20346 1980 20352 2032
rect 20404 2020 20410 2032
rect 23474 2020 23480 2032
rect 20404 1992 23480 2020
rect 20404 1980 20410 1992
rect 23474 1980 23480 1992
rect 23532 1980 23538 2032
rect 23566 1408 23572 1420
rect 23527 1380 23572 1408
rect 23566 1368 23572 1380
rect 23624 1368 23630 1420
<< via1 >>
rect 10140 22516 10192 22568
rect 10600 22516 10652 22568
rect 11612 22516 11664 22568
rect 15108 22516 15160 22568
rect 16212 22516 16264 22568
rect 9864 22448 9916 22500
rect 17408 22448 17460 22500
rect 18420 22448 18472 22500
rect 5448 22380 5500 22432
rect 5908 22380 5960 22432
rect 6644 22380 6696 22432
rect 9956 22380 10008 22432
rect 12256 22380 12308 22432
rect 15016 22380 15068 22432
rect 18880 22380 18932 22432
rect 8446 22278 8498 22330
rect 8510 22278 8562 22330
rect 8574 22278 8626 22330
rect 8638 22278 8690 22330
rect 15910 22278 15962 22330
rect 15974 22278 16026 22330
rect 16038 22278 16090 22330
rect 16102 22278 16154 22330
rect 5908 22108 5960 22160
rect 7472 22176 7524 22228
rect 11704 22176 11756 22228
rect 14464 22176 14516 22228
rect 15016 22176 15068 22228
rect 296 22040 348 22092
rect 1584 22083 1636 22092
rect 1584 22049 1593 22083
rect 1593 22049 1627 22083
rect 1627 22049 1636 22083
rect 1584 22040 1636 22049
rect 1952 22083 2004 22092
rect 1952 22049 1961 22083
rect 1961 22049 1995 22083
rect 1995 22049 2004 22083
rect 1952 22040 2004 22049
rect 2320 22083 2372 22092
rect 2320 22049 2329 22083
rect 2329 22049 2363 22083
rect 2363 22049 2372 22083
rect 2320 22040 2372 22049
rect 2688 22083 2740 22092
rect 2688 22049 2697 22083
rect 2697 22049 2731 22083
rect 2731 22049 2740 22083
rect 2688 22040 2740 22049
rect 2872 22083 2924 22092
rect 2872 22049 2881 22083
rect 2881 22049 2915 22083
rect 2915 22049 2924 22083
rect 2872 22040 2924 22049
rect 3332 22040 3384 22092
rect 940 21972 992 22024
rect 2228 21972 2280 22024
rect 2596 21972 2648 22024
rect 4160 22040 4212 22092
rect 4804 22083 4856 22092
rect 4804 22049 4813 22083
rect 4813 22049 4847 22083
rect 4847 22049 4856 22083
rect 4804 22040 4856 22049
rect 5356 22083 5408 22092
rect 4528 21972 4580 22024
rect 5356 22049 5365 22083
rect 5365 22049 5399 22083
rect 5399 22049 5408 22083
rect 5356 22040 5408 22049
rect 8300 22108 8352 22160
rect 9588 22108 9640 22160
rect 10784 22151 10836 22160
rect 1676 21904 1728 21956
rect 3516 21904 3568 21956
rect 2412 21836 2464 21888
rect 5356 21836 5408 21888
rect 5448 21836 5500 21888
rect 6276 22040 6328 22092
rect 7012 22083 7064 22092
rect 7012 22049 7021 22083
rect 7021 22049 7055 22083
rect 7055 22049 7064 22083
rect 7012 22040 7064 22049
rect 7380 22083 7432 22092
rect 7380 22049 7389 22083
rect 7389 22049 7423 22083
rect 7423 22049 7432 22083
rect 7380 22040 7432 22049
rect 7840 22040 7892 22092
rect 7564 22015 7616 22024
rect 7564 21981 7573 22015
rect 7573 21981 7607 22015
rect 7607 21981 7616 22015
rect 7564 21972 7616 21981
rect 7748 22015 7800 22024
rect 7748 21981 7757 22015
rect 7757 21981 7791 22015
rect 7791 21981 7800 22015
rect 7748 21972 7800 21981
rect 7932 21972 7984 22024
rect 6092 21836 6144 21888
rect 6276 21879 6328 21888
rect 6276 21845 6285 21879
rect 6285 21845 6319 21879
rect 6319 21845 6328 21879
rect 6276 21836 6328 21845
rect 6552 21879 6604 21888
rect 6552 21845 6561 21879
rect 6561 21845 6595 21879
rect 6595 21845 6604 21879
rect 6552 21836 6604 21845
rect 6644 21836 6696 21888
rect 7104 21836 7156 21888
rect 8116 21904 8168 21956
rect 9680 22040 9732 22092
rect 10784 22117 10793 22151
rect 10793 22117 10827 22151
rect 10827 22117 10836 22151
rect 10784 22108 10836 22117
rect 13636 22108 13688 22160
rect 13820 22108 13872 22160
rect 18880 22219 18932 22228
rect 18880 22185 18889 22219
rect 18889 22185 18923 22219
rect 18923 22185 18932 22219
rect 18880 22176 18932 22185
rect 11612 22083 11664 22092
rect 11612 22049 11621 22083
rect 11621 22049 11655 22083
rect 11655 22049 11664 22083
rect 11612 22040 11664 22049
rect 11888 22040 11940 22092
rect 12256 22040 12308 22092
rect 12716 22083 12768 22092
rect 12716 22049 12725 22083
rect 12725 22049 12759 22083
rect 12759 22049 12768 22083
rect 12716 22040 12768 22049
rect 12808 22083 12860 22092
rect 12808 22049 12817 22083
rect 12817 22049 12851 22083
rect 12851 22049 12860 22083
rect 12808 22040 12860 22049
rect 12992 22040 13044 22092
rect 13176 22040 13228 22092
rect 14372 22083 14424 22092
rect 14372 22049 14381 22083
rect 14381 22049 14415 22083
rect 14415 22049 14424 22083
rect 14372 22040 14424 22049
rect 15016 22083 15068 22092
rect 8760 21972 8812 22024
rect 9128 21972 9180 22024
rect 9772 22015 9824 22024
rect 9772 21981 9781 22015
rect 9781 21981 9815 22015
rect 9815 21981 9824 22015
rect 9772 21972 9824 21981
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 10600 21972 10652 22024
rect 11060 21972 11112 22024
rect 13728 21972 13780 22024
rect 13912 22015 13964 22024
rect 13912 21981 13921 22015
rect 13921 21981 13955 22015
rect 13955 21981 13964 22015
rect 13912 21972 13964 21981
rect 10048 21904 10100 21956
rect 11428 21947 11480 21956
rect 11428 21913 11437 21947
rect 11437 21913 11471 21947
rect 11471 21913 11480 21947
rect 11428 21904 11480 21913
rect 13176 21904 13228 21956
rect 15016 22049 15025 22083
rect 15025 22049 15059 22083
rect 15059 22049 15068 22083
rect 15016 22040 15068 22049
rect 15384 22083 15436 22092
rect 15384 22049 15393 22083
rect 15393 22049 15427 22083
rect 15427 22049 15436 22083
rect 15384 22040 15436 22049
rect 16212 22108 16264 22160
rect 17408 22151 17460 22160
rect 17408 22117 17417 22151
rect 17417 22117 17451 22151
rect 17451 22117 17460 22151
rect 17408 22108 17460 22117
rect 17960 22108 18012 22160
rect 16028 22040 16080 22092
rect 16488 22083 16540 22092
rect 16488 22049 16497 22083
rect 16497 22049 16531 22083
rect 16531 22049 16540 22083
rect 16488 22040 16540 22049
rect 16580 22083 16632 22092
rect 16580 22049 16589 22083
rect 16589 22049 16623 22083
rect 16623 22049 16632 22083
rect 17040 22083 17092 22092
rect 16580 22040 16632 22049
rect 17040 22049 17049 22083
rect 17049 22049 17083 22083
rect 17083 22049 17092 22083
rect 17040 22040 17092 22049
rect 19064 22040 19116 22092
rect 20168 22108 20220 22160
rect 22284 22176 22336 22228
rect 18788 21972 18840 22024
rect 19340 22040 19392 22092
rect 19432 22040 19484 22092
rect 19616 22040 19668 22092
rect 20076 22083 20128 22092
rect 20076 22049 20085 22083
rect 20085 22049 20119 22083
rect 20119 22049 20128 22083
rect 20076 22040 20128 22049
rect 20260 22083 20312 22092
rect 20260 22049 20269 22083
rect 20269 22049 20303 22083
rect 20303 22049 20312 22083
rect 20260 22040 20312 22049
rect 20812 22083 20864 22092
rect 20812 22049 20821 22083
rect 20821 22049 20855 22083
rect 20855 22049 20864 22083
rect 20812 22040 20864 22049
rect 20904 22083 20956 22092
rect 20904 22049 20913 22083
rect 20913 22049 20947 22083
rect 20947 22049 20956 22083
rect 21088 22083 21140 22092
rect 20904 22040 20956 22049
rect 21088 22049 21097 22083
rect 21097 22049 21131 22083
rect 21131 22049 21140 22083
rect 21088 22040 21140 22049
rect 21456 22083 21508 22092
rect 21456 22049 21465 22083
rect 21465 22049 21499 22083
rect 21499 22049 21508 22083
rect 21456 22040 21508 22049
rect 21640 22083 21692 22092
rect 21640 22049 21649 22083
rect 21649 22049 21683 22083
rect 21683 22049 21692 22083
rect 21640 22040 21692 22049
rect 21824 22083 21876 22092
rect 21824 22049 21833 22083
rect 21833 22049 21867 22083
rect 21867 22049 21876 22083
rect 21824 22040 21876 22049
rect 21916 22040 21968 22092
rect 23112 22083 23164 22092
rect 23112 22049 23121 22083
rect 23121 22049 23155 22083
rect 23155 22049 23164 22083
rect 23112 22040 23164 22049
rect 19248 21972 19300 22024
rect 21548 21972 21600 22024
rect 22008 21972 22060 22024
rect 17684 21904 17736 21956
rect 22192 21904 22244 21956
rect 9864 21836 9916 21888
rect 11244 21879 11296 21888
rect 11244 21845 11253 21879
rect 11253 21845 11287 21879
rect 11287 21845 11296 21879
rect 11244 21836 11296 21845
rect 11612 21836 11664 21888
rect 12532 21879 12584 21888
rect 12532 21845 12541 21879
rect 12541 21845 12575 21879
rect 12575 21845 12584 21879
rect 12532 21836 12584 21845
rect 13084 21836 13136 21888
rect 13268 21879 13320 21888
rect 13268 21845 13277 21879
rect 13277 21845 13311 21879
rect 13311 21845 13320 21879
rect 13268 21836 13320 21845
rect 14004 21836 14056 21888
rect 14740 21879 14792 21888
rect 14740 21845 14749 21879
rect 14749 21845 14783 21879
rect 14783 21845 14792 21879
rect 14740 21836 14792 21845
rect 15292 21836 15344 21888
rect 15476 21836 15528 21888
rect 16764 21879 16816 21888
rect 16764 21845 16773 21879
rect 16773 21845 16807 21879
rect 16807 21845 16816 21879
rect 16764 21836 16816 21845
rect 16948 21836 17000 21888
rect 18972 21836 19024 21888
rect 22100 21836 22152 21888
rect 4714 21734 4766 21786
rect 4778 21734 4830 21786
rect 4842 21734 4894 21786
rect 4906 21734 4958 21786
rect 12178 21734 12230 21786
rect 12242 21734 12294 21786
rect 12306 21734 12358 21786
rect 12370 21734 12422 21786
rect 19642 21734 19694 21786
rect 19706 21734 19758 21786
rect 19770 21734 19822 21786
rect 19834 21734 19886 21786
rect 1584 21632 1636 21684
rect 1952 21632 2004 21684
rect 3332 21632 3384 21684
rect 6000 21632 6052 21684
rect 6736 21675 6788 21684
rect 6736 21641 6745 21675
rect 6745 21641 6779 21675
rect 6779 21641 6788 21675
rect 6736 21632 6788 21641
rect 7932 21632 7984 21684
rect 8116 21632 8168 21684
rect 9864 21632 9916 21684
rect 10600 21632 10652 21684
rect 11796 21632 11848 21684
rect 12992 21632 13044 21684
rect 2504 21607 2556 21616
rect 1584 21471 1636 21480
rect 1584 21437 1593 21471
rect 1593 21437 1627 21471
rect 1627 21437 1636 21471
rect 2504 21573 2513 21607
rect 2513 21573 2547 21607
rect 2547 21573 2556 21607
rect 2504 21564 2556 21573
rect 4160 21564 4212 21616
rect 2136 21496 2188 21548
rect 1584 21428 1636 21437
rect 2412 21428 2464 21480
rect 6920 21496 6972 21548
rect 9036 21564 9088 21616
rect 10876 21564 10928 21616
rect 8576 21496 8628 21548
rect 4252 21471 4304 21480
rect 3424 21360 3476 21412
rect 4252 21437 4261 21471
rect 4261 21437 4295 21471
rect 4295 21437 4304 21471
rect 4252 21428 4304 21437
rect 4436 21471 4488 21480
rect 4436 21437 4445 21471
rect 4445 21437 4479 21471
rect 4479 21437 4488 21471
rect 4436 21428 4488 21437
rect 4528 21428 4580 21480
rect 6644 21471 6696 21480
rect 5264 21360 5316 21412
rect 5816 21335 5868 21344
rect 5816 21301 5825 21335
rect 5825 21301 5859 21335
rect 5859 21301 5868 21335
rect 5816 21292 5868 21301
rect 6644 21437 6653 21471
rect 6653 21437 6687 21471
rect 6687 21437 6696 21471
rect 6644 21428 6696 21437
rect 8392 21428 8444 21480
rect 8760 21428 8812 21480
rect 10968 21496 11020 21548
rect 10692 21428 10744 21480
rect 11612 21496 11664 21548
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 15384 21632 15436 21684
rect 14648 21607 14700 21616
rect 14648 21573 14657 21607
rect 14657 21573 14691 21607
rect 14691 21573 14700 21607
rect 14648 21564 14700 21573
rect 16396 21632 16448 21684
rect 16580 21632 16632 21684
rect 18328 21632 18380 21684
rect 22836 21632 22888 21684
rect 16212 21607 16264 21616
rect 16212 21573 16221 21607
rect 16221 21573 16255 21607
rect 16255 21573 16264 21607
rect 16212 21564 16264 21573
rect 18052 21564 18104 21616
rect 20076 21564 20128 21616
rect 23480 21564 23532 21616
rect 11336 21428 11388 21480
rect 7840 21360 7892 21412
rect 8944 21403 8996 21412
rect 8944 21369 8953 21403
rect 8953 21369 8987 21403
rect 8987 21369 8996 21403
rect 8944 21360 8996 21369
rect 9128 21360 9180 21412
rect 10416 21360 10468 21412
rect 10968 21360 11020 21412
rect 12348 21428 12400 21480
rect 12900 21428 12952 21480
rect 14096 21428 14148 21480
rect 16028 21496 16080 21548
rect 12072 21403 12124 21412
rect 12072 21369 12106 21403
rect 12106 21369 12124 21403
rect 12072 21360 12124 21369
rect 11612 21292 11664 21344
rect 12900 21292 12952 21344
rect 13360 21360 13412 21412
rect 14280 21360 14332 21412
rect 15108 21360 15160 21412
rect 15292 21428 15344 21480
rect 16764 21496 16816 21548
rect 16948 21471 17000 21480
rect 16948 21437 16957 21471
rect 16957 21437 16991 21471
rect 16991 21437 17000 21471
rect 16948 21428 17000 21437
rect 18696 21496 18748 21548
rect 19248 21496 19300 21548
rect 23112 21539 23164 21548
rect 23112 21505 23121 21539
rect 23121 21505 23155 21539
rect 23155 21505 23164 21539
rect 23112 21496 23164 21505
rect 18604 21428 18656 21480
rect 20168 21428 20220 21480
rect 21640 21428 21692 21480
rect 17224 21403 17276 21412
rect 17224 21369 17258 21403
rect 17258 21369 17276 21403
rect 17224 21360 17276 21369
rect 17316 21360 17368 21412
rect 18880 21292 18932 21344
rect 19156 21360 19208 21412
rect 21088 21292 21140 21344
rect 21364 21335 21416 21344
rect 21364 21301 21373 21335
rect 21373 21301 21407 21335
rect 21407 21301 21416 21335
rect 21364 21292 21416 21301
rect 21548 21292 21600 21344
rect 22192 21335 22244 21344
rect 22192 21301 22201 21335
rect 22201 21301 22235 21335
rect 22235 21301 22244 21335
rect 22192 21292 22244 21301
rect 8446 21190 8498 21242
rect 8510 21190 8562 21242
rect 8574 21190 8626 21242
rect 8638 21190 8690 21242
rect 15910 21190 15962 21242
rect 15974 21190 16026 21242
rect 16038 21190 16090 21242
rect 16102 21190 16154 21242
rect 2320 21088 2372 21140
rect 2688 21088 2740 21140
rect 5264 21131 5316 21140
rect 5264 21097 5273 21131
rect 5273 21097 5307 21131
rect 5307 21097 5316 21131
rect 5264 21088 5316 21097
rect 5356 21088 5408 21140
rect 2596 21020 2648 21072
rect 4160 21063 4212 21072
rect 4160 21029 4194 21063
rect 4194 21029 4212 21063
rect 4160 21020 4212 21029
rect 5816 21020 5868 21072
rect 8760 21088 8812 21140
rect 8852 21088 8904 21140
rect 9312 21088 9364 21140
rect 2136 20952 2188 21004
rect 2872 20952 2924 21004
rect 3700 20995 3752 21004
rect 3700 20961 3709 20995
rect 3709 20961 3743 20995
rect 3743 20961 3752 20995
rect 3700 20952 3752 20961
rect 4436 20952 4488 21004
rect 6736 20952 6788 21004
rect 6644 20884 6696 20936
rect 1676 20859 1728 20868
rect 1676 20825 1685 20859
rect 1685 20825 1719 20859
rect 1719 20825 1728 20859
rect 1676 20816 1728 20825
rect 3424 20859 3476 20868
rect 3424 20825 3433 20859
rect 3433 20825 3467 20859
rect 3467 20825 3476 20859
rect 3424 20816 3476 20825
rect 8392 21020 8444 21072
rect 9588 21063 9640 21072
rect 9588 21029 9622 21063
rect 9622 21029 9640 21063
rect 9588 21020 9640 21029
rect 9772 21088 9824 21140
rect 11060 21131 11112 21140
rect 11060 21097 11069 21131
rect 11069 21097 11103 21131
rect 11103 21097 11112 21131
rect 11060 21088 11112 21097
rect 11336 21063 11388 21072
rect 11336 21029 11345 21063
rect 11345 21029 11379 21063
rect 11379 21029 11388 21063
rect 11336 21020 11388 21029
rect 13360 21131 13412 21140
rect 13360 21097 13369 21131
rect 13369 21097 13403 21131
rect 13403 21097 13412 21131
rect 13728 21131 13780 21140
rect 13360 21088 13412 21097
rect 13728 21097 13737 21131
rect 13737 21097 13771 21131
rect 13771 21097 13780 21131
rect 13728 21088 13780 21097
rect 13912 21131 13964 21140
rect 13912 21097 13921 21131
rect 13921 21097 13955 21131
rect 13955 21097 13964 21131
rect 13912 21088 13964 21097
rect 14096 21088 14148 21140
rect 12072 21020 12124 21072
rect 8392 20884 8444 20936
rect 10508 20952 10560 21004
rect 12348 20952 12400 21004
rect 12624 20995 12676 21004
rect 12624 20961 12642 20995
rect 12642 20961 12676 20995
rect 12900 20995 12952 21004
rect 12624 20952 12676 20961
rect 12900 20961 12909 20995
rect 12909 20961 12943 20995
rect 12943 20961 12952 20995
rect 12900 20952 12952 20961
rect 14004 21063 14056 21072
rect 14004 21029 14013 21063
rect 14013 21029 14047 21063
rect 14047 21029 14056 21063
rect 14004 21020 14056 21029
rect 14648 21063 14700 21072
rect 14648 21029 14682 21063
rect 14682 21029 14700 21063
rect 14648 21020 14700 21029
rect 15108 21088 15160 21140
rect 18604 21088 18656 21140
rect 18788 21131 18840 21140
rect 18788 21097 18797 21131
rect 18797 21097 18831 21131
rect 18831 21097 18840 21131
rect 18788 21088 18840 21097
rect 19064 21131 19116 21140
rect 19064 21097 19073 21131
rect 19073 21097 19107 21131
rect 19107 21097 19116 21131
rect 19064 21088 19116 21097
rect 19156 21088 19208 21140
rect 21456 21088 21508 21140
rect 22100 21088 22152 21140
rect 24124 21088 24176 21140
rect 15292 21020 15344 21072
rect 15660 21020 15712 21072
rect 15844 21020 15896 21072
rect 16396 21020 16448 21072
rect 14464 20952 14516 21004
rect 19432 21020 19484 21072
rect 18880 20952 18932 21004
rect 20444 20952 20496 21004
rect 22008 21020 22060 21072
rect 21180 20952 21232 21004
rect 21364 20952 21416 21004
rect 21732 20952 21784 21004
rect 22100 20952 22152 21004
rect 9036 20884 9088 20936
rect 13452 20884 13504 20936
rect 14096 20884 14148 20936
rect 15660 20884 15712 20936
rect 16948 20884 17000 20936
rect 18420 20884 18472 20936
rect 22284 20952 22336 21004
rect 4252 20748 4304 20800
rect 6460 20748 6512 20800
rect 6736 20791 6788 20800
rect 6736 20757 6745 20791
rect 6745 20757 6779 20791
rect 6779 20757 6788 20791
rect 6736 20748 6788 20757
rect 7564 20748 7616 20800
rect 8484 20748 8536 20800
rect 11336 20816 11388 20868
rect 11060 20748 11112 20800
rect 14188 20816 14240 20868
rect 18512 20816 18564 20868
rect 21180 20816 21232 20868
rect 21824 20816 21876 20868
rect 21916 20816 21968 20868
rect 22100 20816 22152 20868
rect 23480 20884 23532 20936
rect 22744 20859 22796 20868
rect 22744 20825 22753 20859
rect 22753 20825 22787 20859
rect 22787 20825 22796 20859
rect 22744 20816 22796 20825
rect 13360 20748 13412 20800
rect 15844 20748 15896 20800
rect 16580 20748 16632 20800
rect 17224 20791 17276 20800
rect 17224 20757 17233 20791
rect 17233 20757 17267 20791
rect 17267 20757 17276 20791
rect 17224 20748 17276 20757
rect 18972 20748 19024 20800
rect 23020 20791 23072 20800
rect 23020 20757 23029 20791
rect 23029 20757 23063 20791
rect 23063 20757 23072 20791
rect 23020 20748 23072 20757
rect 4714 20646 4766 20698
rect 4778 20646 4830 20698
rect 4842 20646 4894 20698
rect 4906 20646 4958 20698
rect 12178 20646 12230 20698
rect 12242 20646 12294 20698
rect 12306 20646 12358 20698
rect 12370 20646 12422 20698
rect 19642 20646 19694 20698
rect 19706 20646 19758 20698
rect 19770 20646 19822 20698
rect 19834 20646 19886 20698
rect 2872 20544 2924 20596
rect 2136 20340 2188 20392
rect 2872 20340 2924 20392
rect 6828 20544 6880 20596
rect 9588 20544 9640 20596
rect 10876 20544 10928 20596
rect 11336 20587 11388 20596
rect 11336 20553 11345 20587
rect 11345 20553 11379 20587
rect 11379 20553 11388 20587
rect 11336 20544 11388 20553
rect 12716 20544 12768 20596
rect 13636 20544 13688 20596
rect 16304 20544 16356 20596
rect 17960 20544 18012 20596
rect 18328 20544 18380 20596
rect 19248 20544 19300 20596
rect 19340 20544 19392 20596
rect 21640 20544 21692 20596
rect 22008 20587 22060 20596
rect 22008 20553 22017 20587
rect 22017 20553 22051 20587
rect 22051 20553 22060 20587
rect 22008 20544 22060 20553
rect 4436 20408 4488 20460
rect 4896 20451 4948 20460
rect 4896 20417 4905 20451
rect 4905 20417 4939 20451
rect 4939 20417 4948 20451
rect 4896 20408 4948 20417
rect 5816 20408 5868 20460
rect 6092 20408 6144 20460
rect 6644 20408 6696 20460
rect 4160 20340 4212 20392
rect 6920 20383 6972 20392
rect 6920 20349 6929 20383
rect 6929 20349 6963 20383
rect 6963 20349 6972 20383
rect 6920 20340 6972 20349
rect 7932 20340 7984 20392
rect 14924 20476 14976 20528
rect 1676 20272 1728 20324
rect 3700 20272 3752 20324
rect 6368 20272 6420 20324
rect 4068 20204 4120 20256
rect 4252 20204 4304 20256
rect 4620 20247 4672 20256
rect 4620 20213 4629 20247
rect 4629 20213 4663 20247
rect 4663 20213 4672 20247
rect 4620 20204 4672 20213
rect 4712 20204 4764 20256
rect 5724 20204 5776 20256
rect 5908 20247 5960 20256
rect 5908 20213 5917 20247
rect 5917 20213 5951 20247
rect 5951 20213 5960 20247
rect 5908 20204 5960 20213
rect 8760 20272 8812 20324
rect 10600 20383 10652 20392
rect 10600 20349 10609 20383
rect 10609 20349 10643 20383
rect 10643 20349 10652 20383
rect 10600 20340 10652 20349
rect 11520 20340 11572 20392
rect 12992 20340 13044 20392
rect 13268 20340 13320 20392
rect 10140 20272 10192 20324
rect 10232 20272 10284 20324
rect 10508 20272 10560 20324
rect 12808 20315 12860 20324
rect 12808 20281 12826 20315
rect 12826 20281 12860 20315
rect 12808 20272 12860 20281
rect 13452 20272 13504 20324
rect 14740 20408 14792 20460
rect 16212 20408 16264 20460
rect 14280 20383 14332 20392
rect 14280 20349 14289 20383
rect 14289 20349 14323 20383
rect 14323 20349 14332 20383
rect 14280 20340 14332 20349
rect 14648 20340 14700 20392
rect 15200 20340 15252 20392
rect 13820 20272 13872 20324
rect 6644 20247 6696 20256
rect 6644 20213 6653 20247
rect 6653 20213 6687 20247
rect 6687 20213 6696 20247
rect 6644 20204 6696 20213
rect 6736 20247 6788 20256
rect 6736 20213 6745 20247
rect 6745 20213 6779 20247
rect 6779 20213 6788 20247
rect 6736 20204 6788 20213
rect 6920 20204 6972 20256
rect 8300 20204 8352 20256
rect 9772 20204 9824 20256
rect 12624 20204 12676 20256
rect 12900 20204 12952 20256
rect 15016 20247 15068 20256
rect 15016 20213 15025 20247
rect 15025 20213 15059 20247
rect 15059 20213 15068 20247
rect 15016 20204 15068 20213
rect 16856 20272 16908 20324
rect 21548 20476 21600 20528
rect 18880 20451 18932 20460
rect 18880 20417 18889 20451
rect 18889 20417 18923 20451
rect 18923 20417 18932 20451
rect 18880 20408 18932 20417
rect 18972 20408 19024 20460
rect 18328 20272 18380 20324
rect 18788 20340 18840 20392
rect 20904 20340 20956 20392
rect 16212 20204 16264 20256
rect 16396 20247 16448 20256
rect 16396 20213 16405 20247
rect 16405 20213 16439 20247
rect 16439 20213 16448 20247
rect 21640 20340 21692 20392
rect 22192 20340 22244 20392
rect 22836 20315 22888 20324
rect 16396 20204 16448 20213
rect 18972 20204 19024 20256
rect 19064 20247 19116 20256
rect 19064 20213 19073 20247
rect 19073 20213 19107 20247
rect 19107 20213 19116 20247
rect 19524 20247 19576 20256
rect 19064 20204 19116 20213
rect 19524 20213 19533 20247
rect 19533 20213 19567 20247
rect 19567 20213 19576 20247
rect 19524 20204 19576 20213
rect 20076 20247 20128 20256
rect 20076 20213 20085 20247
rect 20085 20213 20119 20247
rect 20119 20213 20128 20247
rect 20076 20204 20128 20213
rect 20260 20204 20312 20256
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 21180 20247 21232 20256
rect 21180 20213 21189 20247
rect 21189 20213 21223 20247
rect 21223 20213 21232 20247
rect 21180 20204 21232 20213
rect 22100 20204 22152 20256
rect 22836 20281 22845 20315
rect 22845 20281 22879 20315
rect 22879 20281 22888 20315
rect 22836 20272 22888 20281
rect 8446 20102 8498 20154
rect 8510 20102 8562 20154
rect 8574 20102 8626 20154
rect 8638 20102 8690 20154
rect 15910 20102 15962 20154
rect 15974 20102 16026 20154
rect 16038 20102 16090 20154
rect 16102 20102 16154 20154
rect 1676 20000 1728 20052
rect 3700 20043 3752 20052
rect 3700 20009 3709 20043
rect 3709 20009 3743 20043
rect 3743 20009 3752 20043
rect 3700 20000 3752 20009
rect 4620 20000 4672 20052
rect 5632 20000 5684 20052
rect 6368 20043 6420 20052
rect 6368 20009 6377 20043
rect 6377 20009 6411 20043
rect 6411 20009 6420 20043
rect 6368 20000 6420 20009
rect 7840 20000 7892 20052
rect 8760 20043 8812 20052
rect 3056 19864 3108 19916
rect 4068 19932 4120 19984
rect 5724 19932 5776 19984
rect 3516 19907 3568 19916
rect 3516 19873 3525 19907
rect 3525 19873 3559 19907
rect 3559 19873 3568 19907
rect 3516 19864 3568 19873
rect 5172 19864 5224 19916
rect 2964 19839 3016 19848
rect 2964 19805 2973 19839
rect 2973 19805 3007 19839
rect 3007 19805 3016 19839
rect 2964 19796 3016 19805
rect 4528 19839 4580 19848
rect 4528 19805 4537 19839
rect 4537 19805 4571 19839
rect 4571 19805 4580 19839
rect 4528 19796 4580 19805
rect 4896 19839 4948 19848
rect 4896 19805 4905 19839
rect 4905 19805 4939 19839
rect 4939 19805 4948 19839
rect 4896 19796 4948 19805
rect 6736 19932 6788 19984
rect 8300 19932 8352 19984
rect 8760 20009 8769 20043
rect 8769 20009 8803 20043
rect 8803 20009 8812 20043
rect 8760 20000 8812 20009
rect 10508 20000 10560 20052
rect 10784 20000 10836 20052
rect 11980 20043 12032 20052
rect 11980 20009 11989 20043
rect 11989 20009 12023 20043
rect 12023 20009 12032 20043
rect 11980 20000 12032 20009
rect 12900 20043 12952 20052
rect 9864 19932 9916 19984
rect 11060 19932 11112 19984
rect 12900 20009 12909 20043
rect 12909 20009 12943 20043
rect 12943 20009 12952 20043
rect 12900 20000 12952 20009
rect 14372 20000 14424 20052
rect 4712 19728 4764 19780
rect 5080 19728 5132 19780
rect 6828 19864 6880 19916
rect 8944 19864 8996 19916
rect 9312 19864 9364 19916
rect 8760 19796 8812 19848
rect 9036 19796 9088 19848
rect 3148 19703 3200 19712
rect 3148 19669 3157 19703
rect 3157 19669 3191 19703
rect 3191 19669 3200 19703
rect 3148 19660 3200 19669
rect 5540 19660 5592 19712
rect 8576 19660 8628 19712
rect 9404 19660 9456 19712
rect 10968 19796 11020 19848
rect 13820 19932 13872 19984
rect 13912 19932 13964 19984
rect 14556 19932 14608 19984
rect 15016 20000 15068 20052
rect 16396 20043 16448 20052
rect 16396 20009 16405 20043
rect 16405 20009 16439 20043
rect 16439 20009 16448 20043
rect 16396 20000 16448 20009
rect 19064 20000 19116 20052
rect 19248 20000 19300 20052
rect 21456 20000 21508 20052
rect 16488 19932 16540 19984
rect 17960 19932 18012 19984
rect 13176 19864 13228 19916
rect 14832 19907 14884 19916
rect 12808 19839 12860 19848
rect 12808 19805 12817 19839
rect 12817 19805 12851 19839
rect 12851 19805 12860 19839
rect 12808 19796 12860 19805
rect 13084 19796 13136 19848
rect 14832 19873 14841 19907
rect 14841 19873 14875 19907
rect 14875 19873 14884 19907
rect 14832 19864 14884 19873
rect 13912 19796 13964 19848
rect 14740 19796 14792 19848
rect 12900 19728 12952 19780
rect 13452 19728 13504 19780
rect 16212 19864 16264 19916
rect 16580 19864 16632 19916
rect 16856 19907 16908 19916
rect 16856 19873 16865 19907
rect 16865 19873 16899 19907
rect 16899 19873 16908 19907
rect 16856 19864 16908 19873
rect 17408 19864 17460 19916
rect 20076 19932 20128 19984
rect 19984 19907 20036 19916
rect 19984 19873 19993 19907
rect 19993 19873 20027 19907
rect 20027 19873 20036 19907
rect 19984 19864 20036 19873
rect 20628 19864 20680 19916
rect 18972 19839 19024 19848
rect 18972 19805 18981 19839
rect 18981 19805 19015 19839
rect 19015 19805 19024 19839
rect 18972 19796 19024 19805
rect 15568 19728 15620 19780
rect 20076 19796 20128 19848
rect 20720 19728 20772 19780
rect 21088 19864 21140 19916
rect 22376 19864 22428 19916
rect 23204 19864 23256 19916
rect 20996 19839 21048 19848
rect 20996 19805 21005 19839
rect 21005 19805 21039 19839
rect 21039 19805 21048 19839
rect 20996 19796 21048 19805
rect 23112 19771 23164 19780
rect 23112 19737 23121 19771
rect 23121 19737 23155 19771
rect 23155 19737 23164 19771
rect 23112 19728 23164 19737
rect 10600 19660 10652 19712
rect 11060 19703 11112 19712
rect 11060 19669 11069 19703
rect 11069 19669 11103 19703
rect 11103 19669 11112 19703
rect 11060 19660 11112 19669
rect 11152 19660 11204 19712
rect 14464 19660 14516 19712
rect 14924 19660 14976 19712
rect 15200 19703 15252 19712
rect 15200 19669 15209 19703
rect 15209 19669 15243 19703
rect 15243 19669 15252 19703
rect 15200 19660 15252 19669
rect 17040 19703 17092 19712
rect 17040 19669 17049 19703
rect 17049 19669 17083 19703
rect 17083 19669 17092 19703
rect 17040 19660 17092 19669
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 17592 19660 17644 19669
rect 20168 19660 20220 19712
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 22560 19660 22612 19712
rect 4714 19558 4766 19610
rect 4778 19558 4830 19610
rect 4842 19558 4894 19610
rect 4906 19558 4958 19610
rect 12178 19558 12230 19610
rect 12242 19558 12294 19610
rect 12306 19558 12358 19610
rect 12370 19558 12422 19610
rect 19642 19558 19694 19610
rect 19706 19558 19758 19610
rect 19770 19558 19822 19610
rect 19834 19558 19886 19610
rect 3516 19456 3568 19508
rect 5908 19456 5960 19508
rect 3148 19388 3200 19440
rect 4344 19388 4396 19440
rect 9128 19456 9180 19508
rect 11520 19499 11572 19508
rect 11520 19465 11529 19499
rect 11529 19465 11563 19499
rect 11563 19465 11572 19499
rect 11520 19456 11572 19465
rect 13084 19499 13136 19508
rect 13084 19465 13093 19499
rect 13093 19465 13127 19499
rect 13127 19465 13136 19499
rect 13084 19456 13136 19465
rect 20076 19456 20128 19508
rect 22284 19456 22336 19508
rect 11152 19388 11204 19440
rect 4436 19320 4488 19372
rect 4528 19320 4580 19372
rect 5448 19363 5500 19372
rect 5448 19329 5457 19363
rect 5457 19329 5491 19363
rect 5491 19329 5500 19363
rect 5448 19320 5500 19329
rect 6460 19320 6512 19372
rect 6920 19320 6972 19372
rect 5632 19295 5684 19304
rect 5632 19261 5641 19295
rect 5641 19261 5675 19295
rect 5675 19261 5684 19295
rect 5632 19252 5684 19261
rect 5724 19252 5776 19304
rect 6644 19252 6696 19304
rect 7380 19252 7432 19304
rect 1952 19227 2004 19236
rect 1952 19193 1986 19227
rect 1986 19193 2004 19227
rect 1952 19184 2004 19193
rect 2136 19184 2188 19236
rect 2228 19184 2280 19236
rect 3056 19159 3108 19168
rect 3056 19125 3065 19159
rect 3065 19125 3099 19159
rect 3099 19125 3108 19159
rect 3056 19116 3108 19125
rect 3332 19116 3384 19168
rect 5816 19184 5868 19236
rect 8116 19320 8168 19372
rect 8576 19320 8628 19372
rect 7748 19252 7800 19304
rect 9864 19320 9916 19372
rect 10232 19363 10284 19372
rect 10232 19329 10241 19363
rect 10241 19329 10275 19363
rect 10275 19329 10284 19363
rect 10232 19320 10284 19329
rect 10416 19320 10468 19372
rect 10692 19320 10744 19372
rect 11336 19295 11388 19304
rect 11336 19261 11345 19295
rect 11345 19261 11379 19295
rect 11379 19261 11388 19295
rect 11336 19252 11388 19261
rect 12900 19320 12952 19372
rect 13728 19320 13780 19372
rect 14004 19320 14056 19372
rect 11796 19252 11848 19304
rect 4344 19159 4396 19168
rect 4344 19125 4353 19159
rect 4353 19125 4387 19159
rect 4387 19125 4396 19159
rect 4344 19116 4396 19125
rect 4804 19159 4856 19168
rect 4804 19125 4813 19159
rect 4813 19125 4847 19159
rect 4847 19125 4856 19159
rect 4804 19116 4856 19125
rect 5264 19159 5316 19168
rect 5264 19125 5273 19159
rect 5273 19125 5307 19159
rect 5307 19125 5316 19159
rect 9588 19184 9640 19236
rect 11152 19184 11204 19236
rect 13268 19184 13320 19236
rect 5264 19116 5316 19125
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 7472 19116 7524 19168
rect 9312 19116 9364 19168
rect 9680 19159 9732 19168
rect 9680 19125 9689 19159
rect 9689 19125 9723 19159
rect 9723 19125 9732 19159
rect 9680 19116 9732 19125
rect 10140 19159 10192 19168
rect 10140 19125 10149 19159
rect 10149 19125 10183 19159
rect 10183 19125 10192 19159
rect 10140 19116 10192 19125
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 10876 19159 10928 19168
rect 10876 19125 10885 19159
rect 10885 19125 10919 19159
rect 10919 19125 10928 19159
rect 11244 19159 11296 19168
rect 10876 19116 10928 19125
rect 11244 19125 11253 19159
rect 11253 19125 11287 19159
rect 11287 19125 11296 19159
rect 11244 19116 11296 19125
rect 12164 19116 12216 19168
rect 13912 19159 13964 19168
rect 13912 19125 13921 19159
rect 13921 19125 13955 19159
rect 13955 19125 13964 19159
rect 13912 19116 13964 19125
rect 14648 19116 14700 19168
rect 15200 19159 15252 19168
rect 15200 19125 15209 19159
rect 15209 19125 15243 19159
rect 15243 19125 15252 19159
rect 15200 19116 15252 19125
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 17592 19252 17644 19304
rect 18972 19252 19024 19304
rect 19156 19252 19208 19304
rect 20536 19252 20588 19304
rect 21640 19320 21692 19372
rect 22836 19363 22888 19372
rect 22836 19329 22845 19363
rect 22845 19329 22879 19363
rect 22879 19329 22888 19363
rect 22836 19320 22888 19329
rect 23572 19363 23624 19372
rect 23572 19329 23581 19363
rect 23581 19329 23615 19363
rect 23615 19329 23624 19363
rect 23572 19320 23624 19329
rect 21732 19252 21784 19304
rect 21916 19252 21968 19304
rect 22376 19252 22428 19304
rect 20352 19184 20404 19236
rect 21180 19184 21232 19236
rect 15292 19116 15344 19125
rect 15752 19116 15804 19168
rect 16580 19116 16632 19168
rect 16764 19159 16816 19168
rect 16764 19125 16773 19159
rect 16773 19125 16807 19159
rect 16807 19125 16816 19159
rect 16764 19116 16816 19125
rect 16948 19159 17000 19168
rect 16948 19125 16957 19159
rect 16957 19125 16991 19159
rect 16991 19125 17000 19159
rect 16948 19116 17000 19125
rect 19340 19159 19392 19168
rect 19340 19125 19349 19159
rect 19349 19125 19383 19159
rect 19383 19125 19392 19159
rect 19340 19116 19392 19125
rect 19432 19159 19484 19168
rect 19432 19125 19441 19159
rect 19441 19125 19475 19159
rect 19475 19125 19484 19159
rect 19432 19116 19484 19125
rect 21364 19116 21416 19168
rect 21916 19116 21968 19168
rect 23020 19159 23072 19168
rect 23020 19125 23029 19159
rect 23029 19125 23063 19159
rect 23063 19125 23072 19159
rect 23020 19116 23072 19125
rect 8446 19014 8498 19066
rect 8510 19014 8562 19066
rect 8574 19014 8626 19066
rect 8638 19014 8690 19066
rect 15910 19014 15962 19066
rect 15974 19014 16026 19066
rect 16038 19014 16090 19066
rect 16102 19014 16154 19066
rect 1952 18912 2004 18964
rect 4344 18912 4396 18964
rect 5080 18912 5132 18964
rect 5264 18955 5316 18964
rect 5264 18921 5273 18955
rect 5273 18921 5307 18955
rect 5307 18921 5316 18955
rect 5264 18912 5316 18921
rect 8116 18912 8168 18964
rect 9772 18912 9824 18964
rect 10784 18912 10836 18964
rect 11152 18912 11204 18964
rect 13268 18955 13320 18964
rect 13268 18921 13277 18955
rect 13277 18921 13311 18955
rect 13311 18921 13320 18955
rect 13268 18912 13320 18921
rect 14556 18955 14608 18964
rect 2136 18844 2188 18896
rect 2320 18776 2372 18828
rect 3056 18844 3108 18896
rect 6184 18844 6236 18896
rect 7840 18887 7892 18896
rect 7840 18853 7858 18887
rect 7858 18853 7892 18887
rect 7840 18844 7892 18853
rect 9128 18844 9180 18896
rect 11704 18844 11756 18896
rect 3608 18776 3660 18828
rect 4804 18819 4856 18828
rect 4804 18785 4813 18819
rect 4813 18785 4847 18819
rect 4847 18785 4856 18819
rect 4804 18776 4856 18785
rect 6368 18776 6420 18828
rect 7380 18776 7432 18828
rect 4436 18708 4488 18760
rect 5080 18708 5132 18760
rect 6828 18708 6880 18760
rect 8300 18751 8352 18760
rect 8300 18717 8309 18751
rect 8309 18717 8343 18751
rect 8343 18717 8352 18751
rect 8300 18708 8352 18717
rect 9036 18708 9088 18760
rect 9312 18708 9364 18760
rect 9680 18708 9732 18760
rect 10140 18776 10192 18828
rect 11060 18776 11112 18828
rect 12164 18819 12216 18828
rect 10324 18708 10376 18760
rect 12164 18785 12198 18819
rect 12198 18785 12216 18819
rect 12164 18776 12216 18785
rect 11796 18708 11848 18760
rect 14004 18844 14056 18896
rect 13912 18776 13964 18828
rect 14556 18921 14565 18955
rect 14565 18921 14599 18955
rect 14599 18921 14608 18955
rect 14556 18912 14608 18921
rect 14832 18955 14884 18964
rect 14832 18921 14841 18955
rect 14841 18921 14875 18955
rect 14875 18921 14884 18955
rect 14832 18912 14884 18921
rect 16764 18912 16816 18964
rect 15384 18844 15436 18896
rect 14648 18819 14700 18828
rect 14648 18785 14657 18819
rect 14657 18785 14691 18819
rect 14691 18785 14700 18819
rect 14648 18776 14700 18785
rect 14740 18776 14792 18828
rect 15200 18819 15252 18828
rect 15200 18785 15223 18819
rect 15223 18785 15252 18819
rect 18236 18844 18288 18896
rect 20076 18912 20128 18964
rect 20444 18912 20496 18964
rect 22376 18912 22428 18964
rect 21364 18887 21416 18896
rect 21364 18853 21398 18887
rect 21398 18853 21416 18887
rect 21364 18844 21416 18853
rect 21732 18844 21784 18896
rect 23020 18844 23072 18896
rect 15200 18776 15252 18785
rect 17408 18819 17460 18828
rect 17408 18785 17417 18819
rect 17417 18785 17451 18819
rect 17451 18785 17460 18819
rect 17408 18776 17460 18785
rect 20444 18776 20496 18828
rect 14924 18751 14976 18760
rect 8760 18640 8812 18692
rect 10968 18683 11020 18692
rect 10968 18649 10977 18683
rect 10977 18649 11011 18683
rect 11011 18649 11020 18683
rect 10968 18640 11020 18649
rect 1584 18572 1636 18624
rect 4528 18572 4580 18624
rect 6092 18572 6144 18624
rect 7932 18572 7984 18624
rect 8300 18572 8352 18624
rect 8392 18572 8444 18624
rect 9496 18572 9548 18624
rect 14924 18717 14933 18751
rect 14933 18717 14967 18751
rect 14967 18717 14976 18751
rect 14924 18708 14976 18717
rect 16212 18708 16264 18760
rect 17132 18751 17184 18760
rect 17132 18717 17144 18751
rect 17144 18717 17178 18751
rect 17178 18717 17184 18751
rect 17132 18708 17184 18717
rect 13820 18640 13872 18692
rect 13084 18572 13136 18624
rect 14372 18572 14424 18624
rect 16580 18640 16632 18692
rect 16120 18572 16172 18624
rect 16948 18572 17000 18624
rect 19156 18708 19208 18760
rect 20996 18708 21048 18760
rect 19248 18683 19300 18692
rect 19248 18649 19257 18683
rect 19257 18649 19291 18683
rect 19291 18649 19300 18683
rect 19248 18640 19300 18649
rect 18328 18572 18380 18624
rect 20352 18572 20404 18624
rect 4714 18470 4766 18522
rect 4778 18470 4830 18522
rect 4842 18470 4894 18522
rect 4906 18470 4958 18522
rect 12178 18470 12230 18522
rect 12242 18470 12294 18522
rect 12306 18470 12358 18522
rect 12370 18470 12422 18522
rect 19642 18470 19694 18522
rect 19706 18470 19758 18522
rect 19770 18470 19822 18522
rect 19834 18470 19886 18522
rect 2228 18411 2280 18420
rect 2228 18377 2237 18411
rect 2237 18377 2271 18411
rect 2271 18377 2280 18411
rect 2228 18368 2280 18377
rect 3608 18368 3660 18420
rect 1584 18275 1636 18284
rect 1584 18241 1593 18275
rect 1593 18241 1627 18275
rect 1627 18241 1636 18275
rect 1584 18232 1636 18241
rect 3056 18164 3108 18216
rect 3332 18207 3384 18216
rect 3332 18173 3350 18207
rect 3350 18173 3384 18207
rect 3332 18164 3384 18173
rect 4436 18232 4488 18284
rect 5172 18368 5224 18420
rect 7656 18368 7708 18420
rect 10048 18368 10100 18420
rect 13912 18411 13964 18420
rect 9036 18300 9088 18352
rect 4620 18232 4672 18284
rect 3608 18207 3660 18216
rect 3608 18173 3610 18207
rect 3610 18173 3644 18207
rect 3644 18173 3660 18207
rect 3608 18164 3660 18173
rect 3792 18164 3844 18216
rect 8392 18232 8444 18284
rect 8760 18232 8812 18284
rect 10876 18232 10928 18284
rect 11244 18232 11296 18284
rect 5080 18207 5132 18216
rect 5080 18173 5114 18207
rect 5114 18173 5132 18207
rect 5080 18164 5132 18173
rect 9036 18207 9088 18216
rect 9036 18173 9045 18207
rect 9045 18173 9079 18207
rect 9079 18173 9088 18207
rect 9036 18164 9088 18173
rect 9220 18164 9272 18216
rect 9680 18164 9732 18216
rect 6092 18096 6144 18148
rect 12072 18300 12124 18352
rect 13912 18377 13921 18411
rect 13921 18377 13955 18411
rect 13955 18377 13964 18411
rect 13912 18368 13964 18377
rect 14740 18411 14792 18420
rect 14740 18377 14749 18411
rect 14749 18377 14783 18411
rect 14783 18377 14792 18411
rect 14740 18368 14792 18377
rect 16672 18368 16724 18420
rect 18236 18411 18288 18420
rect 18236 18377 18245 18411
rect 18245 18377 18279 18411
rect 18279 18377 18288 18411
rect 18236 18368 18288 18377
rect 22468 18368 22520 18420
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 13728 18232 13780 18284
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 16304 18232 16356 18284
rect 16856 18300 16908 18352
rect 17592 18275 17644 18284
rect 17592 18241 17601 18275
rect 17601 18241 17635 18275
rect 17635 18241 17644 18275
rect 17592 18232 17644 18241
rect 17684 18232 17736 18284
rect 22836 18275 22888 18284
rect 15292 18164 15344 18216
rect 15476 18096 15528 18148
rect 15568 18096 15620 18148
rect 17132 18164 17184 18216
rect 17960 18164 18012 18216
rect 22836 18241 22845 18275
rect 22845 18241 22879 18275
rect 22879 18241 22888 18275
rect 22836 18232 22888 18241
rect 19432 18164 19484 18216
rect 19708 18164 19760 18216
rect 20168 18207 20220 18216
rect 20168 18173 20177 18207
rect 20177 18173 20211 18207
rect 20211 18173 20220 18207
rect 20168 18164 20220 18173
rect 19156 18096 19208 18148
rect 22652 18164 22704 18216
rect 20996 18096 21048 18148
rect 21364 18096 21416 18148
rect 4068 18071 4120 18080
rect 4068 18037 4077 18071
rect 4077 18037 4111 18071
rect 4111 18037 4120 18071
rect 4068 18028 4120 18037
rect 6184 18071 6236 18080
rect 6184 18037 6193 18071
rect 6193 18037 6227 18071
rect 6227 18037 6236 18071
rect 6184 18028 6236 18037
rect 6920 18071 6972 18080
rect 6920 18037 6929 18071
rect 6929 18037 6963 18071
rect 6963 18037 6972 18071
rect 6920 18028 6972 18037
rect 9312 18028 9364 18080
rect 12716 18028 12768 18080
rect 14280 18071 14332 18080
rect 14280 18037 14289 18071
rect 14289 18037 14323 18071
rect 14323 18037 14332 18071
rect 14280 18028 14332 18037
rect 14832 18028 14884 18080
rect 17224 18071 17276 18080
rect 17224 18037 17233 18071
rect 17233 18037 17267 18071
rect 17267 18037 17276 18071
rect 17224 18028 17276 18037
rect 17408 18071 17460 18080
rect 17408 18037 17417 18071
rect 17417 18037 17451 18071
rect 17451 18037 17460 18071
rect 17408 18028 17460 18037
rect 18236 18028 18288 18080
rect 20444 18028 20496 18080
rect 22008 18071 22060 18080
rect 22008 18037 22017 18071
rect 22017 18037 22051 18071
rect 22051 18037 22060 18071
rect 22008 18028 22060 18037
rect 22560 18028 22612 18080
rect 8446 17926 8498 17978
rect 8510 17926 8562 17978
rect 8574 17926 8626 17978
rect 8638 17926 8690 17978
rect 15910 17926 15962 17978
rect 15974 17926 16026 17978
rect 16038 17926 16090 17978
rect 16102 17926 16154 17978
rect 3056 17824 3108 17876
rect 5080 17824 5132 17876
rect 3424 17756 3476 17808
rect 3792 17756 3844 17808
rect 1768 17688 1820 17740
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 3240 17620 3292 17672
rect 4436 17620 4488 17672
rect 6828 17824 6880 17876
rect 7196 17824 7248 17876
rect 11244 17824 11296 17876
rect 13820 17824 13872 17876
rect 15292 17824 15344 17876
rect 18696 17824 18748 17876
rect 19708 17824 19760 17876
rect 20720 17824 20772 17876
rect 6092 17688 6144 17740
rect 7288 17688 7340 17740
rect 7932 17756 7984 17808
rect 8300 17663 8352 17672
rect 8300 17629 8309 17663
rect 8309 17629 8343 17663
rect 8343 17629 8352 17663
rect 8300 17620 8352 17629
rect 11060 17756 11112 17808
rect 14280 17756 14332 17808
rect 14924 17756 14976 17808
rect 16580 17756 16632 17808
rect 17224 17756 17276 17808
rect 4068 17552 4120 17604
rect 7196 17552 7248 17604
rect 6368 17484 6420 17536
rect 7012 17484 7064 17536
rect 9404 17620 9456 17672
rect 12072 17688 12124 17740
rect 13360 17688 13412 17740
rect 14372 17731 14424 17740
rect 14372 17697 14381 17731
rect 14381 17697 14415 17731
rect 14415 17697 14424 17731
rect 14372 17688 14424 17697
rect 16396 17688 16448 17740
rect 11520 17620 11572 17672
rect 12900 17663 12952 17672
rect 10416 17552 10468 17604
rect 12900 17629 12909 17663
rect 12909 17629 12943 17663
rect 12943 17629 12952 17663
rect 12900 17620 12952 17629
rect 13084 17663 13136 17672
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 17408 17688 17460 17740
rect 19524 17756 19576 17808
rect 22560 17756 22612 17808
rect 19064 17688 19116 17740
rect 17684 17620 17736 17672
rect 19340 17620 19392 17672
rect 21088 17731 21140 17740
rect 21088 17697 21097 17731
rect 21097 17697 21131 17731
rect 21131 17697 21140 17731
rect 21088 17688 21140 17697
rect 20996 17663 21048 17672
rect 9312 17484 9364 17536
rect 13544 17484 13596 17536
rect 15476 17552 15528 17604
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 21456 17688 21508 17740
rect 22100 17688 22152 17740
rect 20996 17620 21048 17629
rect 17500 17484 17552 17536
rect 17592 17484 17644 17536
rect 22652 17552 22704 17604
rect 19340 17484 19392 17536
rect 22560 17484 22612 17536
rect 4714 17382 4766 17434
rect 4778 17382 4830 17434
rect 4842 17382 4894 17434
rect 4906 17382 4958 17434
rect 12178 17382 12230 17434
rect 12242 17382 12294 17434
rect 12306 17382 12358 17434
rect 12370 17382 12422 17434
rect 19642 17382 19694 17434
rect 19706 17382 19758 17434
rect 19770 17382 19822 17434
rect 19834 17382 19886 17434
rect 1768 17323 1820 17332
rect 1768 17289 1777 17323
rect 1777 17289 1811 17323
rect 1811 17289 1820 17323
rect 1768 17280 1820 17289
rect 3332 17280 3384 17332
rect 5816 17280 5868 17332
rect 9588 17280 9640 17332
rect 13360 17323 13412 17332
rect 13360 17289 13369 17323
rect 13369 17289 13403 17323
rect 13403 17289 13412 17323
rect 13360 17280 13412 17289
rect 14924 17323 14976 17332
rect 14924 17289 14933 17323
rect 14933 17289 14967 17323
rect 14967 17289 14976 17323
rect 14924 17280 14976 17289
rect 17684 17280 17736 17332
rect 19064 17323 19116 17332
rect 19064 17289 19073 17323
rect 19073 17289 19107 17323
rect 19107 17289 19116 17323
rect 19064 17280 19116 17289
rect 19984 17323 20036 17332
rect 19984 17289 19993 17323
rect 19993 17289 20027 17323
rect 20027 17289 20036 17323
rect 19984 17280 20036 17289
rect 21088 17280 21140 17332
rect 4620 17212 4672 17264
rect 3240 17144 3292 17196
rect 9680 17212 9732 17264
rect 6828 17144 6880 17196
rect 7472 17144 7524 17196
rect 4068 17076 4120 17128
rect 6184 17076 6236 17128
rect 7288 17076 7340 17128
rect 8208 17076 8260 17128
rect 11796 17144 11848 17196
rect 14832 17255 14884 17264
rect 14832 17221 14841 17255
rect 14841 17221 14875 17255
rect 14875 17221 14884 17255
rect 14832 17212 14884 17221
rect 16488 17212 16540 17264
rect 10324 17076 10376 17128
rect 4068 16940 4120 16992
rect 6184 16983 6236 16992
rect 6184 16949 6193 16983
rect 6193 16949 6227 16983
rect 6227 16949 6236 16983
rect 6184 16940 6236 16949
rect 6828 16983 6880 16992
rect 6828 16949 6837 16983
rect 6837 16949 6871 16983
rect 6871 16949 6880 16983
rect 6828 16940 6880 16949
rect 7840 16983 7892 16992
rect 7840 16949 7849 16983
rect 7849 16949 7883 16983
rect 7883 16949 7892 16983
rect 7840 16940 7892 16949
rect 8300 16940 8352 16992
rect 8668 17008 8720 17060
rect 11336 17076 11388 17128
rect 11980 17119 12032 17128
rect 11980 17085 11989 17119
rect 11989 17085 12023 17119
rect 12023 17085 12032 17119
rect 11980 17076 12032 17085
rect 13084 17076 13136 17128
rect 16304 17187 16356 17196
rect 16304 17153 16313 17187
rect 16313 17153 16347 17187
rect 16347 17153 16356 17187
rect 16304 17144 16356 17153
rect 8852 16940 8904 16992
rect 9864 16940 9916 16992
rect 10508 16983 10560 16992
rect 10508 16949 10517 16983
rect 10517 16949 10551 16983
rect 10551 16949 10560 16983
rect 10508 16940 10560 16949
rect 11152 16940 11204 16992
rect 11520 17008 11572 17060
rect 16856 17076 16908 17128
rect 17592 17119 17644 17128
rect 17592 17085 17601 17119
rect 17601 17085 17635 17119
rect 17635 17085 17644 17119
rect 17592 17076 17644 17085
rect 17684 17119 17736 17128
rect 17684 17085 17700 17119
rect 17700 17085 17734 17119
rect 17734 17085 17736 17119
rect 19340 17212 19392 17264
rect 22192 17280 22244 17332
rect 22100 17212 22152 17264
rect 19616 17144 19668 17196
rect 20444 17187 20496 17196
rect 17684 17076 17736 17085
rect 15200 16940 15252 16992
rect 16212 16940 16264 16992
rect 17132 16983 17184 16992
rect 17132 16949 17141 16983
rect 17141 16949 17175 16983
rect 17175 16949 17184 16983
rect 17132 16940 17184 16949
rect 17776 17008 17828 17060
rect 20444 17153 20453 17187
rect 20453 17153 20487 17187
rect 20487 17153 20496 17187
rect 20444 17144 20496 17153
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 20720 17144 20772 17196
rect 22468 17144 22520 17196
rect 22744 17187 22796 17196
rect 22744 17153 22753 17187
rect 22753 17153 22787 17187
rect 22787 17153 22796 17187
rect 22744 17144 22796 17153
rect 20352 17119 20404 17128
rect 20352 17085 20361 17119
rect 20361 17085 20395 17119
rect 20395 17085 20404 17119
rect 20352 17076 20404 17085
rect 20444 17008 20496 17060
rect 21364 17119 21416 17128
rect 21364 17085 21373 17119
rect 21373 17085 21407 17119
rect 21407 17085 21416 17119
rect 21364 17076 21416 17085
rect 21824 17119 21876 17128
rect 21824 17085 21833 17119
rect 21833 17085 21867 17119
rect 21867 17085 21876 17119
rect 21824 17076 21876 17085
rect 22560 17119 22612 17128
rect 22560 17085 22569 17119
rect 22569 17085 22603 17119
rect 22603 17085 22612 17119
rect 22560 17076 22612 17085
rect 21916 17008 21968 17060
rect 19248 16940 19300 16992
rect 19892 16983 19944 16992
rect 19892 16949 19901 16983
rect 19901 16949 19935 16983
rect 19935 16949 19944 16983
rect 19892 16940 19944 16949
rect 22192 16983 22244 16992
rect 22192 16949 22201 16983
rect 22201 16949 22235 16983
rect 22235 16949 22244 16983
rect 22192 16940 22244 16949
rect 8446 16838 8498 16890
rect 8510 16838 8562 16890
rect 8574 16838 8626 16890
rect 8638 16838 8690 16890
rect 15910 16838 15962 16890
rect 15974 16838 16026 16890
rect 16038 16838 16090 16890
rect 16102 16838 16154 16890
rect 3240 16736 3292 16788
rect 2780 16668 2832 16720
rect 6828 16736 6880 16788
rect 6920 16736 6972 16788
rect 7472 16779 7524 16788
rect 7472 16745 7481 16779
rect 7481 16745 7515 16779
rect 7515 16745 7524 16779
rect 7472 16736 7524 16745
rect 7840 16736 7892 16788
rect 6184 16668 6236 16720
rect 6552 16668 6604 16720
rect 4620 16600 4672 16652
rect 6368 16600 6420 16652
rect 7012 16600 7064 16652
rect 8484 16668 8536 16720
rect 8944 16668 8996 16720
rect 13084 16736 13136 16788
rect 14464 16736 14516 16788
rect 16212 16736 16264 16788
rect 17776 16736 17828 16788
rect 9772 16668 9824 16720
rect 6184 16575 6236 16584
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 7196 16532 7248 16584
rect 8024 16600 8076 16652
rect 11796 16668 11848 16720
rect 13636 16711 13688 16720
rect 13636 16677 13645 16711
rect 13645 16677 13679 16711
rect 13679 16677 13688 16711
rect 13636 16668 13688 16677
rect 14556 16711 14608 16720
rect 14556 16677 14565 16711
rect 14565 16677 14599 16711
rect 14599 16677 14608 16711
rect 14556 16668 14608 16677
rect 16948 16668 17000 16720
rect 17500 16668 17552 16720
rect 19800 16736 19852 16788
rect 19892 16736 19944 16788
rect 18052 16668 18104 16720
rect 19432 16668 19484 16720
rect 22008 16668 22060 16720
rect 11704 16600 11756 16652
rect 13176 16643 13228 16652
rect 13176 16609 13185 16643
rect 13185 16609 13219 16643
rect 13219 16609 13228 16643
rect 13176 16600 13228 16609
rect 15476 16643 15528 16652
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 15660 16600 15712 16652
rect 16304 16600 16356 16652
rect 18880 16600 18932 16652
rect 19064 16643 19116 16652
rect 19064 16609 19073 16643
rect 19073 16609 19107 16643
rect 19107 16609 19116 16643
rect 19064 16600 19116 16609
rect 19984 16643 20036 16652
rect 8852 16575 8904 16584
rect 8852 16541 8861 16575
rect 8861 16541 8895 16575
rect 8895 16541 8904 16575
rect 8852 16532 8904 16541
rect 4068 16396 4120 16448
rect 4528 16439 4580 16448
rect 4528 16405 4537 16439
rect 4537 16405 4571 16439
rect 4571 16405 4580 16439
rect 4528 16396 4580 16405
rect 5448 16396 5500 16448
rect 8116 16396 8168 16448
rect 11152 16575 11204 16584
rect 10784 16396 10836 16448
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 12900 16575 12952 16584
rect 12900 16541 12909 16575
rect 12909 16541 12943 16575
rect 12943 16541 12952 16575
rect 12900 16532 12952 16541
rect 14464 16575 14516 16584
rect 14464 16541 14473 16575
rect 14473 16541 14507 16575
rect 14507 16541 14516 16575
rect 14464 16532 14516 16541
rect 14648 16575 14700 16584
rect 14648 16541 14657 16575
rect 14657 16541 14691 16575
rect 14691 16541 14700 16575
rect 14648 16532 14700 16541
rect 18972 16575 19024 16584
rect 18972 16541 18981 16575
rect 18981 16541 19015 16575
rect 19015 16541 19024 16575
rect 18972 16532 19024 16541
rect 16304 16396 16356 16448
rect 17408 16396 17460 16448
rect 19432 16532 19484 16584
rect 19340 16464 19392 16516
rect 19984 16609 19993 16643
rect 19993 16609 20027 16643
rect 20027 16609 20036 16643
rect 19984 16600 20036 16609
rect 20536 16600 20588 16652
rect 21456 16643 21508 16652
rect 21456 16609 21465 16643
rect 21465 16609 21499 16643
rect 21499 16609 21508 16643
rect 21456 16600 21508 16609
rect 23112 16643 23164 16652
rect 23112 16609 23121 16643
rect 23121 16609 23155 16643
rect 23155 16609 23164 16643
rect 23112 16600 23164 16609
rect 20720 16532 20772 16584
rect 20904 16575 20956 16584
rect 20904 16541 20913 16575
rect 20913 16541 20947 16575
rect 20947 16541 20956 16575
rect 20904 16532 20956 16541
rect 21456 16396 21508 16448
rect 22836 16439 22888 16448
rect 22836 16405 22845 16439
rect 22845 16405 22879 16439
rect 22879 16405 22888 16439
rect 22836 16396 22888 16405
rect 22928 16439 22980 16448
rect 22928 16405 22937 16439
rect 22937 16405 22971 16439
rect 22971 16405 22980 16439
rect 22928 16396 22980 16405
rect 4714 16294 4766 16346
rect 4778 16294 4830 16346
rect 4842 16294 4894 16346
rect 4906 16294 4958 16346
rect 12178 16294 12230 16346
rect 12242 16294 12294 16346
rect 12306 16294 12358 16346
rect 12370 16294 12422 16346
rect 19642 16294 19694 16346
rect 19706 16294 19758 16346
rect 19770 16294 19822 16346
rect 19834 16294 19886 16346
rect 3424 16235 3476 16244
rect 3424 16201 3433 16235
rect 3433 16201 3467 16235
rect 3467 16201 3476 16235
rect 3424 16192 3476 16201
rect 7564 16192 7616 16244
rect 8300 16192 8352 16244
rect 4620 16124 4672 16176
rect 5448 16056 5500 16108
rect 6000 16056 6052 16108
rect 2780 15988 2832 16040
rect 4528 15988 4580 16040
rect 6920 16124 6972 16176
rect 8944 16099 8996 16108
rect 1584 15963 1636 15972
rect 1584 15929 1593 15963
rect 1593 15929 1627 15963
rect 1627 15929 1636 15963
rect 1584 15920 1636 15929
rect 1768 15920 1820 15972
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 4160 15895 4212 15904
rect 4160 15861 4169 15895
rect 4169 15861 4203 15895
rect 4203 15861 4212 15895
rect 4160 15852 4212 15861
rect 6736 15988 6788 16040
rect 8024 15988 8076 16040
rect 6368 15920 6420 15972
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5816 15895 5868 15904
rect 5172 15852 5224 15861
rect 5816 15861 5825 15895
rect 5825 15861 5859 15895
rect 5859 15861 5868 15895
rect 5816 15852 5868 15861
rect 5908 15895 5960 15904
rect 5908 15861 5917 15895
rect 5917 15861 5951 15895
rect 5951 15861 5960 15895
rect 7012 15920 7064 15972
rect 8208 15920 8260 15972
rect 8944 16065 8953 16099
rect 8953 16065 8987 16099
rect 8987 16065 8996 16099
rect 8944 16056 8996 16065
rect 9128 16056 9180 16108
rect 14556 16192 14608 16244
rect 17316 16192 17368 16244
rect 18880 16192 18932 16244
rect 12164 16124 12216 16176
rect 14280 16124 14332 16176
rect 9864 16099 9916 16108
rect 9864 16065 9876 16099
rect 9876 16065 9910 16099
rect 9910 16065 9916 16099
rect 9864 16056 9916 16065
rect 10324 16056 10376 16108
rect 11980 15988 12032 16040
rect 12900 15988 12952 16040
rect 5908 15852 5960 15861
rect 8760 15895 8812 15904
rect 8760 15861 8769 15895
rect 8769 15861 8803 15895
rect 8803 15861 8812 15895
rect 8760 15852 8812 15861
rect 8852 15895 8904 15904
rect 8852 15861 8861 15895
rect 8861 15861 8895 15895
rect 8895 15861 8904 15895
rect 9312 15895 9364 15904
rect 8852 15852 8904 15861
rect 9312 15861 9321 15895
rect 9321 15861 9355 15895
rect 9355 15861 9364 15895
rect 9312 15852 9364 15861
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 11336 15895 11388 15904
rect 11336 15861 11345 15895
rect 11345 15861 11379 15895
rect 11379 15861 11388 15895
rect 12624 15920 12676 15972
rect 13176 15920 13228 15972
rect 11336 15852 11388 15861
rect 12716 15852 12768 15904
rect 13360 15852 13412 15904
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 15752 16056 15804 16108
rect 15660 16031 15712 16040
rect 14096 15920 14148 15972
rect 15660 15997 15669 16031
rect 15669 15997 15703 16031
rect 15703 15997 15712 16031
rect 15660 15988 15712 15997
rect 17132 15988 17184 16040
rect 17500 16031 17552 16040
rect 17500 15997 17509 16031
rect 17509 15997 17543 16031
rect 17543 15997 17552 16031
rect 17500 15988 17552 15997
rect 17592 16031 17644 16040
rect 17592 15997 17601 16031
rect 17601 15997 17635 16031
rect 17635 15997 17644 16031
rect 17868 16031 17920 16040
rect 17592 15988 17644 15997
rect 17868 15997 17902 16031
rect 17902 15997 17920 16031
rect 19616 16124 19668 16176
rect 19524 16099 19576 16108
rect 19524 16065 19533 16099
rect 19533 16065 19567 16099
rect 19567 16065 19576 16099
rect 19524 16056 19576 16065
rect 19984 16192 20036 16244
rect 20904 16192 20956 16244
rect 21824 16235 21876 16244
rect 21824 16201 21833 16235
rect 21833 16201 21867 16235
rect 21867 16201 21876 16235
rect 21824 16192 21876 16201
rect 19800 16124 19852 16176
rect 23112 16192 23164 16244
rect 20076 16056 20128 16108
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 22376 16099 22428 16108
rect 17868 15988 17920 15997
rect 19340 15988 19392 16040
rect 20720 15988 20772 16040
rect 21456 16031 21508 16040
rect 21456 15997 21465 16031
rect 21465 15997 21499 16031
rect 21499 15997 21508 16031
rect 21456 15988 21508 15997
rect 13728 15852 13780 15904
rect 14188 15852 14240 15904
rect 15384 15895 15436 15904
rect 18512 15920 18564 15972
rect 15384 15861 15399 15895
rect 15399 15861 15433 15895
rect 15433 15861 15436 15895
rect 15384 15852 15436 15861
rect 17224 15852 17276 15904
rect 17592 15852 17644 15904
rect 18880 15852 18932 15904
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 22192 15988 22244 16040
rect 22744 15920 22796 15972
rect 19800 15895 19852 15904
rect 19800 15861 19809 15895
rect 19809 15861 19843 15895
rect 19843 15861 19852 15895
rect 19800 15852 19852 15861
rect 20076 15852 20128 15904
rect 8446 15750 8498 15802
rect 8510 15750 8562 15802
rect 8574 15750 8626 15802
rect 8638 15750 8690 15802
rect 15910 15750 15962 15802
rect 15974 15750 16026 15802
rect 16038 15750 16090 15802
rect 16102 15750 16154 15802
rect 2780 15648 2832 15700
rect 3516 15648 3568 15700
rect 4068 15648 4120 15700
rect 1768 15555 1820 15564
rect 1768 15521 1802 15555
rect 1802 15521 1820 15555
rect 1768 15512 1820 15521
rect 5448 15580 5500 15632
rect 8208 15691 8260 15700
rect 8208 15657 8217 15691
rect 8217 15657 8251 15691
rect 8251 15657 8260 15691
rect 8208 15648 8260 15657
rect 8760 15648 8812 15700
rect 9680 15648 9732 15700
rect 9864 15691 9916 15700
rect 9864 15657 9873 15691
rect 9873 15657 9907 15691
rect 9907 15657 9916 15691
rect 9864 15648 9916 15657
rect 10048 15648 10100 15700
rect 10508 15648 10560 15700
rect 10600 15648 10652 15700
rect 11244 15648 11296 15700
rect 3700 15512 3752 15564
rect 3976 15512 4028 15564
rect 4528 15512 4580 15564
rect 6000 15512 6052 15564
rect 6828 15580 6880 15632
rect 11336 15580 11388 15632
rect 7564 15512 7616 15564
rect 3240 15487 3292 15496
rect 3240 15453 3249 15487
rect 3249 15453 3283 15487
rect 3283 15453 3292 15487
rect 3240 15444 3292 15453
rect 6736 15444 6788 15496
rect 7932 15444 7984 15496
rect 9772 15444 9824 15496
rect 11520 15512 11572 15564
rect 12624 15648 12676 15700
rect 12716 15691 12768 15700
rect 12716 15657 12731 15691
rect 12731 15657 12765 15691
rect 12765 15657 12768 15691
rect 14096 15691 14148 15700
rect 12716 15648 12768 15657
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 15660 15648 15712 15700
rect 14188 15580 14240 15632
rect 14464 15580 14516 15632
rect 17868 15648 17920 15700
rect 18972 15691 19024 15700
rect 18972 15657 18981 15691
rect 18981 15657 19015 15691
rect 19015 15657 19024 15691
rect 18972 15648 19024 15657
rect 16120 15580 16172 15632
rect 16304 15580 16356 15632
rect 19800 15648 19852 15700
rect 22744 15691 22796 15700
rect 22744 15657 22753 15691
rect 22753 15657 22787 15691
rect 22787 15657 22796 15691
rect 22744 15648 22796 15657
rect 20260 15580 20312 15632
rect 20536 15580 20588 15632
rect 20720 15623 20772 15632
rect 20720 15589 20738 15623
rect 20738 15589 20772 15623
rect 20720 15580 20772 15589
rect 22284 15580 22336 15632
rect 22836 15580 22888 15632
rect 16396 15512 16448 15564
rect 17500 15512 17552 15564
rect 10600 15444 10652 15496
rect 10784 15487 10836 15496
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 10784 15444 10836 15453
rect 12164 15444 12216 15496
rect 12716 15487 12768 15496
rect 12716 15453 12728 15487
rect 12728 15453 12762 15487
rect 12762 15453 12768 15487
rect 12716 15444 12768 15453
rect 13728 15444 13780 15496
rect 17592 15444 17644 15496
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 19064 15512 19116 15564
rect 19340 15444 19392 15496
rect 9220 15376 9272 15428
rect 2872 15351 2924 15360
rect 2872 15317 2881 15351
rect 2881 15317 2915 15351
rect 2915 15317 2924 15351
rect 2872 15308 2924 15317
rect 3884 15308 3936 15360
rect 5264 15351 5316 15360
rect 5264 15317 5273 15351
rect 5273 15317 5307 15351
rect 5307 15317 5316 15351
rect 5264 15308 5316 15317
rect 10140 15308 10192 15360
rect 11704 15308 11756 15360
rect 11796 15308 11848 15360
rect 18880 15308 18932 15360
rect 19984 15512 20036 15564
rect 21180 15512 21232 15564
rect 20628 15308 20680 15360
rect 21456 15308 21508 15360
rect 22560 15308 22612 15360
rect 4714 15206 4766 15258
rect 4778 15206 4830 15258
rect 4842 15206 4894 15258
rect 4906 15206 4958 15258
rect 12178 15206 12230 15258
rect 12242 15206 12294 15258
rect 12306 15206 12358 15258
rect 12370 15206 12422 15258
rect 19642 15206 19694 15258
rect 19706 15206 19758 15258
rect 19770 15206 19822 15258
rect 19834 15206 19886 15258
rect 4528 15104 4580 15156
rect 3516 15011 3568 15020
rect 3516 14977 3525 15011
rect 3525 14977 3559 15011
rect 3559 14977 3568 15011
rect 3516 14968 3568 14977
rect 5172 15104 5224 15156
rect 6368 15104 6420 15156
rect 8852 15104 8904 15156
rect 9864 15104 9916 15156
rect 10048 15147 10100 15156
rect 10048 15113 10057 15147
rect 10057 15113 10091 15147
rect 10091 15113 10100 15147
rect 10048 15104 10100 15113
rect 6736 14968 6788 15020
rect 6920 14968 6972 15020
rect 8116 15036 8168 15088
rect 14464 15147 14516 15156
rect 14464 15113 14473 15147
rect 14473 15113 14507 15147
rect 14507 15113 14516 15147
rect 14464 15104 14516 15113
rect 15752 15147 15804 15156
rect 15752 15113 15761 15147
rect 15761 15113 15795 15147
rect 15795 15113 15804 15147
rect 15752 15104 15804 15113
rect 11520 15079 11572 15088
rect 7564 15011 7616 15020
rect 7564 14977 7573 15011
rect 7573 14977 7607 15011
rect 7607 14977 7616 15011
rect 7564 14968 7616 14977
rect 9220 14968 9272 15020
rect 9404 14968 9456 15020
rect 11520 15045 11529 15079
rect 11529 15045 11563 15079
rect 11563 15045 11572 15079
rect 11520 15036 11572 15045
rect 11888 15036 11940 15088
rect 3148 14900 3200 14952
rect 5264 14900 5316 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 7932 14900 7984 14952
rect 2228 14832 2280 14884
rect 4068 14832 4120 14884
rect 6000 14832 6052 14884
rect 9404 14832 9456 14884
rect 10140 15011 10192 15020
rect 10140 14977 10149 15011
rect 10149 14977 10183 15011
rect 10183 14977 10192 15011
rect 10140 14968 10192 14977
rect 11980 14968 12032 15020
rect 18144 15147 18196 15156
rect 18144 15113 18153 15147
rect 18153 15113 18187 15147
rect 18187 15113 18196 15147
rect 18144 15104 18196 15113
rect 18420 15104 18472 15156
rect 19156 15104 19208 15156
rect 20628 15104 20680 15156
rect 20812 15104 20864 15156
rect 16120 15036 16172 15088
rect 16212 15011 16264 15020
rect 16212 14977 16221 15011
rect 16221 14977 16255 15011
rect 16255 14977 16264 15011
rect 16212 14968 16264 14977
rect 16396 15036 16448 15088
rect 17776 14968 17828 15020
rect 22192 15036 22244 15088
rect 22284 15011 22336 15020
rect 11336 14900 11388 14952
rect 11888 14900 11940 14952
rect 12164 14900 12216 14952
rect 12532 14943 12584 14952
rect 12532 14909 12541 14943
rect 12541 14909 12575 14943
rect 12575 14909 12584 14943
rect 12532 14900 12584 14909
rect 13360 14943 13412 14952
rect 13360 14909 13394 14943
rect 13394 14909 13412 14943
rect 13360 14900 13412 14909
rect 15476 14943 15528 14952
rect 15476 14909 15485 14943
rect 15485 14909 15519 14943
rect 15519 14909 15528 14943
rect 17224 14943 17276 14952
rect 15476 14900 15528 14909
rect 17224 14909 17233 14943
rect 17233 14909 17267 14943
rect 17267 14909 17276 14943
rect 17224 14900 17276 14909
rect 18052 14943 18104 14952
rect 18052 14909 18061 14943
rect 18061 14909 18095 14943
rect 18095 14909 18104 14943
rect 18052 14900 18104 14909
rect 19892 14943 19944 14952
rect 12808 14832 12860 14884
rect 13820 14832 13872 14884
rect 10968 14764 11020 14816
rect 11060 14764 11112 14816
rect 11612 14764 11664 14816
rect 11796 14764 11848 14816
rect 12164 14807 12216 14816
rect 12164 14773 12173 14807
rect 12173 14773 12207 14807
rect 12207 14773 12216 14807
rect 12164 14764 12216 14773
rect 13728 14764 13780 14816
rect 14648 14832 14700 14884
rect 17500 14832 17552 14884
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 15568 14764 15620 14816
rect 16304 14764 16356 14816
rect 18420 14764 18472 14816
rect 19892 14909 19901 14943
rect 19901 14909 19935 14943
rect 19935 14909 19944 14943
rect 19892 14900 19944 14909
rect 20720 14900 20772 14952
rect 22284 14977 22293 15011
rect 22293 14977 22327 15011
rect 22327 14977 22336 15011
rect 22284 14968 22336 14977
rect 22928 14968 22980 15020
rect 22100 14900 22152 14952
rect 19248 14832 19300 14884
rect 18880 14764 18932 14816
rect 19524 14764 19576 14816
rect 19984 14832 20036 14884
rect 19892 14764 19944 14816
rect 20444 14764 20496 14816
rect 21364 14807 21416 14816
rect 21364 14773 21373 14807
rect 21373 14773 21407 14807
rect 21407 14773 21416 14807
rect 21364 14764 21416 14773
rect 22468 14764 22520 14816
rect 8446 14662 8498 14714
rect 8510 14662 8562 14714
rect 8574 14662 8626 14714
rect 8638 14662 8690 14714
rect 15910 14662 15962 14714
rect 15974 14662 16026 14714
rect 16038 14662 16090 14714
rect 16102 14662 16154 14714
rect 4160 14560 4212 14612
rect 6000 14603 6052 14612
rect 6000 14569 6009 14603
rect 6009 14569 6043 14603
rect 6043 14569 6052 14603
rect 6000 14560 6052 14569
rect 7288 14560 7340 14612
rect 2872 14535 2924 14544
rect 2872 14501 2890 14535
rect 2890 14501 2924 14535
rect 2872 14492 2924 14501
rect 5264 14492 5316 14544
rect 7196 14492 7248 14544
rect 3148 14467 3200 14476
rect 3148 14433 3157 14467
rect 3157 14433 3191 14467
rect 3191 14433 3200 14467
rect 3148 14424 3200 14433
rect 3884 14467 3936 14476
rect 3884 14433 3893 14467
rect 3893 14433 3927 14467
rect 3927 14433 3936 14467
rect 3884 14424 3936 14433
rect 6276 14424 6328 14476
rect 8760 14467 8812 14476
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 7196 14399 7248 14408
rect 7196 14365 7205 14399
rect 7205 14365 7239 14399
rect 7239 14365 7248 14399
rect 7196 14356 7248 14365
rect 8760 14433 8769 14467
rect 8769 14433 8803 14467
rect 8803 14433 8812 14467
rect 8760 14424 8812 14433
rect 8852 14356 8904 14408
rect 11244 14535 11296 14544
rect 11244 14501 11253 14535
rect 11253 14501 11287 14535
rect 11287 14501 11296 14535
rect 11244 14492 11296 14501
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 11060 14399 11112 14408
rect 11060 14365 11069 14399
rect 11069 14365 11103 14399
rect 11103 14365 11112 14399
rect 11060 14356 11112 14365
rect 11980 14492 12032 14544
rect 12256 14492 12308 14544
rect 13820 14603 13872 14612
rect 13820 14569 13829 14603
rect 13829 14569 13863 14603
rect 13863 14569 13872 14603
rect 13820 14560 13872 14569
rect 14280 14560 14332 14612
rect 15476 14560 15528 14612
rect 17592 14560 17644 14612
rect 17960 14560 18012 14612
rect 11612 14424 11664 14476
rect 11704 14356 11756 14408
rect 14556 14467 14608 14476
rect 9404 14331 9456 14340
rect 9404 14297 9413 14331
rect 9413 14297 9447 14331
rect 9447 14297 9456 14331
rect 9404 14288 9456 14297
rect 2228 14220 2280 14272
rect 3976 14220 4028 14272
rect 8484 14220 8536 14272
rect 12164 14288 12216 14340
rect 12532 14356 12584 14408
rect 14556 14433 14565 14467
rect 14565 14433 14599 14467
rect 14599 14433 14608 14467
rect 14556 14424 14608 14433
rect 13360 14356 13412 14408
rect 16580 14492 16632 14544
rect 19340 14560 19392 14612
rect 19984 14603 20036 14612
rect 19984 14569 19993 14603
rect 19993 14569 20027 14603
rect 20027 14569 20036 14603
rect 19984 14560 20036 14569
rect 20260 14560 20312 14612
rect 20720 14560 20772 14612
rect 22192 14560 22244 14612
rect 22376 14560 22428 14612
rect 22100 14492 22152 14544
rect 15752 14424 15804 14476
rect 16764 14467 16816 14476
rect 16764 14433 16798 14467
rect 16798 14433 16816 14467
rect 16764 14424 16816 14433
rect 18052 14424 18104 14476
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 16212 14356 16264 14408
rect 17868 14356 17920 14408
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 13820 14288 13872 14340
rect 19432 14424 19484 14476
rect 19984 14424 20036 14476
rect 19800 14399 19852 14408
rect 19800 14365 19809 14399
rect 19809 14365 19843 14399
rect 19843 14365 19852 14399
rect 19800 14356 19852 14365
rect 19248 14288 19300 14340
rect 11612 14220 11664 14229
rect 14832 14220 14884 14272
rect 16764 14220 16816 14272
rect 17408 14220 17460 14272
rect 19156 14220 19208 14272
rect 21180 14424 21232 14476
rect 21640 14424 21692 14476
rect 22560 14424 22612 14476
rect 22652 14467 22704 14476
rect 22652 14433 22661 14467
rect 22661 14433 22695 14467
rect 22695 14433 22704 14467
rect 22652 14424 22704 14433
rect 21088 14356 21140 14408
rect 20904 14220 20956 14272
rect 22744 14220 22796 14272
rect 4714 14118 4766 14170
rect 4778 14118 4830 14170
rect 4842 14118 4894 14170
rect 4906 14118 4958 14170
rect 12178 14118 12230 14170
rect 12242 14118 12294 14170
rect 12306 14118 12358 14170
rect 12370 14118 12422 14170
rect 19642 14118 19694 14170
rect 19706 14118 19758 14170
rect 19770 14118 19822 14170
rect 19834 14118 19886 14170
rect 1768 14016 1820 14068
rect 2872 13880 2924 13932
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 3240 14016 3292 14068
rect 3700 14059 3752 14068
rect 3700 14025 3709 14059
rect 3709 14025 3743 14059
rect 3743 14025 3752 14059
rect 3700 14016 3752 14025
rect 5816 14016 5868 14068
rect 5908 14016 5960 14068
rect 8760 14016 8812 14068
rect 10968 14016 11020 14068
rect 11520 14016 11572 14068
rect 11980 14016 12032 14068
rect 3976 13880 4028 13932
rect 4436 13880 4488 13932
rect 5172 13923 5224 13932
rect 5172 13889 5181 13923
rect 5181 13889 5215 13923
rect 5215 13889 5224 13923
rect 5172 13880 5224 13889
rect 5448 13880 5500 13932
rect 4068 13855 4120 13864
rect 2780 13812 2832 13821
rect 2964 13744 3016 13796
rect 4068 13821 4077 13855
rect 4077 13821 4111 13855
rect 4111 13821 4120 13855
rect 4068 13812 4120 13821
rect 4528 13855 4580 13864
rect 4528 13821 4537 13855
rect 4537 13821 4571 13855
rect 4571 13821 4580 13855
rect 4528 13812 4580 13821
rect 5540 13812 5592 13864
rect 8484 13855 8536 13864
rect 8484 13821 8502 13855
rect 8502 13821 8536 13855
rect 8484 13812 8536 13821
rect 8760 13855 8812 13864
rect 8760 13821 8769 13855
rect 8769 13821 8803 13855
rect 8803 13821 8812 13855
rect 9312 13880 9364 13932
rect 10876 13880 10928 13932
rect 13360 14016 13412 14068
rect 13820 14016 13872 14068
rect 14556 13948 14608 14000
rect 15476 13948 15528 14000
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 13360 13880 13412 13932
rect 18604 14016 18656 14068
rect 19248 14059 19300 14068
rect 19248 14025 19257 14059
rect 19257 14025 19291 14059
rect 19291 14025 19300 14059
rect 19248 14016 19300 14025
rect 22192 14059 22244 14068
rect 16396 13948 16448 14000
rect 8760 13812 8812 13821
rect 11704 13812 11756 13864
rect 12808 13855 12860 13864
rect 12808 13821 12826 13855
rect 12826 13821 12860 13855
rect 12808 13812 12860 13821
rect 12992 13812 13044 13864
rect 13728 13855 13780 13864
rect 6552 13744 6604 13796
rect 6184 13676 6236 13728
rect 7656 13676 7708 13728
rect 11336 13787 11388 13796
rect 11336 13753 11345 13787
rect 11345 13753 11379 13787
rect 11379 13753 11388 13787
rect 11336 13744 11388 13753
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 13728 13812 13780 13821
rect 16672 13923 16724 13932
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 17408 13923 17460 13932
rect 16672 13880 16724 13889
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 19432 13948 19484 14000
rect 20260 13948 20312 14000
rect 22192 14025 22201 14059
rect 22201 14025 22235 14059
rect 22235 14025 22244 14059
rect 22192 14016 22244 14025
rect 22284 13948 22336 14000
rect 17500 13880 17552 13889
rect 16488 13812 16540 13864
rect 17132 13812 17184 13864
rect 17776 13855 17828 13864
rect 17776 13821 17785 13855
rect 17785 13821 17819 13855
rect 17819 13821 17828 13855
rect 17776 13812 17828 13821
rect 19156 13880 19208 13932
rect 20076 13880 20128 13932
rect 22560 13880 22612 13932
rect 19248 13812 19300 13864
rect 20352 13812 20404 13864
rect 9864 13676 9916 13728
rect 10508 13719 10560 13728
rect 10508 13685 10517 13719
rect 10517 13685 10551 13719
rect 10551 13685 10560 13719
rect 10508 13676 10560 13685
rect 10784 13676 10836 13728
rect 16948 13719 17000 13728
rect 16948 13685 16957 13719
rect 16957 13685 16991 13719
rect 16991 13685 17000 13719
rect 16948 13676 17000 13685
rect 17316 13719 17368 13728
rect 17316 13685 17325 13719
rect 17325 13685 17359 13719
rect 17359 13685 17368 13719
rect 17316 13676 17368 13685
rect 17500 13676 17552 13728
rect 18328 13744 18380 13796
rect 20168 13787 20220 13796
rect 20168 13753 20177 13787
rect 20177 13753 20211 13787
rect 20211 13753 20220 13787
rect 20168 13744 20220 13753
rect 20444 13744 20496 13796
rect 20720 13812 20772 13864
rect 20904 13855 20956 13864
rect 20904 13821 20938 13855
rect 20938 13821 20956 13855
rect 20904 13812 20956 13821
rect 21456 13744 21508 13796
rect 21824 13744 21876 13796
rect 21640 13676 21692 13728
rect 22468 13744 22520 13796
rect 8446 13574 8498 13626
rect 8510 13574 8562 13626
rect 8574 13574 8626 13626
rect 8638 13574 8690 13626
rect 15910 13574 15962 13626
rect 15974 13574 16026 13626
rect 16038 13574 16090 13626
rect 16102 13574 16154 13626
rect 6184 13515 6236 13524
rect 6184 13481 6193 13515
rect 6193 13481 6227 13515
rect 6227 13481 6236 13515
rect 6184 13472 6236 13481
rect 6552 13515 6604 13524
rect 6552 13481 6561 13515
rect 6561 13481 6595 13515
rect 6595 13481 6604 13515
rect 6552 13472 6604 13481
rect 7932 13472 7984 13524
rect 5172 13404 5224 13456
rect 7656 13447 7708 13456
rect 7656 13413 7690 13447
rect 7690 13413 7708 13447
rect 7656 13404 7708 13413
rect 8300 13404 8352 13456
rect 9036 13472 9088 13524
rect 9864 13515 9916 13524
rect 9864 13481 9873 13515
rect 9873 13481 9907 13515
rect 9907 13481 9916 13515
rect 9864 13472 9916 13481
rect 11796 13472 11848 13524
rect 12808 13472 12860 13524
rect 4252 13379 4304 13388
rect 4252 13345 4261 13379
rect 4261 13345 4295 13379
rect 4295 13345 4304 13379
rect 4252 13336 4304 13345
rect 5448 13336 5500 13388
rect 11612 13404 11664 13456
rect 15108 13472 15160 13524
rect 17316 13472 17368 13524
rect 14924 13404 14976 13456
rect 18328 13472 18380 13524
rect 18604 13472 18656 13524
rect 18696 13404 18748 13456
rect 10600 13379 10652 13388
rect 10600 13345 10609 13379
rect 10609 13345 10643 13379
rect 10643 13345 10652 13379
rect 10600 13336 10652 13345
rect 11152 13336 11204 13388
rect 12532 13379 12584 13388
rect 12532 13345 12541 13379
rect 12541 13345 12575 13379
rect 12575 13345 12584 13379
rect 12532 13336 12584 13345
rect 13452 13336 13504 13388
rect 15016 13336 15068 13388
rect 16028 13379 16080 13388
rect 16028 13345 16037 13379
rect 16037 13345 16071 13379
rect 16071 13345 16080 13379
rect 16028 13336 16080 13345
rect 17408 13336 17460 13388
rect 18328 13336 18380 13388
rect 3240 13311 3292 13320
rect 3240 13277 3249 13311
rect 3249 13277 3283 13311
rect 3283 13277 3292 13311
rect 3240 13268 3292 13277
rect 4344 13311 4396 13320
rect 4344 13277 4353 13311
rect 4353 13277 4387 13311
rect 4387 13277 4396 13311
rect 4344 13268 4396 13277
rect 4436 13311 4488 13320
rect 4436 13277 4445 13311
rect 4445 13277 4479 13311
rect 4479 13277 4488 13311
rect 4436 13268 4488 13277
rect 4620 13268 4672 13320
rect 6644 13311 6696 13320
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 7288 13268 7340 13320
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 10876 13311 10928 13320
rect 10876 13277 10885 13311
rect 10885 13277 10919 13311
rect 10919 13277 10928 13311
rect 10876 13268 10928 13277
rect 17500 13311 17552 13320
rect 4528 13200 4580 13252
rect 10416 13200 10468 13252
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 18696 13268 18748 13320
rect 20812 13336 20864 13388
rect 22008 13336 22060 13388
rect 22376 13379 22428 13388
rect 22376 13345 22385 13379
rect 22385 13345 22419 13379
rect 22419 13345 22428 13379
rect 22376 13336 22428 13345
rect 12716 13243 12768 13252
rect 12716 13209 12725 13243
rect 12725 13209 12759 13243
rect 12759 13209 12768 13243
rect 12716 13200 12768 13209
rect 17132 13200 17184 13252
rect 17316 13200 17368 13252
rect 5908 13132 5960 13184
rect 6920 13132 6972 13184
rect 10232 13175 10284 13184
rect 10232 13141 10241 13175
rect 10241 13141 10275 13175
rect 10275 13141 10284 13175
rect 10232 13132 10284 13141
rect 14648 13132 14700 13184
rect 15752 13175 15804 13184
rect 15752 13141 15761 13175
rect 15761 13141 15795 13175
rect 15795 13141 15804 13175
rect 15752 13132 15804 13141
rect 16396 13132 16448 13184
rect 18880 13175 18932 13184
rect 18880 13141 18889 13175
rect 18889 13141 18923 13175
rect 18923 13141 18932 13175
rect 18880 13132 18932 13141
rect 19524 13132 19576 13184
rect 21088 13268 21140 13320
rect 22468 13311 22520 13320
rect 22468 13277 22477 13311
rect 22477 13277 22511 13311
rect 22511 13277 22520 13311
rect 22468 13268 22520 13277
rect 22836 13311 22888 13320
rect 22836 13277 22845 13311
rect 22845 13277 22879 13311
rect 22879 13277 22888 13311
rect 22836 13268 22888 13277
rect 20444 13132 20496 13184
rect 20812 13132 20864 13184
rect 21824 13175 21876 13184
rect 21824 13141 21833 13175
rect 21833 13141 21867 13175
rect 21867 13141 21876 13175
rect 21824 13132 21876 13141
rect 4714 13030 4766 13082
rect 4778 13030 4830 13082
rect 4842 13030 4894 13082
rect 4906 13030 4958 13082
rect 12178 13030 12230 13082
rect 12242 13030 12294 13082
rect 12306 13030 12358 13082
rect 12370 13030 12422 13082
rect 19642 13030 19694 13082
rect 19706 13030 19758 13082
rect 19770 13030 19822 13082
rect 19834 13030 19886 13082
rect 4344 12928 4396 12980
rect 5540 12971 5592 12980
rect 5540 12937 5549 12971
rect 5549 12937 5583 12971
rect 5583 12937 5592 12971
rect 5540 12928 5592 12937
rect 6552 12928 6604 12980
rect 7932 12971 7984 12980
rect 7932 12937 7941 12971
rect 7941 12937 7975 12971
rect 7975 12937 7984 12971
rect 7932 12928 7984 12937
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 14924 12928 14976 12980
rect 16028 12928 16080 12980
rect 5448 12903 5500 12912
rect 5448 12869 5457 12903
rect 5457 12869 5491 12903
rect 5491 12869 5500 12903
rect 5448 12860 5500 12869
rect 9312 12860 9364 12912
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 3884 12724 3936 12776
rect 4620 12724 4672 12776
rect 5908 12767 5960 12776
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 6736 12792 6788 12844
rect 10876 12792 10928 12844
rect 17776 12928 17828 12980
rect 20168 12928 20220 12980
rect 22560 12928 22612 12980
rect 16488 12792 16540 12844
rect 17132 12835 17184 12844
rect 17132 12801 17141 12835
rect 17141 12801 17175 12835
rect 17175 12801 17184 12835
rect 17132 12792 17184 12801
rect 19248 12860 19300 12912
rect 19524 12792 19576 12844
rect 20720 12860 20772 12912
rect 23480 12860 23532 12912
rect 3056 12656 3108 12708
rect 4252 12588 4304 12640
rect 5264 12656 5316 12708
rect 4436 12588 4488 12640
rect 6644 12724 6696 12776
rect 7288 12656 7340 12708
rect 8760 12724 8812 12776
rect 9036 12767 9088 12776
rect 9036 12733 9054 12767
rect 9054 12733 9088 12767
rect 9036 12724 9088 12733
rect 11152 12767 11204 12776
rect 11152 12733 11161 12767
rect 11161 12733 11195 12767
rect 11195 12733 11204 12767
rect 11152 12724 11204 12733
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 13452 12724 13504 12776
rect 15936 12767 15988 12776
rect 13176 12656 13228 12708
rect 14648 12656 14700 12708
rect 8760 12588 8812 12640
rect 9772 12631 9824 12640
rect 9772 12597 9781 12631
rect 9781 12597 9815 12631
rect 9815 12597 9824 12631
rect 9772 12588 9824 12597
rect 9864 12631 9916 12640
rect 9864 12597 9873 12631
rect 9873 12597 9907 12631
rect 9907 12597 9916 12631
rect 9864 12588 9916 12597
rect 11244 12631 11296 12640
rect 11244 12597 11253 12631
rect 11253 12597 11287 12631
rect 11287 12597 11296 12631
rect 11244 12588 11296 12597
rect 15936 12733 15954 12767
rect 15954 12733 15988 12767
rect 15936 12724 15988 12733
rect 16304 12767 16356 12776
rect 16304 12733 16313 12767
rect 16313 12733 16347 12767
rect 16347 12733 16356 12767
rect 16304 12724 16356 12733
rect 16764 12724 16816 12776
rect 17500 12724 17552 12776
rect 18880 12724 18932 12776
rect 15016 12588 15068 12640
rect 15752 12588 15804 12640
rect 17040 12656 17092 12708
rect 17592 12656 17644 12708
rect 19432 12656 19484 12708
rect 17684 12631 17736 12640
rect 17684 12597 17693 12631
rect 17693 12597 17727 12631
rect 17727 12597 17736 12631
rect 17684 12588 17736 12597
rect 19156 12631 19208 12640
rect 19156 12597 19165 12631
rect 19165 12597 19199 12631
rect 19199 12597 19208 12631
rect 19156 12588 19208 12597
rect 19248 12631 19300 12640
rect 19248 12597 19257 12631
rect 19257 12597 19291 12631
rect 19291 12597 19300 12631
rect 19616 12631 19668 12640
rect 19248 12588 19300 12597
rect 19616 12597 19625 12631
rect 19625 12597 19659 12631
rect 19659 12597 19668 12631
rect 19616 12588 19668 12597
rect 21916 12792 21968 12844
rect 22100 12792 22152 12844
rect 21640 12724 21692 12776
rect 21364 12656 21416 12708
rect 22652 12656 22704 12708
rect 22376 12631 22428 12640
rect 22376 12597 22385 12631
rect 22385 12597 22419 12631
rect 22419 12597 22428 12631
rect 22376 12588 22428 12597
rect 8446 12486 8498 12538
rect 8510 12486 8562 12538
rect 8574 12486 8626 12538
rect 8638 12486 8690 12538
rect 15910 12486 15962 12538
rect 15974 12486 16026 12538
rect 16038 12486 16090 12538
rect 16102 12486 16154 12538
rect 3240 12384 3292 12436
rect 2872 12316 2924 12368
rect 4436 12384 4488 12436
rect 5264 12427 5316 12436
rect 5264 12393 5273 12427
rect 5273 12393 5307 12427
rect 5307 12393 5316 12427
rect 5264 12384 5316 12393
rect 6644 12384 6696 12436
rect 6920 12384 6972 12436
rect 7380 12384 7432 12436
rect 8024 12384 8076 12436
rect 9864 12427 9916 12436
rect 9864 12393 9873 12427
rect 9873 12393 9907 12427
rect 9907 12393 9916 12427
rect 9864 12384 9916 12393
rect 10968 12384 11020 12436
rect 11244 12384 11296 12436
rect 11980 12427 12032 12436
rect 11980 12393 11989 12427
rect 11989 12393 12023 12427
rect 12023 12393 12032 12427
rect 11980 12384 12032 12393
rect 13636 12384 13688 12436
rect 15752 12384 15804 12436
rect 19432 12384 19484 12436
rect 19616 12427 19668 12436
rect 19616 12393 19625 12427
rect 19625 12393 19659 12427
rect 19659 12393 19668 12427
rect 19616 12384 19668 12393
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 4344 12316 4396 12368
rect 5908 12316 5960 12368
rect 7932 12316 7984 12368
rect 3056 12248 3108 12300
rect 4620 12248 4672 12300
rect 8852 12316 8904 12368
rect 8760 12248 8812 12300
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 3884 12223 3936 12232
rect 3884 12189 3893 12223
rect 3893 12189 3927 12223
rect 3927 12189 3936 12223
rect 3884 12180 3936 12189
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 7932 12180 7984 12232
rect 9404 12180 9456 12232
rect 11060 12316 11112 12368
rect 12072 12316 12124 12368
rect 16120 12316 16172 12368
rect 17132 12316 17184 12368
rect 10232 12248 10284 12300
rect 10508 12248 10560 12300
rect 11244 12248 11296 12300
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 13176 12248 13228 12300
rect 14740 12291 14792 12300
rect 14740 12257 14749 12291
rect 14749 12257 14783 12291
rect 14783 12257 14792 12291
rect 14740 12248 14792 12257
rect 15200 12291 15252 12300
rect 15200 12257 15209 12291
rect 15209 12257 15243 12291
rect 15243 12257 15252 12291
rect 15200 12248 15252 12257
rect 15476 12291 15528 12300
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 15660 12248 15712 12300
rect 10416 12180 10468 12232
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 15016 12223 15068 12232
rect 15016 12189 15025 12223
rect 15025 12189 15059 12223
rect 15059 12189 15068 12223
rect 15016 12180 15068 12189
rect 16396 12180 16448 12232
rect 13912 12112 13964 12164
rect 15108 12112 15160 12164
rect 17592 12248 17644 12300
rect 18512 12248 18564 12300
rect 17224 12223 17276 12232
rect 17224 12189 17233 12223
rect 17233 12189 17267 12223
rect 17267 12189 17276 12223
rect 17224 12180 17276 12189
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 16580 12112 16632 12164
rect 17132 12112 17184 12164
rect 17776 12180 17828 12232
rect 8300 12044 8352 12096
rect 8760 12044 8812 12096
rect 11888 12044 11940 12096
rect 14372 12087 14424 12096
rect 14372 12053 14381 12087
rect 14381 12053 14415 12087
rect 14415 12053 14424 12087
rect 14372 12044 14424 12053
rect 15292 12044 15344 12096
rect 16764 12044 16816 12096
rect 17960 12112 18012 12164
rect 21456 12316 21508 12368
rect 20720 12248 20772 12300
rect 21916 12316 21968 12368
rect 22744 12291 22796 12300
rect 22744 12257 22753 12291
rect 22753 12257 22787 12291
rect 22787 12257 22796 12291
rect 22744 12248 22796 12257
rect 22836 12291 22888 12300
rect 22836 12257 22845 12291
rect 22845 12257 22879 12291
rect 22879 12257 22888 12291
rect 22836 12248 22888 12257
rect 19064 12180 19116 12232
rect 17776 12044 17828 12096
rect 19524 12044 19576 12096
rect 19984 12044 20036 12096
rect 20444 12087 20496 12096
rect 20444 12053 20453 12087
rect 20453 12053 20487 12087
rect 20487 12053 20496 12087
rect 20444 12044 20496 12053
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 21364 12044 21416 12096
rect 21732 12044 21784 12096
rect 4714 11942 4766 11994
rect 4778 11942 4830 11994
rect 4842 11942 4894 11994
rect 4906 11942 4958 11994
rect 12178 11942 12230 11994
rect 12242 11942 12294 11994
rect 12306 11942 12358 11994
rect 12370 11942 12422 11994
rect 19642 11942 19694 11994
rect 19706 11942 19758 11994
rect 19770 11942 19822 11994
rect 19834 11942 19886 11994
rect 3056 11840 3108 11892
rect 4068 11840 4120 11892
rect 10508 11840 10560 11892
rect 10600 11840 10652 11892
rect 11060 11840 11112 11892
rect 14740 11840 14792 11892
rect 15108 11840 15160 11892
rect 16028 11840 16080 11892
rect 16120 11840 16172 11892
rect 17224 11840 17276 11892
rect 17868 11840 17920 11892
rect 18052 11883 18104 11892
rect 18052 11849 18061 11883
rect 18061 11849 18095 11883
rect 18095 11849 18104 11883
rect 18052 11840 18104 11849
rect 1400 11636 1452 11688
rect 2596 11636 2648 11688
rect 3884 11772 3936 11824
rect 10416 11772 10468 11824
rect 11152 11815 11204 11824
rect 11152 11781 11161 11815
rect 11161 11781 11195 11815
rect 11195 11781 11204 11815
rect 11152 11772 11204 11781
rect 14832 11772 14884 11824
rect 17960 11815 18012 11824
rect 3148 11568 3200 11620
rect 6920 11636 6972 11688
rect 8208 11636 8260 11688
rect 9404 11636 9456 11688
rect 13452 11747 13504 11756
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 9864 11636 9916 11688
rect 11980 11636 12032 11688
rect 14556 11636 14608 11688
rect 17132 11704 17184 11756
rect 17684 11704 17736 11756
rect 17960 11781 17969 11815
rect 17969 11781 18003 11815
rect 18003 11781 18012 11815
rect 17960 11772 18012 11781
rect 20444 11840 20496 11892
rect 20720 11840 20772 11892
rect 20996 11840 21048 11892
rect 22008 11883 22060 11892
rect 22008 11849 22017 11883
rect 22017 11849 22051 11883
rect 22051 11849 22060 11883
rect 22008 11840 22060 11849
rect 22192 11883 22244 11892
rect 22192 11849 22201 11883
rect 22201 11849 22235 11883
rect 22235 11849 22244 11883
rect 22192 11840 22244 11849
rect 16304 11636 16356 11688
rect 16488 11636 16540 11688
rect 16764 11679 16816 11688
rect 16764 11645 16773 11679
rect 16773 11645 16807 11679
rect 16807 11645 16816 11679
rect 16764 11636 16816 11645
rect 16948 11636 17000 11688
rect 17776 11679 17828 11688
rect 17776 11645 17785 11679
rect 17785 11645 17819 11679
rect 17819 11645 17828 11679
rect 17776 11636 17828 11645
rect 19156 11679 19208 11688
rect 19156 11645 19185 11679
rect 19185 11645 19208 11679
rect 19156 11636 19208 11645
rect 19432 11679 19484 11688
rect 19432 11645 19441 11679
rect 19441 11645 19475 11679
rect 19475 11645 19484 11679
rect 20168 11679 20220 11688
rect 19432 11636 19484 11645
rect 20168 11645 20177 11679
rect 20177 11645 20211 11679
rect 20211 11645 20220 11679
rect 20168 11636 20220 11645
rect 20444 11704 20496 11756
rect 20904 11747 20956 11756
rect 20904 11713 20913 11747
rect 20913 11713 20947 11747
rect 20947 11713 20956 11747
rect 20904 11704 20956 11713
rect 22560 11679 22612 11688
rect 22560 11645 22569 11679
rect 22569 11645 22603 11679
rect 22603 11645 22612 11679
rect 22560 11636 22612 11645
rect 6828 11568 6880 11620
rect 7932 11568 7984 11620
rect 8852 11611 8904 11620
rect 8852 11577 8886 11611
rect 8886 11577 8904 11611
rect 8852 11568 8904 11577
rect 8944 11568 8996 11620
rect 7380 11500 7432 11552
rect 8300 11500 8352 11552
rect 9956 11543 10008 11552
rect 9956 11509 9965 11543
rect 9965 11509 9999 11543
rect 9999 11509 10008 11543
rect 9956 11500 10008 11509
rect 10416 11543 10468 11552
rect 10416 11509 10425 11543
rect 10425 11509 10459 11543
rect 10459 11509 10468 11543
rect 10416 11500 10468 11509
rect 10508 11543 10560 11552
rect 10508 11509 10517 11543
rect 10517 11509 10551 11543
rect 10551 11509 10560 11543
rect 13636 11568 13688 11620
rect 14188 11568 14240 11620
rect 14924 11568 14976 11620
rect 19064 11568 19116 11620
rect 19340 11568 19392 11620
rect 10508 11500 10560 11509
rect 13544 11500 13596 11552
rect 16764 11500 16816 11552
rect 17224 11500 17276 11552
rect 19984 11500 20036 11552
rect 22652 11543 22704 11552
rect 22652 11509 22661 11543
rect 22661 11509 22695 11543
rect 22695 11509 22704 11543
rect 22652 11500 22704 11509
rect 8446 11398 8498 11450
rect 8510 11398 8562 11450
rect 8574 11398 8626 11450
rect 8638 11398 8690 11450
rect 15910 11398 15962 11450
rect 15974 11398 16026 11450
rect 16038 11398 16090 11450
rect 16102 11398 16154 11450
rect 3148 11296 3200 11348
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 8208 11296 8260 11348
rect 10508 11296 10560 11348
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 14188 11339 14240 11348
rect 14188 11305 14197 11339
rect 14197 11305 14231 11339
rect 14231 11305 14240 11339
rect 14188 11296 14240 11305
rect 8024 11228 8076 11280
rect 10416 11228 10468 11280
rect 15660 11271 15712 11280
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 1676 11203 1728 11212
rect 1676 11169 1710 11203
rect 1710 11169 1728 11203
rect 1676 11160 1728 11169
rect 7380 11160 7432 11212
rect 9220 11160 9272 11212
rect 15660 11237 15694 11271
rect 15694 11237 15712 11271
rect 15660 11228 15712 11237
rect 16856 11296 16908 11348
rect 17592 11339 17644 11348
rect 17592 11305 17601 11339
rect 17601 11305 17635 11339
rect 17635 11305 17644 11339
rect 17592 11296 17644 11305
rect 22652 11296 22704 11348
rect 12072 11160 12124 11212
rect 12900 11160 12952 11212
rect 8576 11092 8628 11144
rect 11152 11135 11204 11144
rect 11152 11101 11161 11135
rect 11161 11101 11195 11135
rect 11195 11101 11204 11135
rect 11152 11092 11204 11101
rect 15016 11135 15068 11144
rect 15016 11101 15025 11135
rect 15025 11101 15059 11135
rect 15059 11101 15068 11135
rect 15016 11092 15068 11101
rect 16488 11160 16540 11212
rect 13820 11024 13872 11076
rect 14556 10956 14608 11008
rect 17408 11092 17460 11144
rect 18052 11228 18104 11280
rect 18696 11228 18748 11280
rect 19156 11228 19208 11280
rect 20168 11228 20220 11280
rect 20628 11228 20680 11280
rect 21456 11228 21508 11280
rect 19248 11160 19300 11212
rect 20536 11160 20588 11212
rect 18052 11135 18104 11144
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 19340 11092 19392 11144
rect 19984 11092 20036 11144
rect 22560 11092 22612 11144
rect 16580 10956 16632 11008
rect 19984 10956 20036 11008
rect 20996 10956 21048 11008
rect 21916 10956 21968 11008
rect 22744 10956 22796 11008
rect 4714 10854 4766 10906
rect 4778 10854 4830 10906
rect 4842 10854 4894 10906
rect 4906 10854 4958 10906
rect 12178 10854 12230 10906
rect 12242 10854 12294 10906
rect 12306 10854 12358 10906
rect 12370 10854 12422 10906
rect 19642 10854 19694 10906
rect 19706 10854 19758 10906
rect 19770 10854 19822 10906
rect 19834 10854 19886 10906
rect 9864 10752 9916 10804
rect 10416 10752 10468 10804
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 12900 10752 12952 10804
rect 15660 10752 15712 10804
rect 17500 10752 17552 10804
rect 8576 10659 8628 10668
rect 8576 10625 8585 10659
rect 8585 10625 8619 10659
rect 8619 10625 8628 10659
rect 8576 10616 8628 10625
rect 8300 10591 8352 10600
rect 8300 10557 8318 10591
rect 8318 10557 8352 10591
rect 8300 10548 8352 10557
rect 8760 10548 8812 10600
rect 9220 10591 9272 10600
rect 9220 10557 9229 10591
rect 9229 10557 9263 10591
rect 9263 10557 9272 10591
rect 9220 10548 9272 10557
rect 9956 10548 10008 10600
rect 9404 10480 9456 10532
rect 12072 10616 12124 10668
rect 11428 10548 11480 10600
rect 14648 10548 14700 10600
rect 16672 10616 16724 10668
rect 19432 10752 19484 10804
rect 22376 10752 22428 10804
rect 23204 10684 23256 10736
rect 11244 10480 11296 10532
rect 15752 10480 15804 10532
rect 16304 10480 16356 10532
rect 17132 10548 17184 10600
rect 17224 10480 17276 10532
rect 19432 10616 19484 10668
rect 19800 10616 19852 10668
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 22192 10616 22244 10668
rect 22468 10616 22520 10668
rect 18972 10591 19024 10600
rect 18972 10557 18981 10591
rect 18981 10557 19015 10591
rect 19015 10557 19024 10591
rect 18972 10548 19024 10557
rect 19156 10548 19208 10600
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 19984 10548 20036 10557
rect 8760 10412 8812 10464
rect 14556 10412 14608 10464
rect 16580 10412 16632 10464
rect 17500 10412 17552 10464
rect 18052 10480 18104 10532
rect 18512 10412 18564 10464
rect 18696 10412 18748 10464
rect 18880 10412 18932 10464
rect 19340 10412 19392 10464
rect 19708 10455 19760 10464
rect 19708 10421 19723 10455
rect 19723 10421 19757 10455
rect 19757 10421 19760 10455
rect 19708 10412 19760 10421
rect 19892 10412 19944 10464
rect 22468 10480 22520 10532
rect 22652 10480 22704 10532
rect 20904 10412 20956 10464
rect 22376 10455 22428 10464
rect 22376 10421 22385 10455
rect 22385 10421 22419 10455
rect 22419 10421 22428 10455
rect 22376 10412 22428 10421
rect 8446 10310 8498 10362
rect 8510 10310 8562 10362
rect 8574 10310 8626 10362
rect 8638 10310 8690 10362
rect 15910 10310 15962 10362
rect 15974 10310 16026 10362
rect 16038 10310 16090 10362
rect 16102 10310 16154 10362
rect 8852 10208 8904 10260
rect 9956 10208 10008 10260
rect 10692 10208 10744 10260
rect 12072 10208 12124 10260
rect 15752 10251 15804 10260
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 16396 10208 16448 10260
rect 8760 10140 8812 10192
rect 10508 10140 10560 10192
rect 15292 10140 15344 10192
rect 16856 10183 16908 10192
rect 16856 10149 16874 10183
rect 16874 10149 16908 10183
rect 16856 10140 16908 10149
rect 9220 10072 9272 10124
rect 11152 10072 11204 10124
rect 13452 10072 13504 10124
rect 13544 10072 13596 10124
rect 18788 10208 18840 10260
rect 19984 10208 20036 10260
rect 21456 10208 21508 10260
rect 19432 10140 19484 10192
rect 19616 10140 19668 10192
rect 17408 10115 17460 10124
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 13176 10047 13228 10056
rect 13176 10013 13185 10047
rect 13185 10013 13219 10047
rect 13219 10013 13228 10047
rect 13176 10004 13228 10013
rect 9680 9936 9732 9988
rect 14096 9936 14148 9988
rect 17224 10004 17276 10056
rect 15476 9936 15528 9988
rect 20812 10072 20864 10124
rect 20904 10072 20956 10124
rect 23296 10072 23348 10124
rect 18328 10004 18380 10056
rect 18512 10004 18564 10056
rect 11612 9868 11664 9920
rect 12072 9868 12124 9920
rect 13912 9868 13964 9920
rect 14188 9911 14240 9920
rect 14188 9877 14197 9911
rect 14197 9877 14231 9911
rect 14231 9877 14240 9911
rect 14188 9868 14240 9877
rect 15384 9868 15436 9920
rect 15660 9911 15712 9920
rect 15660 9877 15669 9911
rect 15669 9877 15703 9911
rect 15703 9877 15712 9911
rect 15660 9868 15712 9877
rect 17224 9868 17276 9920
rect 19248 9868 19300 9920
rect 19616 10047 19668 10056
rect 19616 10013 19625 10047
rect 19625 10013 19659 10047
rect 19659 10013 19668 10047
rect 19616 10004 19668 10013
rect 20628 10004 20680 10056
rect 22836 10047 22888 10056
rect 22836 10013 22845 10047
rect 22845 10013 22879 10047
rect 22879 10013 22888 10047
rect 22836 10004 22888 10013
rect 20904 9868 20956 9920
rect 21824 9868 21876 9920
rect 4714 9766 4766 9818
rect 4778 9766 4830 9818
rect 4842 9766 4894 9818
rect 4906 9766 4958 9818
rect 12178 9766 12230 9818
rect 12242 9766 12294 9818
rect 12306 9766 12358 9818
rect 12370 9766 12422 9818
rect 19642 9766 19694 9818
rect 19706 9766 19758 9818
rect 19770 9766 19822 9818
rect 19834 9766 19886 9818
rect 9772 9596 9824 9648
rect 13452 9664 13504 9716
rect 14556 9664 14608 9716
rect 16304 9664 16356 9716
rect 16488 9639 16540 9648
rect 8300 9528 8352 9580
rect 12072 9528 12124 9580
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13176 9528 13228 9537
rect 9404 9460 9456 9512
rect 9864 9503 9916 9512
rect 9864 9469 9873 9503
rect 9873 9469 9907 9503
rect 9907 9469 9916 9503
rect 9864 9460 9916 9469
rect 8760 9392 8812 9444
rect 12164 9460 12216 9512
rect 13820 9528 13872 9580
rect 14004 9571 14056 9580
rect 14004 9537 14013 9571
rect 14013 9537 14047 9571
rect 14047 9537 14056 9571
rect 14004 9528 14056 9537
rect 14188 9528 14240 9580
rect 16488 9605 16497 9639
rect 16497 9605 16531 9639
rect 16531 9605 16540 9639
rect 16488 9596 16540 9605
rect 9680 9324 9732 9376
rect 11888 9324 11940 9376
rect 12716 9324 12768 9376
rect 12900 9435 12952 9444
rect 12900 9401 12918 9435
rect 12918 9401 12952 9435
rect 14372 9460 14424 9512
rect 14556 9460 14608 9512
rect 19340 9664 19392 9716
rect 22376 9664 22428 9716
rect 16856 9596 16908 9648
rect 18604 9639 18656 9648
rect 18604 9605 18613 9639
rect 18613 9605 18647 9639
rect 18647 9605 18656 9639
rect 18604 9596 18656 9605
rect 16304 9503 16356 9512
rect 12900 9392 12952 9401
rect 14004 9392 14056 9444
rect 16304 9469 16313 9503
rect 16313 9469 16347 9503
rect 16347 9469 16356 9503
rect 16304 9460 16356 9469
rect 18420 9528 18472 9580
rect 19064 9596 19116 9648
rect 21640 9596 21692 9648
rect 23388 9596 23440 9648
rect 18788 9528 18840 9580
rect 19432 9528 19484 9580
rect 19984 9528 20036 9580
rect 22744 9571 22796 9580
rect 22744 9537 22753 9571
rect 22753 9537 22787 9571
rect 22787 9537 22796 9571
rect 22744 9528 22796 9537
rect 17040 9460 17092 9512
rect 20076 9460 20128 9512
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 13728 9324 13780 9376
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 15016 9324 15068 9376
rect 16948 9367 17000 9376
rect 16948 9333 16957 9367
rect 16957 9333 16991 9367
rect 16991 9333 17000 9367
rect 16948 9324 17000 9333
rect 17316 9392 17368 9444
rect 17500 9435 17552 9444
rect 17500 9401 17534 9435
rect 17534 9401 17552 9435
rect 17500 9392 17552 9401
rect 17592 9392 17644 9444
rect 18144 9392 18196 9444
rect 19340 9392 19392 9444
rect 18420 9324 18472 9376
rect 18696 9367 18748 9376
rect 18696 9333 18705 9367
rect 18705 9333 18739 9367
rect 18739 9333 18748 9367
rect 18696 9324 18748 9333
rect 19064 9367 19116 9376
rect 19064 9333 19073 9367
rect 19073 9333 19107 9367
rect 19107 9333 19116 9367
rect 19064 9324 19116 9333
rect 19432 9324 19484 9376
rect 20260 9367 20312 9376
rect 20260 9333 20269 9367
rect 20269 9333 20303 9367
rect 20303 9333 20312 9367
rect 20260 9324 20312 9333
rect 22100 9460 22152 9512
rect 20996 9392 21048 9444
rect 21640 9392 21692 9444
rect 21548 9324 21600 9376
rect 22100 9324 22152 9376
rect 23296 9324 23348 9376
rect 8446 9222 8498 9274
rect 8510 9222 8562 9274
rect 8574 9222 8626 9274
rect 8638 9222 8690 9274
rect 15910 9222 15962 9274
rect 15974 9222 16026 9274
rect 16038 9222 16090 9274
rect 16102 9222 16154 9274
rect 1676 9120 1728 9172
rect 12808 9120 12860 9172
rect 13452 9163 13504 9172
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 14004 9120 14056 9172
rect 17500 9120 17552 9172
rect 1400 9027 1452 9036
rect 1400 8993 1409 9027
rect 1409 8993 1443 9027
rect 1443 8993 1452 9027
rect 9680 9052 9732 9104
rect 1400 8984 1452 8993
rect 9220 8984 9272 9036
rect 11336 8984 11388 9036
rect 11612 9052 11664 9104
rect 14096 9052 14148 9104
rect 12532 8984 12584 9036
rect 12716 8984 12768 9036
rect 15200 8984 15252 9036
rect 15752 9027 15804 9036
rect 15752 8993 15761 9027
rect 15761 8993 15795 9027
rect 15795 8993 15804 9027
rect 15752 8984 15804 8993
rect 16948 8984 17000 9036
rect 17960 9052 18012 9104
rect 11060 8916 11112 8968
rect 12900 8916 12952 8968
rect 13544 8916 13596 8968
rect 10508 8823 10560 8832
rect 10508 8789 10517 8823
rect 10517 8789 10551 8823
rect 10551 8789 10560 8823
rect 10508 8780 10560 8789
rect 11428 8780 11480 8832
rect 12624 8780 12676 8832
rect 13728 8848 13780 8900
rect 19340 9052 19392 9104
rect 18880 8984 18932 9036
rect 20076 9120 20128 9172
rect 22192 9120 22244 9172
rect 22468 9120 22520 9172
rect 20260 9052 20312 9104
rect 20904 9027 20956 9036
rect 13544 8780 13596 8832
rect 14648 8780 14700 8832
rect 16304 8823 16356 8832
rect 16304 8789 16313 8823
rect 16313 8789 16347 8823
rect 16347 8789 16356 8823
rect 16304 8780 16356 8789
rect 16580 8823 16632 8832
rect 16580 8789 16589 8823
rect 16589 8789 16623 8823
rect 16623 8789 16632 8823
rect 16580 8780 16632 8789
rect 16672 8780 16724 8832
rect 19524 8848 19576 8900
rect 19892 8848 19944 8900
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 18328 8780 18380 8832
rect 20904 8993 20913 9027
rect 20913 8993 20947 9027
rect 20947 8993 20956 9027
rect 20904 8984 20956 8993
rect 21815 9027 21867 9036
rect 21815 8993 21824 9027
rect 21824 8993 21858 9027
rect 21858 8993 21867 9027
rect 21815 8984 21867 8993
rect 22560 8984 22612 9036
rect 20260 8848 20312 8900
rect 20628 8916 20680 8968
rect 21180 8848 21232 8900
rect 20536 8780 20588 8832
rect 22468 8780 22520 8832
rect 4714 8678 4766 8730
rect 4778 8678 4830 8730
rect 4842 8678 4894 8730
rect 4906 8678 4958 8730
rect 12178 8678 12230 8730
rect 12242 8678 12294 8730
rect 12306 8678 12358 8730
rect 12370 8678 12422 8730
rect 19642 8678 19694 8730
rect 19706 8678 19758 8730
rect 19770 8678 19822 8730
rect 19834 8678 19886 8730
rect 1584 8576 1636 8628
rect 9220 8576 9272 8628
rect 11060 8619 11112 8628
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 11060 8585 11069 8619
rect 11069 8585 11103 8619
rect 11103 8585 11112 8619
rect 11060 8576 11112 8585
rect 13268 8576 13320 8628
rect 14096 8619 14148 8628
rect 14096 8585 14105 8619
rect 14105 8585 14139 8619
rect 14139 8585 14148 8619
rect 14096 8576 14148 8585
rect 18052 8576 18104 8628
rect 18788 8576 18840 8628
rect 21548 8576 21600 8628
rect 21732 8576 21784 8628
rect 22744 8576 22796 8628
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 7380 8372 7432 8424
rect 9680 8372 9732 8424
rect 10508 8372 10560 8424
rect 13084 8415 13136 8424
rect 11612 8304 11664 8356
rect 10784 8236 10836 8288
rect 12440 8304 12492 8356
rect 13084 8381 13093 8415
rect 13093 8381 13127 8415
rect 13127 8381 13136 8415
rect 13084 8372 13136 8381
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 16580 8508 16632 8560
rect 16672 8551 16724 8560
rect 16672 8517 16681 8551
rect 16681 8517 16715 8551
rect 16715 8517 16724 8551
rect 16948 8551 17000 8560
rect 16672 8508 16724 8517
rect 16948 8517 16957 8551
rect 16957 8517 16991 8551
rect 16991 8517 17000 8551
rect 16948 8508 17000 8517
rect 15752 8372 15804 8424
rect 14188 8304 14240 8356
rect 17592 8508 17644 8560
rect 18328 8508 18380 8560
rect 17960 8440 18012 8492
rect 18236 8440 18288 8492
rect 18144 8372 18196 8424
rect 18696 8440 18748 8492
rect 19156 8372 19208 8424
rect 19984 8372 20036 8424
rect 20628 8415 20680 8424
rect 20628 8381 20637 8415
rect 20637 8381 20671 8415
rect 20671 8381 20680 8415
rect 20628 8372 20680 8381
rect 17592 8347 17644 8356
rect 17592 8313 17601 8347
rect 17601 8313 17635 8347
rect 17635 8313 17644 8347
rect 17592 8304 17644 8313
rect 22376 8372 22428 8424
rect 20904 8347 20956 8356
rect 20904 8313 20938 8347
rect 20938 8313 20956 8347
rect 20904 8304 20956 8313
rect 13636 8279 13688 8288
rect 13636 8245 13645 8279
rect 13645 8245 13679 8279
rect 13679 8245 13688 8279
rect 13636 8236 13688 8245
rect 15200 8236 15252 8288
rect 15660 8236 15712 8288
rect 16856 8236 16908 8288
rect 18604 8236 18656 8288
rect 20628 8236 20680 8288
rect 21272 8236 21324 8288
rect 22100 8236 22152 8288
rect 22468 8236 22520 8288
rect 22560 8279 22612 8288
rect 22560 8245 22569 8279
rect 22569 8245 22603 8279
rect 22603 8245 22612 8279
rect 22560 8236 22612 8245
rect 8446 8134 8498 8186
rect 8510 8134 8562 8186
rect 8574 8134 8626 8186
rect 8638 8134 8690 8186
rect 15910 8134 15962 8186
rect 15974 8134 16026 8186
rect 16038 8134 16090 8186
rect 16102 8134 16154 8186
rect 9404 8032 9456 8084
rect 11336 8075 11388 8084
rect 11336 8041 11345 8075
rect 11345 8041 11379 8075
rect 11379 8041 11388 8075
rect 11336 8032 11388 8041
rect 10508 7964 10560 8016
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 13268 8075 13320 8084
rect 12440 8032 12492 8041
rect 13268 8041 13277 8075
rect 13277 8041 13311 8075
rect 13311 8041 13320 8075
rect 13268 8032 13320 8041
rect 14372 8032 14424 8084
rect 7380 7939 7432 7948
rect 7380 7905 7389 7939
rect 7389 7905 7423 7939
rect 7423 7905 7432 7939
rect 7380 7896 7432 7905
rect 10600 7828 10652 7880
rect 10784 7760 10836 7812
rect 10968 7939 11020 7948
rect 10968 7905 10977 7939
rect 10977 7905 11011 7939
rect 11011 7905 11020 7939
rect 11428 7939 11480 7948
rect 10968 7896 11020 7905
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 11980 7896 12032 7948
rect 12716 7896 12768 7948
rect 12900 7896 12952 7948
rect 14004 7939 14056 7948
rect 14004 7905 14013 7939
rect 14013 7905 14047 7939
rect 14047 7905 14056 7939
rect 14004 7896 14056 7905
rect 15200 7896 15252 7948
rect 15292 7939 15344 7948
rect 15292 7905 15301 7939
rect 15301 7905 15335 7939
rect 15335 7905 15344 7939
rect 16856 8032 16908 8084
rect 18328 8075 18380 8084
rect 18328 8041 18337 8075
rect 18337 8041 18371 8075
rect 18371 8041 18380 8075
rect 18328 8032 18380 8041
rect 19064 8032 19116 8084
rect 19432 8075 19484 8084
rect 19432 8041 19441 8075
rect 19441 8041 19475 8075
rect 19475 8041 19484 8075
rect 19432 8032 19484 8041
rect 22560 8032 22612 8084
rect 21732 7964 21784 8016
rect 17224 7939 17276 7948
rect 15292 7896 15344 7905
rect 17224 7905 17233 7939
rect 17233 7905 17267 7939
rect 17267 7905 17276 7939
rect 17224 7896 17276 7905
rect 17316 7896 17368 7948
rect 12992 7828 13044 7880
rect 14556 7871 14608 7880
rect 11888 7692 11940 7744
rect 12072 7735 12124 7744
rect 12072 7701 12081 7735
rect 12081 7701 12115 7735
rect 12115 7701 12124 7735
rect 12072 7692 12124 7701
rect 13636 7760 13688 7812
rect 14188 7735 14240 7744
rect 14188 7701 14197 7735
rect 14197 7701 14231 7735
rect 14231 7701 14240 7735
rect 14188 7692 14240 7701
rect 14556 7837 14565 7871
rect 14565 7837 14599 7871
rect 14599 7837 14608 7871
rect 14556 7828 14608 7837
rect 15016 7871 15068 7880
rect 15016 7837 15028 7871
rect 15028 7837 15062 7871
rect 15062 7837 15068 7871
rect 15016 7828 15068 7837
rect 16488 7871 16540 7880
rect 16488 7837 16497 7871
rect 16497 7837 16531 7871
rect 16531 7837 16540 7871
rect 16488 7828 16540 7837
rect 17592 7828 17644 7880
rect 18880 7871 18932 7880
rect 18880 7837 18889 7871
rect 18889 7837 18923 7871
rect 18923 7837 18932 7871
rect 18880 7828 18932 7837
rect 19156 7896 19208 7948
rect 19708 7828 19760 7880
rect 18144 7760 18196 7812
rect 19248 7760 19300 7812
rect 20076 7828 20128 7880
rect 20444 7828 20496 7880
rect 20628 7871 20680 7880
rect 20628 7837 20637 7871
rect 20637 7837 20671 7871
rect 20671 7837 20680 7871
rect 20628 7828 20680 7837
rect 20812 7828 20864 7880
rect 21272 7828 21324 7880
rect 21824 7939 21876 7948
rect 21824 7905 21833 7939
rect 21833 7905 21867 7939
rect 21867 7905 21876 7939
rect 22468 7939 22520 7948
rect 21824 7896 21876 7905
rect 22468 7905 22477 7939
rect 22477 7905 22511 7939
rect 22511 7905 22520 7939
rect 22468 7896 22520 7905
rect 22376 7871 22428 7880
rect 22376 7837 22385 7871
rect 22385 7837 22419 7871
rect 22419 7837 22428 7871
rect 22376 7828 22428 7837
rect 22928 7828 22980 7880
rect 22652 7760 22704 7812
rect 16948 7692 17000 7744
rect 18604 7692 18656 7744
rect 19156 7692 19208 7744
rect 20076 7692 20128 7744
rect 20444 7692 20496 7744
rect 21640 7692 21692 7744
rect 4714 7590 4766 7642
rect 4778 7590 4830 7642
rect 4842 7590 4894 7642
rect 4906 7590 4958 7642
rect 12178 7590 12230 7642
rect 12242 7590 12294 7642
rect 12306 7590 12358 7642
rect 12370 7590 12422 7642
rect 19642 7590 19694 7642
rect 19706 7590 19758 7642
rect 19770 7590 19822 7642
rect 19834 7590 19886 7642
rect 10508 7531 10560 7540
rect 10508 7497 10517 7531
rect 10517 7497 10551 7531
rect 10551 7497 10560 7531
rect 10508 7488 10560 7497
rect 10968 7488 11020 7540
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 14004 7488 14056 7540
rect 17592 7488 17644 7540
rect 18788 7488 18840 7540
rect 12624 7395 12676 7404
rect 12624 7361 12633 7395
rect 12633 7361 12667 7395
rect 12667 7361 12676 7395
rect 12624 7352 12676 7361
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14188 7352 14240 7361
rect 14372 7395 14424 7404
rect 14372 7361 14381 7395
rect 14381 7361 14415 7395
rect 14415 7361 14424 7395
rect 14372 7352 14424 7361
rect 15384 7352 15436 7404
rect 9404 7327 9456 7336
rect 9404 7293 9438 7327
rect 9438 7293 9456 7327
rect 9404 7284 9456 7293
rect 9680 7216 9732 7268
rect 11152 7216 11204 7268
rect 11244 7148 11296 7200
rect 12072 7284 12124 7336
rect 12256 7216 12308 7268
rect 13820 7259 13872 7268
rect 13820 7225 13829 7259
rect 13829 7225 13863 7259
rect 13863 7225 13872 7259
rect 13820 7216 13872 7225
rect 12992 7148 13044 7200
rect 15844 7352 15896 7404
rect 17132 7352 17184 7404
rect 17224 7352 17276 7404
rect 17592 7395 17644 7404
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 20536 7488 20588 7540
rect 20996 7488 21048 7540
rect 21732 7531 21784 7540
rect 21732 7497 21741 7531
rect 21741 7497 21775 7531
rect 21775 7497 21784 7531
rect 21732 7488 21784 7497
rect 22560 7488 22612 7540
rect 21640 7420 21692 7472
rect 22376 7395 22428 7404
rect 22376 7361 22385 7395
rect 22385 7361 22419 7395
rect 22419 7361 22428 7395
rect 22376 7352 22428 7361
rect 14556 7148 14608 7200
rect 15200 7191 15252 7200
rect 15200 7157 15209 7191
rect 15209 7157 15243 7191
rect 15243 7157 15252 7191
rect 15200 7148 15252 7157
rect 15292 7191 15344 7200
rect 15292 7157 15301 7191
rect 15301 7157 15335 7191
rect 15335 7157 15344 7191
rect 15660 7191 15712 7200
rect 15292 7148 15344 7157
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 16764 7148 16816 7200
rect 19616 7216 19668 7268
rect 19984 7284 20036 7336
rect 22100 7284 22152 7336
rect 20076 7259 20128 7268
rect 20076 7225 20085 7259
rect 20085 7225 20119 7259
rect 20119 7225 20128 7259
rect 20076 7216 20128 7225
rect 17316 7191 17368 7200
rect 17316 7157 17325 7191
rect 17325 7157 17359 7191
rect 17359 7157 17368 7191
rect 17316 7148 17368 7157
rect 17408 7148 17460 7200
rect 20444 7216 20496 7268
rect 20720 7216 20772 7268
rect 20996 7148 21048 7200
rect 21548 7148 21600 7200
rect 22192 7216 22244 7268
rect 8446 7046 8498 7098
rect 8510 7046 8562 7098
rect 8574 7046 8626 7098
rect 8638 7046 8690 7098
rect 15910 7046 15962 7098
rect 15974 7046 16026 7098
rect 16038 7046 16090 7098
rect 16102 7046 16154 7098
rect 10048 6944 10100 6996
rect 11244 6944 11296 6996
rect 12256 6987 12308 6996
rect 12256 6953 12265 6987
rect 12265 6953 12299 6987
rect 12299 6953 12308 6987
rect 12256 6944 12308 6953
rect 12992 6944 13044 6996
rect 10508 6876 10560 6928
rect 9680 6808 9732 6860
rect 11520 6808 11572 6860
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 13360 6808 13412 6860
rect 14372 6876 14424 6928
rect 15384 6808 15436 6860
rect 10600 6740 10652 6792
rect 10784 6740 10836 6792
rect 8944 6604 8996 6656
rect 11060 6740 11112 6792
rect 11152 6672 11204 6724
rect 12532 6740 12584 6792
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 20904 6944 20956 6996
rect 21732 6944 21784 6996
rect 19156 6876 19208 6928
rect 20628 6876 20680 6928
rect 17592 6808 17644 6860
rect 18788 6851 18840 6860
rect 18788 6817 18797 6851
rect 18797 6817 18831 6851
rect 18831 6817 18840 6851
rect 19340 6851 19392 6860
rect 18788 6808 18840 6817
rect 19340 6817 19349 6851
rect 19349 6817 19383 6851
rect 19383 6817 19392 6851
rect 19340 6808 19392 6817
rect 21640 6876 21692 6928
rect 15752 6740 15804 6792
rect 10968 6604 11020 6656
rect 15292 6604 15344 6656
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 17132 6672 17184 6724
rect 16212 6604 16264 6656
rect 16948 6604 17000 6656
rect 19984 6715 20036 6724
rect 19984 6681 19993 6715
rect 19993 6681 20027 6715
rect 20027 6681 20036 6715
rect 19984 6672 20036 6681
rect 20352 6783 20404 6792
rect 20352 6749 20361 6783
rect 20361 6749 20395 6783
rect 20395 6749 20404 6783
rect 20352 6740 20404 6749
rect 20444 6672 20496 6724
rect 20812 6740 20864 6792
rect 20628 6672 20680 6724
rect 21180 6740 21232 6792
rect 20812 6647 20864 6656
rect 20812 6613 20821 6647
rect 20821 6613 20855 6647
rect 20855 6613 20864 6647
rect 20812 6604 20864 6613
rect 21548 6808 21600 6860
rect 21640 6647 21692 6656
rect 21640 6613 21649 6647
rect 21649 6613 21683 6647
rect 21683 6613 21692 6647
rect 21640 6604 21692 6613
rect 22744 6604 22796 6656
rect 22836 6604 22888 6656
rect 4714 6502 4766 6554
rect 4778 6502 4830 6554
rect 4842 6502 4894 6554
rect 4906 6502 4958 6554
rect 12178 6502 12230 6554
rect 12242 6502 12294 6554
rect 12306 6502 12358 6554
rect 12370 6502 12422 6554
rect 19642 6502 19694 6554
rect 19706 6502 19758 6554
rect 19770 6502 19822 6554
rect 19834 6502 19886 6554
rect 10048 6443 10100 6452
rect 10048 6409 10057 6443
rect 10057 6409 10091 6443
rect 10091 6409 10100 6443
rect 10048 6400 10100 6409
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 12624 6400 12676 6452
rect 13820 6400 13872 6452
rect 9680 6264 9732 6316
rect 15384 6400 15436 6452
rect 17316 6400 17368 6452
rect 17960 6400 18012 6452
rect 19156 6400 19208 6452
rect 18880 6332 18932 6384
rect 20444 6400 20496 6452
rect 22652 6400 22704 6452
rect 8944 6239 8996 6248
rect 8944 6205 8978 6239
rect 8978 6205 8996 6239
rect 8944 6196 8996 6205
rect 13084 6196 13136 6248
rect 14372 6196 14424 6248
rect 19156 6264 19208 6316
rect 20720 6332 20772 6384
rect 20812 6332 20864 6384
rect 23112 6332 23164 6384
rect 11060 6128 11112 6180
rect 12532 6128 12584 6180
rect 13360 6128 13412 6180
rect 15476 6196 15528 6248
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 19432 6239 19484 6248
rect 19432 6205 19441 6239
rect 19441 6205 19475 6239
rect 19475 6205 19484 6239
rect 19432 6196 19484 6205
rect 22284 6239 22336 6248
rect 14740 6128 14792 6180
rect 17132 6128 17184 6180
rect 18236 6128 18288 6180
rect 18788 6128 18840 6180
rect 18972 6103 19024 6112
rect 18972 6069 18981 6103
rect 18981 6069 19015 6103
rect 19015 6069 19024 6103
rect 18972 6060 19024 6069
rect 20720 6128 20772 6180
rect 21732 6171 21784 6180
rect 21732 6137 21741 6171
rect 21741 6137 21775 6171
rect 21775 6137 21784 6171
rect 21732 6128 21784 6137
rect 21916 6171 21968 6180
rect 21916 6137 21925 6171
rect 21925 6137 21959 6171
rect 21959 6137 21968 6171
rect 21916 6128 21968 6137
rect 20628 6060 20680 6112
rect 20812 6103 20864 6112
rect 20812 6069 20821 6103
rect 20821 6069 20855 6103
rect 20855 6069 20864 6103
rect 20812 6060 20864 6069
rect 20904 6103 20956 6112
rect 20904 6069 20913 6103
rect 20913 6069 20947 6103
rect 20947 6069 20956 6103
rect 20904 6060 20956 6069
rect 21272 6060 21324 6112
rect 22284 6205 22293 6239
rect 22293 6205 22327 6239
rect 22327 6205 22336 6239
rect 22284 6196 22336 6205
rect 22744 6171 22796 6180
rect 22744 6137 22753 6171
rect 22753 6137 22787 6171
rect 22787 6137 22796 6171
rect 22744 6128 22796 6137
rect 23020 6060 23072 6112
rect 8446 5958 8498 6010
rect 8510 5958 8562 6010
rect 8574 5958 8626 6010
rect 8638 5958 8690 6010
rect 15910 5958 15962 6010
rect 15974 5958 16026 6010
rect 16038 5958 16090 6010
rect 16102 5958 16154 6010
rect 11060 5899 11112 5908
rect 11060 5865 11069 5899
rect 11069 5865 11103 5899
rect 11103 5865 11112 5899
rect 11060 5856 11112 5865
rect 12532 5899 12584 5908
rect 12532 5865 12541 5899
rect 12541 5865 12575 5899
rect 12575 5865 12584 5899
rect 12532 5856 12584 5865
rect 13544 5856 13596 5908
rect 15200 5856 15252 5908
rect 15660 5856 15712 5908
rect 17224 5856 17276 5908
rect 18512 5856 18564 5908
rect 18972 5856 19024 5908
rect 10048 5788 10100 5840
rect 11520 5788 11572 5840
rect 12624 5788 12676 5840
rect 13084 5788 13136 5840
rect 15568 5788 15620 5840
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 14556 5720 14608 5772
rect 14648 5763 14700 5772
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 15384 5763 15436 5772
rect 14648 5720 14700 5729
rect 15384 5729 15393 5763
rect 15393 5729 15427 5763
rect 15427 5729 15436 5763
rect 15384 5720 15436 5729
rect 15752 5652 15804 5704
rect 14740 5584 14792 5636
rect 16028 5720 16080 5772
rect 18052 5788 18104 5840
rect 20352 5856 20404 5908
rect 21548 5899 21600 5908
rect 21088 5831 21140 5840
rect 17868 5720 17920 5772
rect 21088 5797 21097 5831
rect 21097 5797 21131 5831
rect 21131 5797 21140 5831
rect 21088 5788 21140 5797
rect 21548 5865 21557 5899
rect 21557 5865 21591 5899
rect 21591 5865 21600 5899
rect 21548 5856 21600 5865
rect 22468 5788 22520 5840
rect 17684 5652 17736 5704
rect 19156 5720 19208 5772
rect 21640 5720 21692 5772
rect 22836 5720 22888 5772
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 17960 5584 18012 5636
rect 19524 5652 19576 5704
rect 20720 5584 20772 5636
rect 15476 5516 15528 5568
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 18512 5516 18564 5568
rect 20352 5516 20404 5568
rect 21456 5559 21508 5568
rect 21456 5525 21465 5559
rect 21465 5525 21499 5559
rect 21499 5525 21508 5559
rect 21456 5516 21508 5525
rect 22192 5516 22244 5568
rect 4714 5414 4766 5466
rect 4778 5414 4830 5466
rect 4842 5414 4894 5466
rect 4906 5414 4958 5466
rect 12178 5414 12230 5466
rect 12242 5414 12294 5466
rect 12306 5414 12358 5466
rect 12370 5414 12422 5466
rect 19642 5414 19694 5466
rect 19706 5414 19758 5466
rect 19770 5414 19822 5466
rect 19834 5414 19886 5466
rect 13360 5312 13412 5364
rect 17868 5312 17920 5364
rect 14740 5176 14792 5228
rect 15384 5176 15436 5228
rect 16948 5219 17000 5228
rect 16948 5185 16957 5219
rect 16957 5185 16991 5219
rect 16991 5185 17000 5219
rect 16948 5176 17000 5185
rect 18144 5176 18196 5228
rect 22376 5244 22428 5296
rect 13544 5108 13596 5160
rect 16304 5108 16356 5160
rect 17224 5151 17276 5160
rect 17224 5117 17258 5151
rect 17258 5117 17276 5151
rect 17224 5108 17276 5117
rect 18788 5108 18840 5160
rect 20812 5108 20864 5160
rect 20996 5219 21048 5228
rect 20996 5185 21005 5219
rect 21005 5185 21039 5219
rect 21039 5185 21048 5219
rect 20996 5176 21048 5185
rect 21548 5176 21600 5228
rect 22744 5219 22796 5228
rect 22744 5185 22753 5219
rect 22753 5185 22787 5219
rect 22787 5185 22796 5219
rect 22744 5176 22796 5185
rect 17960 4972 18012 5024
rect 18604 4972 18656 5024
rect 19984 4972 20036 5024
rect 20720 5015 20772 5024
rect 20720 4981 20729 5015
rect 20729 4981 20763 5015
rect 20763 4981 20772 5015
rect 20720 4972 20772 4981
rect 21088 4972 21140 5024
rect 22192 5108 22244 5160
rect 22284 5108 22336 5160
rect 21732 4972 21784 5024
rect 22100 4972 22152 5024
rect 22376 5040 22428 5092
rect 23388 5040 23440 5092
rect 22468 4972 22520 5024
rect 8446 4870 8498 4922
rect 8510 4870 8562 4922
rect 8574 4870 8626 4922
rect 8638 4870 8690 4922
rect 15910 4870 15962 4922
rect 15974 4870 16026 4922
rect 16038 4870 16090 4922
rect 16102 4870 16154 4922
rect 17684 4768 17736 4820
rect 18604 4811 18656 4820
rect 18604 4777 18613 4811
rect 18613 4777 18647 4811
rect 18647 4777 18656 4811
rect 18604 4768 18656 4777
rect 17868 4700 17920 4752
rect 20076 4700 20128 4752
rect 21364 4743 21416 4752
rect 21364 4709 21373 4743
rect 21373 4709 21407 4743
rect 21407 4709 21416 4743
rect 21364 4700 21416 4709
rect 22376 4700 22428 4752
rect 16120 4675 16172 4684
rect 16120 4641 16129 4675
rect 16129 4641 16163 4675
rect 16163 4641 16172 4675
rect 16120 4632 16172 4641
rect 17224 4632 17276 4684
rect 18328 4632 18380 4684
rect 18696 4632 18748 4684
rect 22560 4675 22612 4684
rect 22560 4641 22578 4675
rect 22578 4641 22612 4675
rect 22560 4632 22612 4641
rect 22836 4675 22888 4684
rect 22836 4641 22845 4675
rect 22845 4641 22879 4675
rect 22879 4641 22888 4675
rect 22836 4632 22888 4641
rect 23112 4675 23164 4684
rect 23112 4641 23121 4675
rect 23121 4641 23155 4675
rect 23155 4641 23164 4675
rect 23112 4632 23164 4641
rect 17776 4607 17828 4616
rect 17776 4573 17785 4607
rect 17785 4573 17819 4607
rect 17819 4573 17828 4607
rect 17776 4564 17828 4573
rect 18052 4607 18104 4616
rect 18052 4573 18061 4607
rect 18061 4573 18095 4607
rect 18095 4573 18104 4607
rect 18052 4564 18104 4573
rect 19156 4607 19208 4616
rect 19156 4573 19165 4607
rect 19165 4573 19199 4607
rect 19199 4573 19208 4607
rect 19156 4564 19208 4573
rect 19064 4496 19116 4548
rect 19524 4564 19576 4616
rect 20996 4564 21048 4616
rect 21364 4564 21416 4616
rect 20628 4496 20680 4548
rect 16672 4428 16724 4480
rect 20996 4471 21048 4480
rect 20996 4437 21005 4471
rect 21005 4437 21039 4471
rect 21039 4437 21048 4471
rect 20996 4428 21048 4437
rect 21548 4496 21600 4548
rect 4714 4326 4766 4378
rect 4778 4326 4830 4378
rect 4842 4326 4894 4378
rect 4906 4326 4958 4378
rect 12178 4326 12230 4378
rect 12242 4326 12294 4378
rect 12306 4326 12358 4378
rect 12370 4326 12422 4378
rect 19642 4326 19694 4378
rect 19706 4326 19758 4378
rect 19770 4326 19822 4378
rect 19834 4326 19886 4378
rect 16120 4224 16172 4276
rect 18788 4224 18840 4276
rect 21364 4224 21416 4276
rect 22192 4267 22244 4276
rect 18328 4199 18380 4208
rect 18328 4165 18337 4199
rect 18337 4165 18371 4199
rect 18371 4165 18380 4199
rect 18328 4156 18380 4165
rect 16948 4131 17000 4140
rect 16948 4097 16957 4131
rect 16957 4097 16991 4131
rect 16991 4097 17000 4131
rect 16948 4088 17000 4097
rect 19432 4088 19484 4140
rect 20444 4156 20496 4208
rect 20168 4131 20220 4140
rect 20168 4097 20177 4131
rect 20177 4097 20211 4131
rect 20211 4097 20220 4131
rect 20168 4088 20220 4097
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 22192 4233 22201 4267
rect 22201 4233 22235 4267
rect 22235 4233 22244 4267
rect 22192 4224 22244 4233
rect 22468 4156 22520 4208
rect 22284 4088 22336 4140
rect 16672 4020 16724 4072
rect 17224 4063 17276 4072
rect 17224 4029 17258 4063
rect 17258 4029 17276 4063
rect 17224 4020 17276 4029
rect 16488 3927 16540 3936
rect 16488 3893 16497 3927
rect 16497 3893 16531 3927
rect 16531 3893 16540 3927
rect 16488 3884 16540 3893
rect 17776 3952 17828 4004
rect 19524 4020 19576 4072
rect 20352 4063 20404 4072
rect 20352 4029 20361 4063
rect 20361 4029 20395 4063
rect 20395 4029 20404 4063
rect 20352 4020 20404 4029
rect 20628 4063 20680 4072
rect 20628 4029 20637 4063
rect 20637 4029 20671 4063
rect 20671 4029 20680 4063
rect 20628 4020 20680 4029
rect 18696 3995 18748 4004
rect 18696 3961 18730 3995
rect 18730 3961 18748 3995
rect 18696 3952 18748 3961
rect 21640 4020 21692 4072
rect 22560 4063 22612 4072
rect 22560 4029 22569 4063
rect 22569 4029 22603 4063
rect 22603 4029 22612 4063
rect 22560 4020 22612 4029
rect 21548 3952 21600 4004
rect 20076 3884 20128 3936
rect 20812 3884 20864 3936
rect 21180 3884 21232 3936
rect 21732 3884 21784 3936
rect 23296 3884 23348 3936
rect 8446 3782 8498 3834
rect 8510 3782 8562 3834
rect 8574 3782 8626 3834
rect 8638 3782 8690 3834
rect 15910 3782 15962 3834
rect 15974 3782 16026 3834
rect 16038 3782 16090 3834
rect 16102 3782 16154 3834
rect 4068 3612 4120 3664
rect 18328 3612 18380 3664
rect 18696 3680 18748 3732
rect 20352 3680 20404 3732
rect 20720 3680 20772 3732
rect 20904 3680 20956 3732
rect 22560 3680 22612 3732
rect 23020 3680 23072 3732
rect 19892 3655 19944 3664
rect 19892 3621 19901 3655
rect 19901 3621 19935 3655
rect 19935 3621 19944 3655
rect 19892 3612 19944 3621
rect 20260 3655 20312 3664
rect 20260 3621 20294 3655
rect 20294 3621 20312 3655
rect 20260 3612 20312 3621
rect 21088 3612 21140 3664
rect 17776 3544 17828 3596
rect 18512 3544 18564 3596
rect 19156 3544 19208 3596
rect 19524 3544 19576 3596
rect 20628 3544 20680 3596
rect 20812 3544 20864 3596
rect 22744 3612 22796 3664
rect 21732 3587 21784 3596
rect 21732 3553 21766 3587
rect 21766 3553 21784 3587
rect 21732 3544 21784 3553
rect 22100 3544 22152 3596
rect 3700 3383 3752 3392
rect 3700 3349 3709 3383
rect 3709 3349 3743 3383
rect 3743 3349 3752 3383
rect 3700 3340 3752 3349
rect 17224 3340 17276 3392
rect 19340 3340 19392 3392
rect 22836 3340 22888 3392
rect 4714 3238 4766 3290
rect 4778 3238 4830 3290
rect 4842 3238 4894 3290
rect 4906 3238 4958 3290
rect 12178 3238 12230 3290
rect 12242 3238 12294 3290
rect 12306 3238 12358 3290
rect 12370 3238 12422 3290
rect 19642 3238 19694 3290
rect 19706 3238 19758 3290
rect 19770 3238 19822 3290
rect 19834 3238 19886 3290
rect 1400 3111 1452 3120
rect 1400 3077 1409 3111
rect 1409 3077 1443 3111
rect 1443 3077 1452 3111
rect 1400 3068 1452 3077
rect 3700 3136 3752 3188
rect 16488 3136 16540 3188
rect 19340 3179 19392 3188
rect 19340 3145 19349 3179
rect 19349 3145 19383 3179
rect 19383 3145 19392 3179
rect 19340 3136 19392 3145
rect 20168 3136 20220 3188
rect 20444 3136 20496 3188
rect 17960 3068 18012 3120
rect 21180 3136 21232 3188
rect 19064 3043 19116 3052
rect 19064 3009 19073 3043
rect 19073 3009 19107 3043
rect 19107 3009 19116 3043
rect 19064 3000 19116 3009
rect 19432 3000 19484 3052
rect 21364 3000 21416 3052
rect 6092 2975 6144 2984
rect 2504 2839 2556 2848
rect 2504 2805 2513 2839
rect 2513 2805 2547 2839
rect 2547 2805 2556 2839
rect 2504 2796 2556 2805
rect 6092 2941 6101 2975
rect 6101 2941 6135 2975
rect 6135 2941 6144 2975
rect 6092 2932 6144 2941
rect 16948 2975 17000 2984
rect 16948 2941 16957 2975
rect 16957 2941 16991 2975
rect 16991 2941 17000 2975
rect 16948 2932 17000 2941
rect 17224 2975 17276 2984
rect 17224 2941 17258 2975
rect 17258 2941 17276 2975
rect 17224 2932 17276 2941
rect 20260 2932 20312 2984
rect 20812 2975 20864 2984
rect 20812 2941 20821 2975
rect 20821 2941 20855 2975
rect 20855 2941 20864 2975
rect 20812 2932 20864 2941
rect 20996 2932 21048 2984
rect 22836 2932 22888 2984
rect 3700 2864 3752 2916
rect 18236 2864 18288 2916
rect 19248 2864 19300 2916
rect 20444 2864 20496 2916
rect 22008 2864 22060 2916
rect 10692 2796 10744 2848
rect 17960 2796 18012 2848
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 20076 2796 20128 2848
rect 21916 2839 21968 2848
rect 21916 2805 21925 2839
rect 21925 2805 21959 2839
rect 21959 2805 21968 2839
rect 21916 2796 21968 2805
rect 23020 2839 23072 2848
rect 23020 2805 23029 2839
rect 23029 2805 23063 2839
rect 23063 2805 23072 2839
rect 23020 2796 23072 2805
rect 8446 2694 8498 2746
rect 8510 2694 8562 2746
rect 8574 2694 8626 2746
rect 8638 2694 8690 2746
rect 15910 2694 15962 2746
rect 15974 2694 16026 2746
rect 16038 2694 16090 2746
rect 16102 2694 16154 2746
rect 10692 2635 10744 2644
rect 10692 2601 10701 2635
rect 10701 2601 10735 2635
rect 10735 2601 10744 2635
rect 10692 2592 10744 2601
rect 18512 2592 18564 2644
rect 19156 2635 19208 2644
rect 19156 2601 19165 2635
rect 19165 2601 19199 2635
rect 19199 2601 19208 2635
rect 19156 2592 19208 2601
rect 22468 2592 22520 2644
rect 22652 2592 22704 2644
rect 2504 2524 2556 2576
rect 6092 2524 6144 2576
rect 18328 2524 18380 2576
rect 2044 2363 2096 2372
rect 2044 2329 2053 2363
rect 2053 2329 2087 2363
rect 2087 2329 2096 2363
rect 2044 2320 2096 2329
rect 6092 2363 6144 2372
rect 6092 2329 6101 2363
rect 6101 2329 6135 2363
rect 6135 2329 6144 2363
rect 6092 2320 6144 2329
rect 10232 2363 10284 2372
rect 10232 2329 10241 2363
rect 10241 2329 10275 2363
rect 10275 2329 10284 2363
rect 10232 2320 10284 2329
rect 14280 2252 14332 2304
rect 16948 2456 17000 2508
rect 17776 2456 17828 2508
rect 22008 2524 22060 2576
rect 19984 2499 20036 2508
rect 18420 2320 18472 2372
rect 19984 2465 19993 2499
rect 19993 2465 20027 2499
rect 20027 2465 20036 2499
rect 19984 2456 20036 2465
rect 20352 2499 20404 2508
rect 20352 2465 20361 2499
rect 20361 2465 20395 2499
rect 20395 2465 20404 2499
rect 20352 2456 20404 2465
rect 20720 2456 20772 2508
rect 20904 2499 20956 2508
rect 20904 2465 20938 2499
rect 20938 2465 20956 2499
rect 20904 2456 20956 2465
rect 21456 2456 21508 2508
rect 22192 2499 22244 2508
rect 22192 2465 22201 2499
rect 22201 2465 22235 2499
rect 22235 2465 22244 2499
rect 23204 2524 23256 2576
rect 22192 2456 22244 2465
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 22008 2388 22060 2440
rect 22836 2388 22888 2440
rect 20352 2320 20404 2372
rect 19432 2295 19484 2304
rect 19432 2261 19441 2295
rect 19441 2261 19475 2295
rect 19475 2261 19484 2295
rect 19432 2252 19484 2261
rect 21272 2252 21324 2304
rect 21732 2252 21784 2304
rect 4714 2150 4766 2202
rect 4778 2150 4830 2202
rect 4842 2150 4894 2202
rect 4906 2150 4958 2202
rect 12178 2150 12230 2202
rect 12242 2150 12294 2202
rect 12306 2150 12358 2202
rect 12370 2150 12422 2202
rect 19642 2150 19694 2202
rect 19706 2150 19758 2202
rect 19770 2150 19822 2202
rect 19834 2150 19886 2202
rect 19432 2048 19484 2100
rect 22192 2048 22244 2100
rect 20352 1980 20404 2032
rect 23480 1980 23532 2032
rect 23572 1411 23624 1420
rect 23572 1377 23581 1411
rect 23581 1377 23615 1411
rect 23615 1377 23624 1411
rect 23572 1368 23624 1377
<< metal2 >>
rect 294 23800 350 24600
rect 938 23800 994 24600
rect 1582 23800 1638 24600
rect 2226 23800 2282 24600
rect 2870 23800 2926 24600
rect 3514 23800 3570 24600
rect 4158 23800 4214 24600
rect 4802 23800 4858 24600
rect 5446 23800 5502 24600
rect 6090 23800 6146 24600
rect 6734 23800 6790 24600
rect 7378 23800 7434 24600
rect 8022 23800 8078 24600
rect 8666 23800 8722 24600
rect 9310 23800 9366 24600
rect 9954 23800 10010 24600
rect 10598 23800 10654 24600
rect 11242 23800 11298 24600
rect 11886 23800 11942 24600
rect 12530 23800 12586 24600
rect 13174 23800 13230 24600
rect 13818 23800 13874 24600
rect 14462 23800 14518 24600
rect 15106 23800 15162 24600
rect 15750 23800 15806 24600
rect 16394 23800 16450 24600
rect 17038 23800 17094 24600
rect 17682 23800 17738 24600
rect 18326 23800 18382 24600
rect 18970 23800 19026 24600
rect 19614 23800 19670 24600
rect 20258 23800 20314 24600
rect 20902 23800 20958 24600
rect 21546 23800 21602 24600
rect 21822 24304 21878 24313
rect 21822 24239 21878 24248
rect 308 22098 336 23800
rect 296 22092 348 22098
rect 296 22034 348 22040
rect 952 22030 980 23800
rect 1596 22250 1624 23800
rect 1596 22222 1716 22250
rect 1584 22092 1636 22098
rect 1584 22034 1636 22040
rect 940 22024 992 22030
rect 940 21966 992 21972
rect 1596 21690 1624 22034
rect 1688 21962 1716 22222
rect 1952 22092 2004 22098
rect 1952 22034 2004 22040
rect 1676 21956 1728 21962
rect 1676 21898 1728 21904
rect 1964 21690 1992 22034
rect 2240 22030 2268 23800
rect 2884 22098 2912 23800
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2688 22092 2740 22098
rect 2688 22034 2740 22040
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 3332 22092 3384 22098
rect 3332 22034 3384 22040
rect 2228 22024 2280 22030
rect 2228 21966 2280 21972
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1952 21684 2004 21690
rect 1952 21626 2004 21632
rect 2136 21548 2188 21554
rect 2136 21490 2188 21496
rect 1584 21480 1636 21486
rect 1582 21448 1584 21457
rect 1636 21448 1638 21457
rect 1582 21383 1638 21392
rect 2148 21010 2176 21490
rect 2332 21146 2360 22034
rect 2596 22024 2648 22030
rect 2596 21966 2648 21972
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 2424 21486 2452 21830
rect 2504 21616 2556 21622
rect 2502 21584 2504 21593
rect 2556 21584 2558 21593
rect 2502 21519 2558 21528
rect 2412 21480 2464 21486
rect 2412 21422 2464 21428
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2608 21078 2636 21966
rect 2700 21146 2728 22034
rect 3344 21690 3372 22034
rect 3528 21962 3556 23800
rect 4172 22098 4200 23800
rect 4816 22098 4844 23800
rect 5460 22438 5488 23800
rect 5448 22432 5500 22438
rect 5448 22374 5500 22380
rect 5908 22432 5960 22438
rect 5908 22374 5960 22380
rect 5920 22166 5948 22374
rect 5908 22160 5960 22166
rect 5908 22102 5960 22108
rect 4160 22092 4212 22098
rect 4160 22034 4212 22040
rect 4804 22092 4856 22098
rect 4804 22034 4856 22040
rect 5356 22092 5408 22098
rect 5356 22034 5408 22040
rect 6104 22080 6132 23800
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6276 22092 6328 22098
rect 6104 22052 6276 22080
rect 4528 22024 4580 22030
rect 3698 21992 3754 22001
rect 3516 21956 3568 21962
rect 4528 21966 4580 21972
rect 5368 21978 5396 22034
rect 3698 21927 3754 21936
rect 3516 21898 3568 21904
rect 3332 21684 3384 21690
rect 3332 21626 3384 21632
rect 3424 21412 3476 21418
rect 3424 21354 3476 21360
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 2596 21072 2648 21078
rect 2596 21014 2648 21020
rect 2136 21004 2188 21010
rect 2136 20946 2188 20952
rect 2872 21004 2924 21010
rect 2872 20946 2924 20952
rect 1674 20904 1730 20913
rect 1674 20839 1676 20848
rect 1728 20839 1730 20848
rect 1676 20810 1728 20816
rect 2148 20398 2176 20946
rect 2884 20602 2912 20946
rect 3436 20874 3464 21354
rect 3712 21010 3740 21927
rect 4160 21616 4212 21622
rect 4160 21558 4212 21564
rect 4172 21078 4200 21558
rect 4540 21486 4568 21966
rect 5368 21950 5580 21978
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 5448 21888 5500 21894
rect 5448 21830 5500 21836
rect 4688 21788 4984 21808
rect 4744 21786 4768 21788
rect 4824 21786 4848 21788
rect 4904 21786 4928 21788
rect 4766 21734 4768 21786
rect 4830 21734 4842 21786
rect 4904 21734 4906 21786
rect 4744 21732 4768 21734
rect 4824 21732 4848 21734
rect 4904 21732 4928 21734
rect 4688 21712 4984 21732
rect 4252 21480 4304 21486
rect 4436 21480 4488 21486
rect 4304 21440 4384 21468
rect 4252 21422 4304 21428
rect 4160 21072 4212 21078
rect 4160 21014 4212 21020
rect 3700 21004 3752 21010
rect 3700 20946 3752 20952
rect 3424 20868 3476 20874
rect 3424 20810 3476 20816
rect 2872 20596 2924 20602
rect 2872 20538 2924 20544
rect 4172 20398 4200 21014
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 2136 20392 2188 20398
rect 2136 20334 2188 20340
rect 2872 20392 2924 20398
rect 2872 20334 2924 20340
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 1676 20324 1728 20330
rect 1676 20266 1728 20272
rect 1688 20058 1716 20266
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 2148 19242 2176 20334
rect 2884 19836 2912 20334
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3712 20058 3740 20266
rect 4264 20262 4292 20742
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4252 20256 4304 20262
rect 4252 20198 4304 20204
rect 3700 20052 3752 20058
rect 3700 19994 3752 20000
rect 4080 19990 4108 20198
rect 4068 19984 4120 19990
rect 4068 19926 4120 19932
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 3516 19916 3568 19922
rect 3516 19858 3568 19864
rect 2964 19848 3016 19854
rect 2884 19808 2964 19836
rect 2964 19790 3016 19796
rect 1952 19236 2004 19242
rect 1952 19178 2004 19184
rect 2136 19236 2188 19242
rect 2136 19178 2188 19184
rect 2228 19236 2280 19242
rect 2228 19178 2280 19184
rect 1964 18970 1992 19178
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2148 18902 2176 19178
rect 2136 18896 2188 18902
rect 2136 18838 2188 18844
rect 1584 18624 1636 18630
rect 1584 18566 1636 18572
rect 1596 18290 1624 18566
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1780 17338 1808 17682
rect 2148 17678 2176 18838
rect 2240 18816 2268 19178
rect 3068 19174 3096 19858
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 19446 3188 19654
rect 3528 19514 3556 19858
rect 3516 19508 3568 19514
rect 3516 19450 3568 19456
rect 4356 19446 4384 21440
rect 4436 21422 4488 21428
rect 4528 21480 4580 21486
rect 4528 21422 4580 21428
rect 4448 21010 4476 21422
rect 5264 21412 5316 21418
rect 5264 21354 5316 21360
rect 5276 21146 5304 21354
rect 5368 21146 5396 21830
rect 5264 21140 5316 21146
rect 5264 21082 5316 21088
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 4688 20700 4984 20720
rect 4744 20698 4768 20700
rect 4824 20698 4848 20700
rect 4904 20698 4928 20700
rect 4766 20646 4768 20698
rect 4830 20646 4842 20698
rect 4904 20646 4906 20698
rect 4744 20644 4768 20646
rect 4824 20644 4848 20646
rect 4904 20644 4928 20646
rect 4688 20624 4984 20644
rect 4436 20460 4488 20466
rect 4436 20402 4488 20408
rect 4896 20460 4948 20466
rect 4896 20402 4948 20408
rect 3148 19440 3200 19446
rect 3148 19382 3200 19388
rect 4344 19440 4396 19446
rect 4344 19382 4396 19388
rect 4448 19378 4476 20402
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4632 20058 4660 20198
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4540 19378 4568 19790
rect 4724 19786 4752 20198
rect 4908 19854 4936 20402
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 4688 19612 4984 19632
rect 4744 19610 4768 19612
rect 4824 19610 4848 19612
rect 4904 19610 4928 19612
rect 4766 19558 4768 19610
rect 4830 19558 4842 19610
rect 4904 19558 4906 19610
rect 4744 19556 4768 19558
rect 4824 19556 4848 19558
rect 4904 19556 4928 19558
rect 4688 19536 4984 19556
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4528 19372 4580 19378
rect 4528 19314 4580 19320
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 3068 18902 3096 19110
rect 3056 18896 3108 18902
rect 3056 18838 3108 18844
rect 2320 18828 2372 18834
rect 2240 18788 2320 18816
rect 2240 18426 2268 18788
rect 2320 18770 2372 18776
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 3344 18222 3372 19110
rect 4356 18970 4384 19110
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3620 18426 3648 18770
rect 4448 18766 4476 19314
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3620 18222 3648 18362
rect 4448 18290 4476 18702
rect 4540 18630 4568 19314
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4816 18834 4844 19110
rect 5092 18970 5120 19722
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 4688 18524 4984 18544
rect 4744 18522 4768 18524
rect 4824 18522 4848 18524
rect 4904 18522 4928 18524
rect 4766 18470 4768 18522
rect 4830 18470 4842 18522
rect 4904 18470 4906 18522
rect 4744 18468 4768 18470
rect 4824 18468 4848 18470
rect 4904 18468 4928 18470
rect 4688 18448 4984 18468
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 3056 18216 3108 18222
rect 3056 18158 3108 18164
rect 3332 18216 3384 18222
rect 3332 18158 3384 18164
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3068 17882 3096 18158
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1780 15978 1808 17274
rect 3252 17202 3280 17614
rect 3344 17338 3372 18158
rect 3804 17814 3832 18158
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 3424 17808 3476 17814
rect 3424 17750 3476 17756
rect 3792 17808 3844 17814
rect 3792 17750 3844 17756
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3252 16794 3280 17138
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 2780 16720 2832 16726
rect 2780 16662 2832 16668
rect 2792 16046 2820 16662
rect 3436 16250 3464 17750
rect 4080 17610 4108 18022
rect 4448 17678 4476 18226
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 4080 17134 4108 17546
rect 4632 17270 4660 18226
rect 5092 18222 5120 18702
rect 5184 18426 5212 19858
rect 5460 19378 5488 21830
rect 5552 19718 5580 21950
rect 6104 21894 6132 22052
rect 6276 22034 6328 22040
rect 6656 21978 6684 22374
rect 6748 22094 6776 23800
rect 7392 22098 7420 23800
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7012 22094 7064 22098
rect 6748 22092 7064 22094
rect 6748 22066 7012 22092
rect 6656 21950 6776 21978
rect 6092 21888 6144 21894
rect 6092 21830 6144 21836
rect 6276 21888 6328 21894
rect 6276 21830 6328 21836
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5828 21078 5856 21286
rect 5816 21072 5868 21078
rect 5816 21014 5868 21020
rect 5828 20466 5856 21014
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5644 19310 5672 19994
rect 5736 19990 5764 20198
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 5736 19310 5764 19926
rect 5920 19514 5948 20198
rect 5908 19508 5960 19514
rect 5908 19450 5960 19456
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5724 19304 5776 19310
rect 5724 19246 5776 19252
rect 5816 19236 5868 19242
rect 5816 19178 5868 19184
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5276 18970 5304 19110
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5092 17882 5120 18158
rect 5080 17876 5132 17882
rect 5080 17818 5132 17824
rect 4688 17436 4984 17456
rect 4744 17434 4768 17436
rect 4824 17434 4848 17436
rect 4904 17434 4928 17436
rect 4766 17382 4768 17434
rect 4830 17382 4842 17434
rect 4904 17382 4906 17434
rect 4744 17380 4768 17382
rect 4824 17380 4848 17382
rect 4904 17380 4928 17382
rect 4688 17360 4984 17380
rect 5828 17338 5856 19178
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 4080 16454 4108 16934
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 1584 15972 1636 15978
rect 1584 15914 1636 15920
rect 1768 15972 1820 15978
rect 1768 15914 1820 15920
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15337 1532 15846
rect 1490 15328 1546 15337
rect 1490 15263 1546 15272
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11218 1440 11630
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1412 9042 1440 9143
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1596 8634 1624 15914
rect 2792 15706 2820 15982
rect 4080 15706 4108 16390
rect 4540 16046 4568 16390
rect 4632 16182 4660 16594
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 4688 16348 4984 16368
rect 4744 16346 4768 16348
rect 4824 16346 4848 16348
rect 4904 16346 4928 16348
rect 4766 16294 4768 16346
rect 4830 16294 4842 16346
rect 4904 16294 4906 16346
rect 4744 16292 4768 16294
rect 4824 16292 4848 16294
rect 4904 16292 4928 16294
rect 4688 16272 4984 16292
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 5460 16114 5488 16390
rect 6012 16114 6040 21626
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 6104 18630 6132 20402
rect 6184 18896 6236 18902
rect 6184 18838 6236 18844
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 6104 18154 6132 18566
rect 6092 18148 6144 18154
rect 6092 18090 6144 18096
rect 6104 17746 6132 18090
rect 6196 18086 6224 18838
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6104 16572 6132 17682
rect 6196 17134 6224 18022
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6196 16726 6224 16934
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6184 16584 6236 16590
rect 6104 16544 6184 16572
rect 6184 16526 6236 16532
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 6000 16108 6052 16114
rect 6000 16050 6052 16056
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 3516 15700 3568 15706
rect 4068 15700 4120 15706
rect 3516 15642 3568 15648
rect 3988 15660 4068 15688
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 1780 14074 1808 15506
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 2240 14278 2268 14826
rect 2884 14550 2912 15302
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2884 14090 2912 14486
rect 3160 14482 3188 14894
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 1768 14068 1820 14074
rect 2884 14062 3004 14090
rect 3252 14074 3280 15438
rect 3528 15026 3556 15642
rect 3988 15570 4016 15660
rect 4068 15642 4120 15648
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3712 14074 3740 15506
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3896 14482 3924 15302
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 3884 14476 3936 14482
rect 3884 14418 3936 14424
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 1768 14010 1820 14016
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2596 12776 2648 12782
rect 2792 12764 2820 13806
rect 2648 12736 2820 12764
rect 2596 12718 2648 12724
rect 2608 11694 2636 12718
rect 2884 12374 2912 13874
rect 2976 13802 3004 14062
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3988 13938 4016 14214
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 4080 13870 4108 14826
rect 4172 14618 4200 15846
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4540 15162 4568 15506
rect 4688 15260 4984 15280
rect 4744 15258 4768 15260
rect 4824 15258 4848 15260
rect 4904 15258 4928 15260
rect 4766 15206 4768 15258
rect 4830 15206 4842 15258
rect 4904 15206 4906 15258
rect 4744 15204 4768 15206
rect 4824 15204 4848 15206
rect 4904 15204 4928 15206
rect 4688 15184 4984 15204
rect 5184 15162 5212 15846
rect 5460 15638 5488 16050
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5908 15904 5960 15910
rect 5908 15846 5960 15852
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 5276 14958 5304 15302
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 5276 14550 5304 14894
rect 5264 14544 5316 14550
rect 5264 14486 5316 14492
rect 4688 14172 4984 14192
rect 4744 14170 4768 14172
rect 4824 14170 4848 14172
rect 4904 14170 4928 14172
rect 4766 14118 4768 14170
rect 4830 14118 4842 14170
rect 4904 14118 4906 14170
rect 4744 14116 4768 14118
rect 4824 14116 4848 14118
rect 4904 14116 4928 14118
rect 4688 14096 4984 14116
rect 5460 13938 5488 15574
rect 5828 14074 5856 15846
rect 5920 14074 5948 15846
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 6012 14890 6040 15506
rect 6000 14884 6052 14890
rect 6000 14826 6052 14832
rect 6012 14618 6040 14826
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 6288 14482 6316 21830
rect 6460 20800 6512 20806
rect 6460 20742 6512 20748
rect 6368 20324 6420 20330
rect 6368 20266 6420 20272
rect 6380 20058 6408 20266
rect 6368 20052 6420 20058
rect 6368 19994 6420 20000
rect 6472 19378 6500 20742
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6380 17542 6408 18770
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6380 16658 6408 17478
rect 6564 16726 6592 21830
rect 6656 21486 6684 21830
rect 6748 21690 6776 21950
rect 6736 21684 6788 21690
rect 6736 21626 6788 21632
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6644 20936 6696 20942
rect 6644 20878 6696 20884
rect 6656 20466 6684 20878
rect 6748 20806 6776 20946
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6840 20602 6868 22066
rect 7012 22034 7064 22040
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 6932 20398 6960 21490
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6656 19310 6684 20198
rect 6748 19990 6776 20198
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6840 18766 6868 19858
rect 6932 19378 6960 20198
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6840 17882 6868 18702
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6840 17202 6868 17818
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6840 16794 6868 16934
rect 6932 16794 6960 18022
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6552 16720 6604 16726
rect 6552 16662 6604 16668
rect 7024 16658 7052 17478
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6368 15972 6420 15978
rect 6368 15914 6420 15920
rect 6380 15162 6408 15914
rect 6748 15502 6776 15982
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6748 14414 6776 14962
rect 6840 14958 6868 15574
rect 6932 15026 6960 16118
rect 7012 15972 7064 15978
rect 7116 15960 7144 21830
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7208 17882 7236 19110
rect 7392 18834 7420 19246
rect 7484 19174 7512 22170
rect 7840 22092 7892 22098
rect 7840 22034 7892 22040
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7576 21457 7604 21966
rect 7562 21448 7618 21457
rect 7562 21383 7618 21392
rect 7576 20806 7604 21383
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7760 19310 7788 21966
rect 7852 21418 7880 22034
rect 7932 22024 7984 22030
rect 7932 21966 7984 21972
rect 7944 21690 7972 21966
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 7840 21412 7892 21418
rect 7840 21354 7892 21360
rect 7944 20398 7972 21626
rect 8036 20754 8064 23800
rect 8680 22930 8708 23800
rect 8680 22902 8892 22930
rect 8420 22332 8716 22352
rect 8476 22330 8500 22332
rect 8556 22330 8580 22332
rect 8636 22330 8660 22332
rect 8498 22278 8500 22330
rect 8562 22278 8574 22330
rect 8636 22278 8638 22330
rect 8476 22276 8500 22278
rect 8556 22276 8580 22278
rect 8636 22276 8660 22278
rect 8420 22256 8716 22276
rect 8300 22160 8352 22166
rect 8300 22102 8352 22108
rect 8116 21956 8168 21962
rect 8116 21898 8168 21904
rect 8128 21690 8156 21898
rect 8116 21684 8168 21690
rect 8116 21626 8168 21632
rect 8312 21060 8340 22102
rect 8760 22024 8812 22030
rect 8758 21992 8760 22001
rect 8812 21992 8814 22001
rect 8758 21927 8814 21936
rect 8574 21584 8630 21593
rect 8574 21519 8576 21528
rect 8628 21519 8630 21528
rect 8576 21490 8628 21496
rect 8392 21480 8444 21486
rect 8390 21448 8392 21457
rect 8760 21480 8812 21486
rect 8444 21448 8446 21457
rect 8760 21422 8812 21428
rect 8390 21383 8446 21392
rect 8420 21244 8716 21264
rect 8476 21242 8500 21244
rect 8556 21242 8580 21244
rect 8636 21242 8660 21244
rect 8498 21190 8500 21242
rect 8562 21190 8574 21242
rect 8636 21190 8638 21242
rect 8476 21188 8500 21190
rect 8556 21188 8580 21190
rect 8636 21188 8660 21190
rect 8420 21168 8716 21188
rect 8772 21146 8800 21422
rect 8864 21146 8892 22902
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 9036 21616 9088 21622
rect 9036 21558 9088 21564
rect 8944 21412 8996 21418
rect 8944 21354 8996 21360
rect 8760 21140 8812 21146
rect 8760 21082 8812 21088
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 8392 21072 8444 21078
rect 8312 21032 8392 21060
rect 8392 21014 8444 21020
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 8482 20904 8538 20913
rect 8404 20754 8432 20878
rect 8482 20839 8538 20848
rect 8496 20806 8524 20839
rect 8036 20726 8432 20754
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 7932 20392 7984 20398
rect 7932 20334 7984 20340
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 7840 20052 7892 20058
rect 7840 19994 7892 20000
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7380 18828 7432 18834
rect 7380 18770 7432 18776
rect 7760 18442 7788 19246
rect 7852 18902 7880 19994
rect 8312 19990 8340 20198
rect 8420 20156 8716 20176
rect 8476 20154 8500 20156
rect 8556 20154 8580 20156
rect 8636 20154 8660 20156
rect 8498 20102 8500 20154
rect 8562 20102 8574 20154
rect 8636 20102 8638 20154
rect 8476 20100 8500 20102
rect 8556 20100 8580 20102
rect 8636 20100 8660 20102
rect 8420 20080 8716 20100
rect 8772 20058 8800 20266
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 8128 18970 8156 19314
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 7840 18896 7892 18902
rect 7840 18838 7892 18844
rect 8312 18766 8340 19926
rect 8956 19922 8984 21354
rect 9048 20942 9076 21558
rect 9140 21418 9168 21966
rect 9128 21412 9180 21418
rect 9128 21354 9180 21360
rect 9324 21146 9352 23800
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9588 22160 9640 22166
rect 9588 22102 9640 22108
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 9600 21078 9628 22102
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9588 21072 9640 21078
rect 9588 21014 9640 21020
rect 9036 20936 9088 20942
rect 9036 20878 9088 20884
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 9048 19854 9076 20878
rect 9600 20602 9628 21014
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8588 19378 8616 19654
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8420 19068 8716 19088
rect 8476 19066 8500 19068
rect 8556 19066 8580 19068
rect 8636 19066 8660 19068
rect 8498 19014 8500 19066
rect 8562 19014 8574 19066
rect 8636 19014 8638 19066
rect 8476 19012 8500 19014
rect 8556 19012 8580 19014
rect 8636 19012 8660 19014
rect 8420 18992 8716 19012
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8772 18698 8800 19790
rect 9324 19666 9352 19858
rect 9232 19638 9352 19666
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9140 18902 9168 19450
rect 9128 18896 9180 18902
rect 9128 18838 9180 18844
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 7668 18426 7788 18442
rect 7656 18420 7788 18426
rect 7708 18414 7788 18420
rect 7656 18362 7708 18368
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7944 17814 7972 18566
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7196 17604 7248 17610
rect 7196 17546 7248 17552
rect 7208 16590 7236 17546
rect 7300 17134 7328 17682
rect 8312 17678 8340 18566
rect 8404 18290 8432 18566
rect 9048 18358 9076 18702
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8420 17980 8716 18000
rect 8476 17978 8500 17980
rect 8556 17978 8580 17980
rect 8636 17978 8660 17980
rect 8498 17926 8500 17978
rect 8562 17926 8574 17978
rect 8636 17926 8638 17978
rect 8476 17924 8500 17926
rect 8556 17924 8580 17926
rect 8636 17924 8660 17926
rect 8420 17904 8716 17924
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7196 16584 7248 16590
rect 7196 16526 7248 16532
rect 7064 15932 7144 15960
rect 7012 15914 7064 15920
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 7208 14550 7236 16526
rect 7300 14618 7328 17070
rect 7484 16794 7512 17138
rect 8208 17128 8260 17134
rect 8260 17076 8708 17082
rect 8208 17070 8708 17076
rect 8220 17066 8708 17070
rect 8220 17060 8720 17066
rect 8220 17054 8668 17060
rect 8668 17002 8720 17008
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 8300 16992 8352 16998
rect 8300 16934 8352 16940
rect 7852 16794 7880 16934
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7576 15570 7604 16186
rect 8036 16046 8064 16594
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7576 15026 7604 15506
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7944 14958 7972 15438
rect 8128 15094 8156 16390
rect 8312 16250 8340 16934
rect 8420 16892 8716 16912
rect 8476 16890 8500 16892
rect 8556 16890 8580 16892
rect 8636 16890 8660 16892
rect 8498 16838 8500 16890
rect 8562 16838 8574 16890
rect 8636 16838 8638 16890
rect 8476 16836 8500 16838
rect 8556 16836 8580 16838
rect 8636 16836 8660 16838
rect 8420 16816 8716 16836
rect 8484 16720 8536 16726
rect 8772 16674 8800 18226
rect 9048 18222 9076 18294
rect 9232 18222 9260 19638
rect 9416 19530 9444 19654
rect 9324 19502 9444 19530
rect 9324 19174 9352 19502
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9324 18766 9352 19110
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9036 18216 9088 18222
rect 9220 18216 9272 18222
rect 9088 18164 9168 18170
rect 9036 18158 9168 18164
rect 9220 18158 9272 18164
rect 9048 18142 9168 18158
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8536 16668 8800 16674
rect 8484 16662 8800 16668
rect 8496 16646 8800 16662
rect 8864 16590 8892 16934
rect 8944 16720 8996 16726
rect 8944 16662 8996 16668
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8956 16114 8984 16662
rect 9140 16114 9168 18142
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8220 15706 8248 15914
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8420 15804 8716 15824
rect 8476 15802 8500 15804
rect 8556 15802 8580 15804
rect 8636 15802 8660 15804
rect 8498 15750 8500 15802
rect 8562 15750 8574 15802
rect 8636 15750 8638 15802
rect 8476 15748 8500 15750
rect 8556 15748 8580 15750
rect 8636 15748 8660 15750
rect 8420 15728 8716 15748
rect 8772 15706 8800 15846
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8864 15162 8892 15846
rect 9232 15434 9260 18158
rect 9324 18086 9352 18702
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9324 17542 9352 18022
rect 9508 17898 9536 18566
rect 9416 17870 9536 17898
rect 9416 17678 9444 17870
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9324 15910 9352 17478
rect 9600 17338 9628 19178
rect 9692 19174 9720 22034
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9784 21146 9812 21966
rect 9876 21894 9904 22442
rect 9968 22438 9996 23800
rect 10612 22574 10640 23800
rect 10140 22568 10192 22574
rect 10140 22510 10192 22516
rect 10600 22568 10652 22574
rect 10600 22510 10652 22516
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 10046 22128 10102 22137
rect 10046 22063 10102 22072
rect 10060 21962 10088 22063
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9784 18970 9812 20198
rect 9876 19990 9904 21626
rect 10152 20330 10180 22510
rect 10784 22160 10836 22166
rect 10784 22102 10836 22108
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10428 21321 10456 21354
rect 10414 21312 10470 21321
rect 10414 21247 10470 21256
rect 10520 21010 10548 21966
rect 10612 21690 10640 21966
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10692 21480 10744 21486
rect 10690 21448 10692 21457
rect 10744 21448 10746 21457
rect 10690 21383 10746 21392
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10600 20392 10652 20398
rect 10600 20334 10652 20340
rect 10140 20324 10192 20330
rect 10140 20266 10192 20272
rect 10232 20324 10284 20330
rect 10232 20266 10284 20272
rect 10508 20324 10560 20330
rect 10508 20266 10560 20272
rect 9864 19984 9916 19990
rect 9864 19926 9916 19932
rect 10244 19378 10272 20266
rect 10520 20058 10548 20266
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 10612 19718 10640 20334
rect 10796 20058 10824 22102
rect 11060 22024 11112 22030
rect 11256 22001 11284 23800
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11624 22098 11652 22510
rect 11704 22228 11756 22234
rect 11704 22170 11756 22176
rect 11716 22137 11744 22170
rect 11702 22128 11758 22137
rect 11612 22092 11664 22098
rect 11900 22098 11928 23800
rect 12256 22432 12308 22438
rect 12256 22374 12308 22380
rect 12268 22098 12296 22374
rect 11702 22063 11758 22072
rect 11888 22092 11940 22098
rect 11612 22034 11664 22040
rect 12256 22092 12308 22098
rect 11888 22034 11940 22040
rect 11992 22052 12256 22080
rect 11060 21966 11112 21972
rect 11242 21992 11298 22001
rect 10876 21616 10928 21622
rect 10876 21558 10928 21564
rect 10966 21584 11022 21593
rect 10888 20602 10916 21558
rect 10966 21519 10968 21528
rect 11020 21519 11022 21528
rect 10968 21490 11020 21496
rect 10968 21412 11020 21418
rect 10968 21354 11020 21360
rect 10980 21026 11008 21354
rect 11072 21146 11100 21966
rect 11242 21927 11298 21936
rect 11428 21956 11480 21962
rect 11428 21898 11480 21904
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11256 21457 11284 21830
rect 11336 21480 11388 21486
rect 11242 21448 11298 21457
rect 11336 21422 11388 21428
rect 11242 21383 11298 21392
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11348 21078 11376 21422
rect 11336 21072 11388 21078
rect 10980 20998 11100 21026
rect 11336 21014 11388 21020
rect 11072 20806 11100 20998
rect 11336 20868 11388 20874
rect 11336 20810 11388 20816
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 11072 19990 11100 20742
rect 11348 20602 11376 20810
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11060 19984 11112 19990
rect 11060 19926 11112 19932
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10690 19408 10746 19417
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 10232 19372 10284 19378
rect 10232 19314 10284 19320
rect 10416 19372 10468 19378
rect 10690 19343 10692 19352
rect 10416 19314 10468 19320
rect 10744 19343 10746 19352
rect 10692 19314 10744 19320
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9692 18222 9720 18702
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9692 15706 9720 17206
rect 9876 16998 9904 19314
rect 10140 19168 10192 19174
rect 10140 19110 10192 19116
rect 10152 18834 10180 19110
rect 10140 18828 10192 18834
rect 10060 18788 10140 18816
rect 10060 18426 10088 18788
rect 10140 18770 10192 18776
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 10336 17134 10364 18702
rect 10428 17610 10456 19314
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10796 18970 10824 19110
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10888 18290 10916 19110
rect 10980 18698 11008 19790
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11072 18834 11100 19654
rect 11164 19446 11192 19654
rect 11152 19440 11204 19446
rect 11152 19382 11204 19388
rect 11336 19304 11388 19310
rect 11336 19246 11388 19252
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11164 18970 11192 19178
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 11072 17814 11100 18770
rect 11256 18290 11284 19110
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11060 17808 11112 17814
rect 11060 17750 11112 17756
rect 10416 17604 10468 17610
rect 10416 17546 10468 17552
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9784 15502 9812 16662
rect 10336 16114 10364 17070
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 9876 15706 9904 16050
rect 10520 15706 10548 16934
rect 11164 16590 11192 16934
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9862 15192 9918 15201
rect 8852 15156 8904 15162
rect 10060 15162 10088 15642
rect 10612 15502 10640 15642
rect 10796 15502 10824 16390
rect 11256 15994 11284 17818
rect 11348 17134 11376 19246
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11164 15966 11284 15994
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 9862 15127 9864 15136
rect 8852 15098 8904 15104
rect 9916 15127 9918 15136
rect 10048 15156 10100 15162
rect 9864 15098 9916 15104
rect 10048 15098 10100 15104
rect 8116 15088 8168 15094
rect 8116 15030 8168 15036
rect 9416 15026 9536 15042
rect 10152 15026 10180 15302
rect 11164 15201 11192 15966
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11256 15706 11284 15846
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11348 15638 11376 15846
rect 11336 15632 11388 15638
rect 11336 15574 11388 15580
rect 11150 15192 11206 15201
rect 11150 15127 11206 15136
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9404 15020 9536 15026
rect 9456 15014 9536 15020
rect 9404 14962 9456 14968
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 8420 14716 8716 14736
rect 8476 14714 8500 14716
rect 8556 14714 8580 14716
rect 8636 14714 8660 14716
rect 8498 14662 8500 14714
rect 8562 14662 8574 14714
rect 8636 14662 8638 14714
rect 8476 14660 8500 14662
rect 8556 14660 8580 14662
rect 8636 14660 8660 14662
rect 8420 14640 8716 14660
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 4068 13864 4120 13870
rect 4068 13806 4120 13812
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 3068 12306 3096 12650
rect 3252 12442 3280 13262
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3068 11898 3096 12242
rect 3896 12238 3924 12718
rect 4264 12646 4292 13330
rect 4448 13326 4476 13874
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4356 12986 4384 13262
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4356 12374 4384 12922
rect 4448 12646 4476 13262
rect 4540 13258 4568 13806
rect 5184 13462 5212 13874
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4632 12782 4660 13262
rect 4688 13084 4984 13104
rect 4744 13082 4768 13084
rect 4824 13082 4848 13084
rect 4904 13082 4928 13084
rect 4766 13030 4768 13082
rect 4830 13030 4842 13082
rect 4904 13030 4906 13082
rect 4744 13028 4768 13030
rect 4824 13028 4848 13030
rect 4904 13028 4928 13030
rect 4688 13008 4984 13028
rect 5460 12918 5488 13330
rect 5552 12986 5580 13806
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13530 6224 13670
rect 6564 13530 6592 13738
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5920 12782 5948 13126
rect 6564 12986 6592 13466
rect 6748 13326 6776 14350
rect 7208 13410 7236 14350
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8496 13870 8524 14214
rect 8772 14074 8800 14418
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 13462 7696 13670
rect 8420 13628 8716 13648
rect 8476 13626 8500 13628
rect 8556 13626 8580 13628
rect 8636 13626 8660 13628
rect 8498 13574 8500 13626
rect 8562 13574 8574 13626
rect 8636 13574 8638 13626
rect 8476 13572 8500 13574
rect 8556 13572 8580 13574
rect 8636 13572 8660 13574
rect 8420 13552 8716 13572
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7656 13456 7708 13462
rect 7208 13382 7328 13410
rect 7656 13398 7708 13404
rect 7300 13326 7328 13382
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6656 12782 6684 13262
rect 6748 12850 6776 13262
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6644 12776 6696 12782
rect 6644 12718 6696 12724
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4448 12442 4476 12582
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4632 12306 4660 12718
rect 5264 12708 5316 12714
rect 5264 12650 5316 12656
rect 5276 12442 5304 12650
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5920 12374 5948 12718
rect 6656 12442 6684 12718
rect 6932 12442 6960 13126
rect 7300 12714 7328 13262
rect 7944 12986 7972 13466
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 5908 12368 5960 12374
rect 7300 12322 7328 12650
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 5908 12310 5960 12316
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 6932 12294 7328 12322
rect 6932 12238 6960 12294
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 3160 11626 3188 12174
rect 3896 11830 3924 12174
rect 4688 11996 4984 12016
rect 4744 11994 4768 11996
rect 4824 11994 4848 11996
rect 4904 11994 4928 11996
rect 4766 11942 4768 11994
rect 4830 11942 4842 11994
rect 4904 11942 4906 11994
rect 4744 11940 4768 11942
rect 4824 11940 4848 11942
rect 4904 11940 4928 11942
rect 4688 11920 4984 11940
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 3884 11824 3936 11830
rect 3884 11766 3936 11772
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 3160 11354 3188 11562
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1688 9178 1716 11154
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 4080 3670 4108 11834
rect 6932 11694 6960 12174
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6840 11354 6868 11562
rect 7392 11558 7420 12378
rect 7944 12374 7972 12922
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7944 11626 7972 12174
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 7392 11218 7420 11494
rect 8036 11286 8064 12378
rect 8312 12102 8340 13398
rect 8772 12782 8800 13806
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8420 12540 8716 12560
rect 8476 12538 8500 12540
rect 8556 12538 8580 12540
rect 8636 12538 8660 12540
rect 8498 12486 8500 12538
rect 8562 12486 8574 12538
rect 8636 12486 8638 12538
rect 8476 12484 8500 12486
rect 8556 12484 8580 12486
rect 8636 12484 8660 12486
rect 8420 12464 8716 12484
rect 8772 12306 8800 12582
rect 8864 12434 8892 14350
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9048 12782 9076 13466
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8864 12406 8984 12434
rect 8864 12374 8892 12406
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8220 11354 8248 11630
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8024 11280 8076 11286
rect 8024 11222 8076 11228
rect 7380 11212 7432 11218
rect 7380 11154 7432 11160
rect 4688 10908 4984 10928
rect 4744 10906 4768 10908
rect 4824 10906 4848 10908
rect 4904 10906 4928 10908
rect 4766 10854 4768 10906
rect 4830 10854 4842 10906
rect 4904 10854 4906 10906
rect 4744 10852 4768 10854
rect 4824 10852 4848 10854
rect 4904 10852 4928 10854
rect 4688 10832 4984 10852
rect 8312 10606 8340 11494
rect 8420 11452 8716 11472
rect 8476 11450 8500 11452
rect 8556 11450 8580 11452
rect 8636 11450 8660 11452
rect 8498 11398 8500 11450
rect 8562 11398 8574 11450
rect 8636 11398 8638 11450
rect 8476 11396 8500 11398
rect 8556 11396 8580 11398
rect 8636 11396 8660 11398
rect 8420 11376 8716 11396
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8588 10674 8616 11086
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8772 10606 8800 12038
rect 8956 11626 8984 12406
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 4688 9820 4984 9840
rect 4744 9818 4768 9820
rect 4824 9818 4848 9820
rect 4904 9818 4928 9820
rect 4766 9766 4768 9818
rect 4830 9766 4842 9818
rect 4904 9766 4906 9818
rect 4744 9764 4768 9766
rect 4824 9764 4848 9766
rect 4904 9764 4928 9766
rect 4688 9744 4984 9764
rect 8312 9586 8340 10542
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8420 10364 8716 10384
rect 8476 10362 8500 10364
rect 8556 10362 8580 10364
rect 8636 10362 8660 10364
rect 8498 10310 8500 10362
rect 8562 10310 8574 10362
rect 8636 10310 8638 10362
rect 8476 10308 8500 10310
rect 8556 10308 8580 10310
rect 8636 10308 8660 10310
rect 8420 10288 8716 10308
rect 8772 10198 8800 10406
rect 8864 10266 8892 11562
rect 9232 11218 9260 14962
rect 9508 14940 9536 15014
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 11336 14952 11388 14958
rect 9508 14912 9720 14940
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9416 14346 9444 14826
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9324 13326 9352 13874
rect 9692 13433 9720 14912
rect 11336 14894 11388 14900
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10980 14521 11008 14758
rect 10966 14512 11022 14521
rect 10966 14447 11022 14456
rect 11072 14414 11100 14758
rect 11244 14544 11296 14550
rect 11244 14486 11296 14492
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10796 13977 10824 14350
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10782 13968 10838 13977
rect 10782 13903 10838 13912
rect 10876 13932 10928 13938
rect 10796 13818 10824 13903
rect 10876 13874 10928 13880
rect 10428 13790 10824 13818
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 13530 9904 13670
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9678 13424 9734 13433
rect 9678 13359 9734 13368
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9324 12918 9352 13262
rect 10428 13258 10456 13790
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10416 13252 10468 13258
rect 10416 13194 10468 13200
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9324 12434 9352 12854
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9324 12406 9444 12434
rect 9416 12238 9444 12406
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9416 11694 9444 12174
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8772 9450 8800 10134
rect 9232 10130 9260 10542
rect 9416 10538 9444 11630
rect 9404 10532 9456 10538
rect 9404 10474 9456 10480
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9416 10062 9444 10474
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9416 9518 9444 9998
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 9692 9382 9720 9930
rect 9784 9654 9812 12582
rect 9876 12442 9904 12582
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 10244 12306 10272 13126
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10428 12238 10456 13194
rect 10520 12306 10548 13670
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10506 12200 10562 12209
rect 10428 11830 10456 12174
rect 10506 12135 10562 12144
rect 10520 11898 10548 12135
rect 10612 11898 10640 13330
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10508 11892 10560 11898
rect 10508 11834 10560 11840
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9876 10810 9904 11630
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9876 9518 9904 10746
rect 9968 10606 9996 11494
rect 10428 11286 10456 11494
rect 10520 11354 10548 11494
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10428 10810 10456 11222
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9968 10266 9996 10542
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10520 10198 10548 11290
rect 10704 10266 10732 13262
rect 10796 12986 10824 13670
rect 10888 13326 10916 13874
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10888 12850 10916 13262
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10980 12442 11008 14010
rect 11256 13512 11284 14486
rect 11348 13802 11376 14894
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11072 13484 11284 13512
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 11072 12374 11100 13484
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11164 12782 11192 13330
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 11164 11914 11192 12718
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11256 12442 11284 12582
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11072 11898 11192 11914
rect 11060 11892 11192 11898
rect 11112 11886 11192 11892
rect 11060 11834 11112 11840
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11164 11150 11192 11766
rect 11256 11354 11284 12242
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 11164 10130 11192 11086
rect 11256 10538 11284 11290
rect 11440 10606 11468 21898
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11624 21554 11652 21830
rect 11796 21684 11848 21690
rect 11900 21672 11928 22034
rect 11848 21644 11928 21672
rect 11796 21626 11848 21632
rect 11702 21584 11758 21593
rect 11612 21548 11664 21554
rect 11702 21519 11704 21528
rect 11612 21490 11664 21496
rect 11756 21519 11758 21528
rect 11704 21490 11756 21496
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11520 20392 11572 20398
rect 11520 20334 11572 20340
rect 11532 19514 11560 20334
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 11532 17066 11560 17614
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11532 15094 11560 15506
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 11624 14822 11652 21286
rect 11992 20058 12020 22052
rect 12544 22094 12572 23800
rect 13188 22098 13216 23800
rect 13832 22166 13860 23800
rect 14476 22234 14504 23800
rect 15120 22574 15148 23800
rect 15108 22568 15160 22574
rect 15108 22510 15160 22516
rect 15016 22432 15068 22438
rect 15016 22374 15068 22380
rect 15028 22234 15056 22374
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 15016 22228 15068 22234
rect 15016 22170 15068 22176
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 12716 22094 12768 22098
rect 12544 22092 12768 22094
rect 12544 22066 12716 22092
rect 12256 22034 12308 22040
rect 12716 22034 12768 22040
rect 12808 22092 12860 22098
rect 12808 22034 12860 22040
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 13176 22092 13228 22098
rect 13176 22034 13228 22040
rect 12532 21888 12584 21894
rect 12532 21830 12584 21836
rect 12152 21788 12448 21808
rect 12208 21786 12232 21788
rect 12288 21786 12312 21788
rect 12368 21786 12392 21788
rect 12230 21734 12232 21786
rect 12294 21734 12306 21786
rect 12368 21734 12370 21786
rect 12208 21732 12232 21734
rect 12288 21732 12312 21734
rect 12368 21732 12392 21734
rect 12152 21712 12448 21732
rect 12346 21584 12402 21593
rect 12346 21519 12402 21528
rect 12360 21486 12388 21519
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12072 21412 12124 21418
rect 12072 21354 12124 21360
rect 12084 21078 12112 21354
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 12346 21040 12402 21049
rect 12346 20975 12348 20984
rect 12400 20975 12402 20984
rect 12348 20946 12400 20952
rect 12152 20700 12448 20720
rect 12208 20698 12232 20700
rect 12288 20698 12312 20700
rect 12368 20698 12392 20700
rect 12230 20646 12232 20698
rect 12294 20646 12306 20698
rect 12368 20646 12370 20698
rect 12208 20644 12232 20646
rect 12288 20644 12312 20646
rect 12368 20644 12392 20646
rect 12152 20624 12448 20644
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12152 19612 12448 19632
rect 12208 19610 12232 19612
rect 12288 19610 12312 19612
rect 12368 19610 12392 19612
rect 12230 19558 12232 19610
rect 12294 19558 12306 19610
rect 12368 19558 12370 19610
rect 12208 19556 12232 19558
rect 12288 19556 12312 19558
rect 12368 19556 12392 19558
rect 12152 19536 12448 19556
rect 11796 19304 11848 19310
rect 11702 19272 11758 19281
rect 11796 19246 11848 19252
rect 11702 19207 11758 19216
rect 11716 18902 11744 19207
rect 11704 18896 11756 18902
rect 11704 18838 11756 18844
rect 11808 18766 11836 19246
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12176 18834 12204 19110
rect 12164 18828 12216 18834
rect 12084 18788 12164 18816
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 12084 18358 12112 18788
rect 12164 18770 12216 18776
rect 12152 18524 12448 18544
rect 12208 18522 12232 18524
rect 12288 18522 12312 18524
rect 12368 18522 12392 18524
rect 12230 18470 12232 18522
rect 12294 18470 12306 18522
rect 12368 18470 12370 18522
rect 12208 18468 12232 18470
rect 12288 18468 12312 18470
rect 12368 18468 12392 18470
rect 12152 18448 12448 18468
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11808 16726 11836 17138
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11716 15366 11744 16594
rect 11808 15366 11836 16662
rect 11992 16046 12020 17070
rect 11980 16040 12032 16046
rect 11900 16000 11980 16028
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11900 15094 11928 16000
rect 11980 15982 12032 15988
rect 11888 15088 11940 15094
rect 11888 15030 11940 15036
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11624 14634 11652 14758
rect 11624 14606 11744 14634
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11624 14362 11652 14418
rect 11716 14414 11744 14606
rect 11532 14334 11652 14362
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11532 14074 11560 14334
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11624 13462 11652 14214
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11716 10810 11744 13806
rect 11808 13530 11836 14758
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11900 12102 11928 14894
rect 11992 14550 12020 14962
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11992 14074 12020 14486
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11992 11694 12020 12378
rect 12084 12374 12112 17682
rect 12152 17436 12448 17456
rect 12208 17434 12232 17436
rect 12288 17434 12312 17436
rect 12368 17434 12392 17436
rect 12230 17382 12232 17434
rect 12294 17382 12306 17434
rect 12368 17382 12370 17434
rect 12208 17380 12232 17382
rect 12288 17380 12312 17382
rect 12368 17380 12392 17382
rect 12152 17360 12448 17380
rect 12152 16348 12448 16368
rect 12208 16346 12232 16348
rect 12288 16346 12312 16348
rect 12368 16346 12392 16348
rect 12230 16294 12232 16346
rect 12294 16294 12306 16346
rect 12368 16294 12370 16346
rect 12208 16292 12232 16294
rect 12288 16292 12312 16294
rect 12368 16292 12392 16294
rect 12152 16272 12448 16292
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12176 15502 12204 16118
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12152 15260 12448 15280
rect 12208 15258 12232 15260
rect 12288 15258 12312 15260
rect 12368 15258 12392 15260
rect 12230 15206 12232 15258
rect 12294 15206 12306 15258
rect 12368 15206 12370 15258
rect 12208 15204 12232 15206
rect 12288 15204 12312 15206
rect 12368 15204 12392 15206
rect 12152 15184 12448 15204
rect 12544 14958 12572 21830
rect 12624 21004 12676 21010
rect 12624 20946 12676 20952
rect 12636 20262 12664 20946
rect 12728 20602 12756 22034
rect 12820 22001 12848 22034
rect 12806 21992 12862 22001
rect 12806 21927 12862 21936
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12820 20482 12848 21927
rect 13004 21690 13032 22034
rect 13176 21956 13228 21962
rect 13176 21898 13228 21904
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12912 21350 12940 21422
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12912 21010 12940 21286
rect 12900 21004 12952 21010
rect 12900 20946 12952 20952
rect 12728 20454 12848 20482
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12728 18086 12756 20454
rect 12912 20380 12940 20946
rect 12992 20392 13044 20398
rect 12912 20352 12992 20380
rect 12992 20334 13044 20340
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 12820 19854 12848 20266
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12912 20058 12940 20198
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 13096 19938 13124 21830
rect 13004 19910 13124 19938
rect 13188 19922 13216 21898
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13280 20398 13308 21830
rect 13542 21584 13598 21593
rect 13542 21519 13598 21528
rect 13360 21412 13412 21418
rect 13360 21354 13412 21360
rect 13372 21146 13400 21354
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13358 21040 13414 21049
rect 13358 20975 13414 20984
rect 13372 20806 13400 20975
rect 13452 20936 13504 20942
rect 13452 20878 13504 20884
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13268 20392 13320 20398
rect 13268 20334 13320 20340
rect 13464 20330 13492 20878
rect 13556 20482 13584 21519
rect 13648 20602 13676 22102
rect 15028 22098 15056 22170
rect 14372 22092 14424 22098
rect 14372 22034 14424 22040
rect 15016 22092 15068 22098
rect 15016 22034 15068 22040
rect 15384 22092 15436 22098
rect 15764 22094 15792 23800
rect 16212 22568 16264 22574
rect 16212 22510 16264 22516
rect 15884 22332 16180 22352
rect 15940 22330 15964 22332
rect 16020 22330 16044 22332
rect 16100 22330 16124 22332
rect 15962 22278 15964 22330
rect 16026 22278 16038 22330
rect 16100 22278 16102 22330
rect 15940 22276 15964 22278
rect 16020 22276 16044 22278
rect 16100 22276 16124 22278
rect 15884 22256 16180 22276
rect 16224 22166 16252 22510
rect 16212 22160 16264 22166
rect 16264 22120 16344 22148
rect 16212 22102 16264 22108
rect 15384 22034 15436 22040
rect 15580 22080 15792 22094
rect 16028 22092 16080 22098
rect 15580 22066 16028 22080
rect 13728 22024 13780 22030
rect 13728 21966 13780 21972
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13740 21146 13768 21966
rect 13924 21146 13952 21966
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13556 20454 13676 20482
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 13176 19916 13228 19922
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12900 19780 12952 19786
rect 12900 19722 12952 19728
rect 12912 19378 12940 19722
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12912 17678 12940 19314
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12912 16046 12940 16526
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12624 15972 12676 15978
rect 12624 15914 12676 15920
rect 12636 15706 12664 15914
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12728 15706 12756 15846
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12716 15700 12768 15706
rect 12716 15642 12768 15648
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12164 14952 12216 14958
rect 12532 14952 12584 14958
rect 12216 14912 12296 14940
rect 12164 14894 12216 14900
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12176 14346 12204 14758
rect 12268 14550 12296 14912
rect 12532 14894 12584 14900
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12152 14172 12448 14192
rect 12208 14170 12232 14172
rect 12288 14170 12312 14172
rect 12368 14170 12392 14172
rect 12230 14118 12232 14170
rect 12294 14118 12306 14170
rect 12368 14118 12370 14170
rect 12208 14116 12232 14118
rect 12288 14116 12312 14118
rect 12368 14116 12392 14118
rect 12152 14096 12448 14116
rect 12544 13394 12572 14350
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12728 13258 12756 15438
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12820 13870 12848 14826
rect 13004 13870 13032 19910
rect 13176 19858 13228 19864
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13096 19514 13124 19790
rect 13464 19786 13492 20266
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13268 19236 13320 19242
rect 13268 19178 13320 19184
rect 13280 18970 13308 19178
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13096 18290 13124 18566
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13096 17134 13124 17614
rect 13372 17338 13400 17682
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 13096 16794 13124 17070
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13176 16652 13228 16658
rect 13176 16594 13228 16600
rect 13188 15978 13216 16594
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 14958 13400 15846
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13372 14074 13400 14350
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13082 13968 13138 13977
rect 13082 13903 13084 13912
rect 13136 13903 13138 13912
rect 13360 13932 13412 13938
rect 13084 13874 13136 13880
rect 13360 13874 13412 13880
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 12820 13530 12848 13806
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12152 13084 12448 13104
rect 12208 13082 12232 13084
rect 12288 13082 12312 13084
rect 12368 13082 12392 13084
rect 12230 13030 12232 13082
rect 12294 13030 12306 13082
rect 12368 13030 12370 13082
rect 12208 13028 12232 13030
rect 12288 13028 12312 13030
rect 12368 13028 12392 13030
rect 12152 13008 12448 13028
rect 13372 12782 13400 13874
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13464 12782 13492 13330
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 13188 12306 13216 12650
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 12268 12209 12296 12242
rect 12254 12200 12310 12209
rect 12254 12135 12310 12144
rect 12152 11996 12448 12016
rect 12208 11994 12232 11996
rect 12288 11994 12312 11996
rect 12368 11994 12392 11996
rect 12230 11942 12232 11994
rect 12294 11942 12306 11994
rect 12368 11942 12370 11994
rect 12208 11940 12232 11942
rect 12288 11940 12312 11942
rect 12368 11940 12392 11942
rect 12152 11920 12448 11940
rect 13464 11762 13492 12718
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 13556 11558 13584 17478
rect 13648 16726 13676 20454
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 13832 19990 13860 20266
rect 13924 19990 13952 21082
rect 14016 21078 14044 21830
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 14108 21146 14136 21422
rect 14280 21412 14332 21418
rect 14280 21354 14332 21360
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 14004 21072 14056 21078
rect 14004 21014 14056 21020
rect 14108 20942 14136 21082
rect 14186 21040 14242 21049
rect 14186 20975 14242 20984
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14200 20874 14228 20975
rect 14188 20868 14240 20874
rect 14188 20810 14240 20816
rect 14292 20398 14320 21354
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14384 20058 14412 22034
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 14648 21616 14700 21622
rect 14648 21558 14700 21564
rect 14462 21312 14518 21321
rect 14462 21247 14518 21256
rect 14476 21010 14504 21247
rect 14660 21078 14688 21558
rect 14648 21072 14700 21078
rect 14648 21014 14700 21020
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14660 20398 14688 21014
rect 14752 20466 14780 21830
rect 15304 21486 15332 21830
rect 15396 21690 15424 22034
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15108 21412 15160 21418
rect 15108 21354 15160 21360
rect 15120 21146 15148 21354
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15292 21072 15344 21078
rect 15292 21014 15344 21020
rect 14924 20528 14976 20534
rect 14924 20470 14976 20476
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13912 19984 13964 19990
rect 14556 19984 14608 19990
rect 13964 19932 14044 19938
rect 13912 19926 14044 19932
rect 14556 19926 14608 19932
rect 13924 19910 14044 19926
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13740 18290 13768 19314
rect 13924 19174 13952 19790
rect 14016 19378 14044 19910
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 13912 19168 13964 19174
rect 13912 19110 13964 19116
rect 14016 18902 14044 19314
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13820 18692 13872 18698
rect 13820 18634 13872 18640
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13832 17882 13860 18634
rect 13924 18426 13952 18770
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 14292 17814 14320 18022
rect 14280 17808 14332 17814
rect 14280 17750 14332 17756
rect 14384 17746 14412 18566
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14476 16794 14504 19654
rect 14568 18970 14596 19926
rect 14752 19854 14780 20402
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14660 18834 14688 19110
rect 14844 18970 14872 19858
rect 14936 19718 14964 20470
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15016 20256 15068 20262
rect 15016 20198 15068 20204
rect 15028 20058 15056 20198
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 15212 19718 15240 20334
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15304 19334 15332 21014
rect 14936 19306 15332 19334
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14752 18426 14780 18770
rect 14936 18766 14964 19306
rect 15488 19281 15516 21830
rect 15580 19786 15608 22066
rect 15764 22052 16028 22066
rect 16028 22034 16080 22040
rect 16212 21616 16264 21622
rect 16212 21558 16264 21564
rect 16028 21548 16080 21554
rect 16028 21490 16080 21496
rect 16040 21332 16068 21490
rect 15764 21304 16068 21332
rect 15660 21072 15712 21078
rect 15764 21060 15792 21304
rect 15884 21244 16180 21264
rect 15940 21242 15964 21244
rect 16020 21242 16044 21244
rect 16100 21242 16124 21244
rect 15962 21190 15964 21242
rect 16026 21190 16038 21242
rect 16100 21190 16102 21242
rect 15940 21188 15964 21190
rect 16020 21188 16044 21190
rect 16100 21188 16124 21190
rect 15884 21168 16180 21188
rect 15712 21032 15792 21060
rect 15844 21072 15896 21078
rect 15660 21014 15712 21020
rect 15844 21014 15896 21020
rect 15672 20942 15700 21014
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15856 20806 15884 21014
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 16224 20466 16252 21558
rect 16316 20602 16344 22120
rect 16408 22094 16436 23800
rect 17052 22098 17080 23800
rect 17408 22500 17460 22506
rect 17408 22442 17460 22448
rect 17420 22166 17448 22442
rect 17408 22160 17460 22166
rect 17408 22102 17460 22108
rect 16488 22094 16540 22098
rect 16408 22092 16540 22094
rect 16408 22066 16488 22092
rect 16488 22034 16540 22040
rect 16580 22092 16632 22098
rect 16580 22034 16632 22040
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16408 21078 16436 21626
rect 16396 21072 16448 21078
rect 16396 21014 16448 21020
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 15884 20156 16180 20176
rect 15940 20154 15964 20156
rect 16020 20154 16044 20156
rect 16100 20154 16124 20156
rect 15962 20102 15964 20154
rect 16026 20102 16038 20154
rect 16100 20102 16102 20154
rect 15940 20100 15964 20102
rect 16020 20100 16044 20102
rect 16100 20100 16124 20102
rect 15884 20080 16180 20100
rect 16224 19922 16252 20198
rect 16408 20058 16436 20198
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16500 19990 16528 22034
rect 16592 21690 16620 22034
rect 17696 21962 17724 23800
rect 17960 22160 18012 22166
rect 17960 22102 18012 22108
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 16764 21888 16816 21894
rect 16948 21888 17000 21894
rect 16764 21830 16816 21836
rect 16868 21848 16948 21876
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16776 21554 16804 21830
rect 16764 21548 16816 21554
rect 16764 21490 16816 21496
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16488 19984 16540 19990
rect 16488 19926 16540 19932
rect 16592 19922 16620 20742
rect 16868 20482 16896 21848
rect 16948 21830 17000 21836
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16960 20942 16988 21422
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 17316 21412 17368 21418
rect 17316 21354 17368 21360
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 17236 20806 17264 21354
rect 17328 21049 17356 21354
rect 17314 21040 17370 21049
rect 17314 20975 17370 20984
rect 17224 20800 17276 20806
rect 17224 20742 17276 20748
rect 17972 20602 18000 22102
rect 18340 21690 18368 23800
rect 18420 22500 18472 22506
rect 18420 22442 18472 22448
rect 18328 21684 18380 21690
rect 18328 21626 18380 21632
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 18064 21457 18092 21558
rect 18050 21448 18106 21457
rect 18050 21383 18106 21392
rect 18432 20942 18460 22442
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18892 22234 18920 22374
rect 18880 22228 18932 22234
rect 18880 22170 18932 22176
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18616 21146 18644 21422
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18512 20868 18564 20874
rect 18512 20810 18564 20816
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 18328 20596 18380 20602
rect 18328 20538 18380 20544
rect 16684 20454 16896 20482
rect 16212 19916 16264 19922
rect 16212 19858 16264 19864
rect 16580 19916 16632 19922
rect 16580 19858 16632 19864
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15474 19272 15530 19281
rect 15474 19207 15530 19216
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15292 19168 15344 19174
rect 15752 19168 15804 19174
rect 15292 19110 15344 19116
rect 15488 19116 15752 19122
rect 15488 19110 15804 19116
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 15212 18834 15240 19110
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 15304 18222 15332 19110
rect 15488 19094 15792 19110
rect 15384 18896 15436 18902
rect 15384 18838 15436 18844
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14844 17270 14872 18022
rect 15304 17882 15332 18158
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 14936 17338 14964 17750
rect 14924 17332 14976 17338
rect 14924 17274 14976 17280
rect 14832 17264 14884 17270
rect 14832 17206 14884 17212
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14280 16176 14332 16182
rect 14280 16118 14332 16124
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 13740 15502 13768 15846
rect 14108 15706 14136 15914
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 14200 15638 14228 15846
rect 14188 15632 14240 15638
rect 14188 15574 14240 15580
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13740 13870 13768 14758
rect 13832 14618 13860 14826
rect 14292 14618 14320 16118
rect 14476 15638 14504 16526
rect 14568 16250 14596 16662
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14660 16114 14688 16526
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14464 15632 14516 15638
rect 14464 15574 14516 15580
rect 14476 15162 14504 15574
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13832 14074 13860 14282
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13636 12436 13688 12442
rect 13832 12434 13860 14010
rect 14568 14006 14596 14418
rect 14556 14000 14608 14006
rect 14556 13942 14608 13948
rect 14660 13190 14688 14826
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 12714 14688 13126
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14844 12434 14872 14214
rect 14936 13462 14964 14758
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 14924 13456 14976 13462
rect 14924 13398 14976 13404
rect 14936 12986 14964 13398
rect 15028 13394 15056 14350
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 15016 12640 15068 12646
rect 15120 12628 15148 13466
rect 15212 13297 15240 16934
rect 15396 15910 15424 18838
rect 15488 18154 15516 19094
rect 15884 19068 16180 19088
rect 15940 19066 15964 19068
rect 16020 19066 16044 19068
rect 16100 19066 16124 19068
rect 15962 19014 15964 19066
rect 16026 19014 16038 19066
rect 16100 19014 16102 19066
rect 15940 19012 15964 19014
rect 16020 19012 16044 19014
rect 16100 19012 16124 19014
rect 15884 18992 16180 19012
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16132 18290 16160 18566
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 15568 18148 15620 18154
rect 15568 18090 15620 18096
rect 15488 17610 15516 18090
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15474 16688 15530 16697
rect 15474 16623 15476 16632
rect 15528 16623 15530 16632
rect 15476 16594 15528 16600
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15198 13288 15254 13297
rect 15198 13223 15254 13232
rect 15068 12600 15148 12628
rect 15016 12582 15068 12588
rect 13832 12406 13952 12434
rect 14844 12406 14964 12434
rect 13636 12378 13688 12384
rect 13648 11626 13676 12378
rect 13924 12170 13952 12406
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 13912 12164 13964 12170
rect 13912 12106 13964 12112
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 12084 10674 12112 11154
rect 12152 10908 12448 10928
rect 12208 10906 12232 10908
rect 12288 10906 12312 10908
rect 12368 10906 12392 10908
rect 12230 10854 12232 10906
rect 12294 10854 12306 10906
rect 12368 10854 12370 10906
rect 12208 10852 12232 10854
rect 12288 10852 12312 10854
rect 12368 10852 12392 10854
rect 12152 10832 12448 10852
rect 12912 10810 12940 11154
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 11244 10532 11296 10538
rect 11244 10474 11296 10480
rect 12084 10266 12112 10610
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 8420 9276 8716 9296
rect 8476 9274 8500 9276
rect 8556 9274 8580 9276
rect 8636 9274 8660 9276
rect 8498 9222 8500 9274
rect 8562 9222 8574 9274
rect 8636 9222 8638 9274
rect 8476 9220 8500 9222
rect 8556 9220 8580 9222
rect 8636 9220 8660 9222
rect 8420 9200 8716 9220
rect 9692 9110 9720 9318
rect 11624 9110 11652 9862
rect 12084 9586 12112 9862
rect 12152 9820 12448 9840
rect 12208 9818 12232 9820
rect 12288 9818 12312 9820
rect 12368 9818 12392 9820
rect 12230 9766 12232 9818
rect 12294 9766 12306 9818
rect 12368 9766 12370 9818
rect 12208 9764 12232 9766
rect 12288 9764 12312 9766
rect 12368 9764 12392 9766
rect 12152 9744 12448 9764
rect 13188 9586 13216 9998
rect 13464 9722 13492 10066
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 11888 9376 11940 9382
rect 12176 9364 12204 9454
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 11940 9336 12204 9364
rect 12716 9376 12768 9382
rect 11888 9318 11940 9324
rect 12716 9318 12768 9324
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 4688 8732 4984 8752
rect 4744 8730 4768 8732
rect 4824 8730 4848 8732
rect 4904 8730 4928 8732
rect 4766 8678 4768 8730
rect 4830 8678 4842 8730
rect 4904 8678 4906 8730
rect 4744 8676 4768 8678
rect 4824 8676 4848 8678
rect 4904 8676 4928 8678
rect 4688 8656 4984 8676
rect 9232 8634 9260 8978
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9692 8430 9720 9046
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 7392 7954 7420 8366
rect 8420 8188 8716 8208
rect 8476 8186 8500 8188
rect 8556 8186 8580 8188
rect 8636 8186 8660 8188
rect 8498 8134 8500 8186
rect 8562 8134 8574 8186
rect 8636 8134 8638 8186
rect 8476 8132 8500 8134
rect 8556 8132 8580 8134
rect 8636 8132 8660 8134
rect 8420 8112 8716 8132
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 4688 7644 4984 7664
rect 4744 7642 4768 7644
rect 4824 7642 4848 7644
rect 4904 7642 4928 7644
rect 4766 7590 4768 7642
rect 4830 7590 4842 7642
rect 4904 7590 4906 7642
rect 4744 7588 4768 7590
rect 4824 7588 4848 7590
rect 4904 7588 4928 7590
rect 4688 7568 4984 7588
rect 9416 7342 9444 8026
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9692 7274 9720 8366
rect 10428 7834 10456 8434
rect 10520 8430 10548 8774
rect 11072 8634 11100 8910
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10520 8022 10548 8366
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10600 7880 10652 7886
rect 10428 7828 10600 7834
rect 10428 7822 10652 7828
rect 10428 7806 10640 7822
rect 10796 7818 10824 8230
rect 11348 8090 11376 8978
rect 11428 8832 11480 8838
rect 11428 8774 11480 8780
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11440 7954 11468 8774
rect 11624 8362 11652 9046
rect 12728 9042 12756 9318
rect 12808 9172 12860 9178
rect 12912 9160 12940 9386
rect 13464 9178 13492 9658
rect 12860 9132 12940 9160
rect 13452 9172 13504 9178
rect 12808 9114 12860 9120
rect 13452 9114 13504 9120
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12152 8732 12448 8752
rect 12208 8730 12232 8732
rect 12288 8730 12312 8732
rect 12368 8730 12392 8732
rect 12230 8678 12232 8730
rect 12294 8678 12306 8730
rect 12368 8678 12370 8730
rect 12208 8676 12232 8678
rect 12288 8676 12312 8678
rect 12368 8676 12392 8678
rect 12152 8656 12448 8676
rect 12544 8514 12572 8978
rect 12820 8922 12848 9114
rect 13556 8974 13584 10066
rect 13832 9586 13860 11018
rect 13924 9926 13952 12106
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14200 11354 14228 11562
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 14004 9580 14056 9586
rect 14004 9522 14056 9528
rect 14016 9450 14044 9522
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 12728 8894 12848 8922
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12452 8486 12572 8514
rect 12452 8362 12480 8486
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12452 8090 12480 8298
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 8420 7100 8716 7120
rect 8476 7098 8500 7100
rect 8556 7098 8580 7100
rect 8636 7098 8660 7100
rect 8498 7046 8500 7098
rect 8562 7046 8574 7098
rect 8636 7046 8638 7098
rect 8476 7044 8500 7046
rect 8556 7044 8580 7046
rect 8636 7044 8660 7046
rect 8420 7024 8716 7044
rect 9692 6866 9720 7210
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 4688 6556 4984 6576
rect 4744 6554 4768 6556
rect 4824 6554 4848 6556
rect 4904 6554 4928 6556
rect 4766 6502 4768 6554
rect 4830 6502 4842 6554
rect 4904 6502 4906 6554
rect 4744 6500 4768 6502
rect 4824 6500 4848 6502
rect 4904 6500 4928 6502
rect 4688 6480 4984 6500
rect 8956 6254 8984 6598
rect 9692 6322 9720 6802
rect 10060 6458 10088 6938
rect 10520 6934 10548 7482
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10612 6798 10640 7806
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 10980 7546 11008 7890
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11900 7313 11928 7686
rect 11992 7546 12020 7890
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 12084 7342 12112 7686
rect 12152 7644 12448 7664
rect 12208 7642 12232 7644
rect 12288 7642 12312 7644
rect 12368 7642 12392 7644
rect 12230 7590 12232 7642
rect 12294 7590 12306 7642
rect 12368 7590 12370 7642
rect 12208 7588 12232 7590
rect 12288 7588 12312 7590
rect 12368 7588 12392 7590
rect 12152 7568 12448 7588
rect 12636 7410 12664 8774
rect 12728 7954 12756 8894
rect 12912 7954 12940 8910
rect 13740 8906 13768 9318
rect 14016 9178 14044 9386
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14108 9110 14136 9930
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14200 9586 14228 9862
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14384 9518 14412 12038
rect 14752 11898 14780 12242
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14844 11830 14872 12174
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14556 11688 14608 11694
rect 14556 11630 14608 11636
rect 14568 11014 14596 11630
rect 14936 11626 14964 12406
rect 15028 12345 15056 12582
rect 15212 12434 15240 13223
rect 15212 12406 15332 12434
rect 15014 12336 15070 12345
rect 15014 12271 15070 12280
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 15028 11150 15056 12174
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15120 11898 15148 12106
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14568 10470 14596 10950
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14568 9722 14596 10406
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14568 9518 14596 9658
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12072 7336 12124 7342
rect 11886 7304 11942 7313
rect 11152 7268 11204 7274
rect 12072 7278 12124 7284
rect 11886 7239 11942 7248
rect 12256 7268 12308 7274
rect 11152 7210 11204 7216
rect 12256 7210 12308 7216
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10784 6792 10836 6798
rect 11060 6792 11112 6798
rect 10836 6740 11008 6746
rect 10784 6734 11008 6740
rect 11060 6734 11112 6740
rect 10796 6718 11008 6734
rect 10980 6662 11008 6718
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8420 6012 8716 6032
rect 8476 6010 8500 6012
rect 8556 6010 8580 6012
rect 8636 6010 8660 6012
rect 8498 5958 8500 6010
rect 8562 5958 8574 6010
rect 8636 5958 8638 6010
rect 8476 5956 8500 5958
rect 8556 5956 8580 5958
rect 8636 5956 8660 5958
rect 8420 5936 8716 5956
rect 9692 5778 9720 6258
rect 10060 5846 10088 6394
rect 11072 6186 11100 6734
rect 11164 6730 11192 7210
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11256 7002 11284 7142
rect 12268 7002 12296 7210
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11532 6458 11560 6802
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12152 6556 12448 6576
rect 12208 6554 12232 6556
rect 12288 6554 12312 6556
rect 12368 6554 12392 6556
rect 12230 6502 12232 6554
rect 12294 6502 12306 6554
rect 12368 6502 12370 6554
rect 12208 6500 12232 6502
rect 12288 6500 12312 6502
rect 12368 6500 12392 6502
rect 12152 6480 12448 6500
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11072 5914 11100 6122
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11532 5846 11560 6394
rect 12544 6186 12572 6734
rect 12636 6458 12664 6802
rect 12912 6798 12940 7890
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13004 7410 13032 7822
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 13004 7002 13032 7142
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12544 5914 12572 6122
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 12636 5846 12664 6394
rect 13096 6254 13124 8366
rect 13280 8090 13308 8570
rect 13556 8430 13584 8774
rect 13740 8498 13768 8842
rect 14108 8634 14136 9046
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 14200 8362 14228 9318
rect 14660 8838 14688 10542
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14188 8356 14240 8362
rect 14188 8298 14240 8304
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13268 8084 13320 8090
rect 13268 8026 13320 8032
rect 13648 7818 13676 8230
rect 14372 8084 14424 8090
rect 14372 8026 14424 8032
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 14016 7546 14044 7890
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14200 7410 14228 7686
rect 14384 7410 14412 8026
rect 14556 7880 14608 7886
rect 14554 7848 14556 7857
rect 14608 7848 14610 7857
rect 14554 7783 14610 7792
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 13096 5846 13124 6190
rect 13372 6186 13400 6802
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 11520 5840 11572 5846
rect 11520 5782 11572 5788
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 4688 5468 4984 5488
rect 4744 5466 4768 5468
rect 4824 5466 4848 5468
rect 4904 5466 4928 5468
rect 4766 5414 4768 5466
rect 4830 5414 4842 5466
rect 4904 5414 4906 5466
rect 4744 5412 4768 5414
rect 4824 5412 4848 5414
rect 4904 5412 4928 5414
rect 4688 5392 4984 5412
rect 12152 5468 12448 5488
rect 12208 5466 12232 5468
rect 12288 5466 12312 5468
rect 12368 5466 12392 5468
rect 12230 5414 12232 5466
rect 12294 5414 12306 5466
rect 12368 5414 12370 5466
rect 12208 5412 12232 5414
rect 12288 5412 12312 5414
rect 12368 5412 12392 5414
rect 12152 5392 12448 5412
rect 13372 5370 13400 6122
rect 13556 5914 13584 6734
rect 13832 6458 13860 7210
rect 14384 6934 14412 7346
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14384 6254 14412 6734
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13556 5166 13584 5850
rect 14568 5778 14596 7142
rect 14660 5778 14688 8774
rect 15028 7886 15056 9318
rect 15212 9042 15240 12242
rect 15304 12102 15332 12406
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 15200 8288 15252 8294
rect 15200 8230 15252 8236
rect 15212 7954 15240 8230
rect 15304 7993 15332 10134
rect 15396 9926 15424 15846
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14618 15516 14894
rect 15580 14822 15608 18090
rect 15884 17980 16180 18000
rect 15940 17978 15964 17980
rect 16020 17978 16044 17980
rect 16100 17978 16124 17980
rect 15962 17926 15964 17978
rect 16026 17926 16038 17978
rect 16100 17926 16102 17978
rect 15940 17924 15964 17926
rect 16020 17924 16044 17926
rect 16100 17924 16124 17926
rect 15884 17904 16180 17924
rect 16224 16998 16252 18702
rect 16592 18698 16620 19110
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16316 17728 16344 18226
rect 16592 17814 16620 18634
rect 16684 18426 16712 20454
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 16868 19922 16896 20266
rect 17972 19990 18000 20538
rect 18340 20330 18368 20538
rect 18328 20324 18380 20330
rect 18328 20266 18380 20272
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17040 19712 17092 19718
rect 17092 19672 17172 19700
rect 17040 19654 17092 19660
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16776 18970 16804 19110
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16960 18630 16988 19110
rect 17144 18766 17172 19672
rect 17420 18834 17448 19858
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17604 19310 17632 19654
rect 18524 19334 18552 20810
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 18432 19306 18552 19334
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16856 18352 16908 18358
rect 16856 18294 16908 18300
rect 16580 17808 16632 17814
rect 16580 17750 16632 17756
rect 16396 17740 16448 17746
rect 16316 17700 16396 17728
rect 16316 17202 16344 17700
rect 16396 17682 16448 17688
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 15884 16892 16180 16912
rect 15940 16890 15964 16892
rect 16020 16890 16044 16892
rect 16100 16890 16124 16892
rect 15962 16838 15964 16890
rect 16026 16838 16038 16890
rect 16100 16838 16102 16890
rect 15940 16836 15964 16838
rect 16020 16836 16044 16838
rect 16100 16836 16124 16838
rect 15884 16816 16180 16836
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15672 16046 15700 16594
rect 15752 16108 15804 16114
rect 15752 16050 15804 16056
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15488 12306 15516 13942
rect 15672 12434 15700 15642
rect 15764 15162 15792 16050
rect 15884 15804 16180 15824
rect 15940 15802 15964 15804
rect 16020 15802 16044 15804
rect 16100 15802 16124 15804
rect 15962 15750 15964 15802
rect 16026 15750 16038 15802
rect 16100 15750 16102 15802
rect 15940 15748 15964 15750
rect 16020 15748 16044 15750
rect 16100 15748 16124 15750
rect 15884 15728 16180 15748
rect 16120 15632 16172 15638
rect 16120 15574 16172 15580
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 16132 15094 16160 15574
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 16224 15026 16252 16730
rect 16316 16658 16344 17138
rect 16304 16652 16356 16658
rect 16356 16612 16436 16640
rect 16304 16594 16356 16600
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16316 15638 16344 16390
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16408 15570 16436 16612
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16396 15088 16448 15094
rect 16396 15030 16448 15036
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 15884 14716 16180 14736
rect 15940 14714 15964 14716
rect 16020 14714 16044 14716
rect 16100 14714 16124 14716
rect 15962 14662 15964 14714
rect 16026 14662 16038 14714
rect 16100 14662 16102 14714
rect 15940 14660 15964 14662
rect 16020 14660 16044 14662
rect 16100 14660 16124 14662
rect 15884 14640 16180 14660
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15764 13190 15792 14418
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 15884 13628 16180 13648
rect 15940 13626 15964 13628
rect 16020 13626 16044 13628
rect 16100 13626 16124 13628
rect 15962 13574 15964 13626
rect 16026 13574 16038 13626
rect 16100 13574 16102 13626
rect 15940 13572 15964 13574
rect 16020 13572 16044 13574
rect 16100 13572 16124 13574
rect 15884 13552 16180 13572
rect 16224 13512 16252 14350
rect 16040 13484 16252 13512
rect 16040 13394 16068 13484
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 16040 12986 16068 13330
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16316 12782 16344 14758
rect 16408 14006 16436 15030
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16500 13870 16528 17206
rect 16868 17134 16896 18294
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16580 14544 16632 14550
rect 16580 14486 16632 14492
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16396 13184 16448 13190
rect 16448 13144 16528 13172
rect 16396 13126 16448 13132
rect 16500 12850 16528 13144
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 15936 12776 15988 12782
rect 15934 12744 15936 12753
rect 16304 12776 16356 12782
rect 15988 12744 15990 12753
rect 16304 12718 16356 12724
rect 15934 12679 15990 12688
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15764 12442 15792 12582
rect 15884 12540 16180 12560
rect 15940 12538 15964 12540
rect 16020 12538 16044 12540
rect 16100 12538 16124 12540
rect 15962 12486 15964 12538
rect 16026 12486 16038 12538
rect 16100 12486 16102 12538
rect 15940 12484 15964 12486
rect 16020 12484 16044 12486
rect 16100 12484 16124 12486
rect 15884 12464 16180 12484
rect 15580 12406 15700 12434
rect 15752 12436 15804 12442
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15476 9988 15528 9994
rect 15476 9930 15528 9936
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15290 7984 15346 7993
rect 15200 7948 15252 7954
rect 15290 7919 15292 7928
rect 15200 7890 15252 7896
rect 15344 7919 15346 7928
rect 15292 7890 15344 7896
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14752 5642 14780 6122
rect 15212 5914 15240 7142
rect 15304 6662 15332 7142
rect 15396 6866 15424 7346
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15396 6458 15424 6802
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15488 6254 15516 9930
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 14740 5636 14792 5642
rect 14740 5578 14792 5584
rect 14752 5234 14780 5578
rect 15396 5234 15424 5714
rect 15488 5574 15516 6190
rect 15580 5846 15608 12406
rect 15752 12378 15804 12384
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 11286 15700 12242
rect 16132 11898 16160 12310
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16040 11676 16068 11834
rect 16304 11688 16356 11694
rect 16040 11648 16304 11676
rect 16304 11630 16356 11636
rect 15884 11452 16180 11472
rect 15940 11450 15964 11452
rect 16020 11450 16044 11452
rect 16100 11450 16124 11452
rect 15962 11398 15964 11450
rect 16026 11398 16038 11450
rect 16100 11398 16102 11450
rect 15940 11396 15964 11398
rect 16020 11396 16044 11398
rect 16100 11396 16124 11398
rect 15884 11376 16180 11396
rect 15660 11280 15712 11286
rect 16408 11268 16436 12174
rect 16592 12170 16620 14486
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16670 14376 16726 14385
rect 16670 14311 16726 14320
rect 16684 13938 16712 14311
rect 16776 14278 16804 14418
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16776 12782 16804 14214
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16868 12628 16896 17070
rect 16960 16726 16988 18566
rect 17144 18222 17172 18702
rect 17132 18216 17184 18222
rect 17420 18170 17448 18770
rect 17604 18290 17632 19246
rect 18236 18896 18288 18902
rect 18236 18838 18288 18844
rect 18248 18426 18276 18838
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 18340 18306 18368 18566
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 18248 18278 18368 18306
rect 17132 18158 17184 18164
rect 17328 18142 17448 18170
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17236 17814 17264 18022
rect 17224 17808 17276 17814
rect 17224 17750 17276 17756
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 17144 16046 17172 16934
rect 17328 16250 17356 18142
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17420 17746 17448 18022
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17420 16454 17448 17682
rect 17696 17678 17724 18226
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17512 16726 17540 17478
rect 17604 17134 17632 17478
rect 17696 17338 17724 17614
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17696 17134 17724 17274
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17604 16266 17632 17070
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17420 16238 17632 16266
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17224 15904 17276 15910
rect 17224 15846 17276 15852
rect 17236 14958 17264 15846
rect 17224 14952 17276 14958
rect 17420 14929 17448 16238
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17592 16040 17644 16046
rect 17696 16028 17724 17070
rect 17776 17060 17828 17066
rect 17776 17002 17828 17008
rect 17788 16794 17816 17002
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17644 16000 17724 16028
rect 17868 16040 17920 16046
rect 17592 15982 17644 15988
rect 17868 15982 17920 15988
rect 17512 15570 17540 15982
rect 17604 15910 17632 15982
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17500 15564 17552 15570
rect 17500 15506 17552 15512
rect 17604 15502 17632 15846
rect 17880 15706 17908 15982
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17774 15056 17830 15065
rect 17774 14991 17776 15000
rect 17828 14991 17830 15000
rect 17776 14962 17828 14968
rect 17224 14894 17276 14900
rect 17406 14920 17462 14929
rect 17406 14855 17462 14864
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17420 13938 17448 14214
rect 17512 13938 17540 14826
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 16948 13728 17000 13734
rect 16948 13670 17000 13676
rect 16684 12600 16896 12628
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16488 11688 16540 11694
rect 16540 11648 16620 11676
rect 16488 11630 16540 11636
rect 15660 11222 15712 11228
rect 16316 11240 16436 11268
rect 15672 10810 15700 11222
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 16316 10538 16344 11240
rect 16488 11212 16540 11218
rect 16408 11172 16488 11200
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 16304 10532 16356 10538
rect 16304 10474 16356 10480
rect 15764 10266 15792 10474
rect 15884 10364 16180 10384
rect 15940 10362 15964 10364
rect 16020 10362 16044 10364
rect 16100 10362 16124 10364
rect 15962 10310 15964 10362
rect 16026 10310 16038 10362
rect 16100 10310 16102 10362
rect 15940 10308 15964 10310
rect 16020 10308 16044 10310
rect 16100 10308 16124 10310
rect 15884 10288 16180 10308
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15672 8294 15700 9862
rect 16316 9722 16344 10474
rect 16408 10266 16436 11172
rect 16488 11154 16540 11160
rect 16592 11014 16620 11648
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16592 10470 16620 10950
rect 16684 10674 16712 12600
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16776 11694 16804 12038
rect 16960 11694 16988 13670
rect 17144 13258 17172 13806
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17328 13530 17356 13670
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17420 13394 17448 13874
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17512 13326 17540 13670
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17144 12850 17172 13194
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17130 12744 17186 12753
rect 17040 12708 17092 12714
rect 17130 12679 17186 12688
rect 17040 12650 17092 12656
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16580 10464 16632 10470
rect 16486 10432 16542 10441
rect 16580 10406 16632 10412
rect 16486 10367 16542 10376
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16500 9654 16528 10367
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 15884 9276 16180 9296
rect 15940 9274 15964 9276
rect 16020 9274 16044 9276
rect 16100 9274 16124 9276
rect 15962 9222 15964 9274
rect 16026 9222 16038 9274
rect 16100 9222 16102 9274
rect 15940 9220 15964 9222
rect 16020 9220 16044 9222
rect 16100 9220 16124 9222
rect 15884 9200 16180 9220
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15764 8430 15792 8978
rect 16316 8838 16344 9454
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15672 5914 15700 7142
rect 15764 6798 15792 8366
rect 15884 8188 16180 8208
rect 15940 8186 15964 8188
rect 16020 8186 16044 8188
rect 16100 8186 16124 8188
rect 15962 8134 15964 8186
rect 16026 8134 16038 8186
rect 16100 8134 16102 8186
rect 15940 8132 15964 8134
rect 16020 8132 16044 8134
rect 16100 8132 16124 8134
rect 15884 8112 16180 8132
rect 15842 7440 15898 7449
rect 15842 7375 15844 7384
rect 15896 7375 15898 7384
rect 15844 7346 15896 7352
rect 15884 7100 16180 7120
rect 15940 7098 15964 7100
rect 16020 7098 16044 7100
rect 16100 7098 16124 7100
rect 15962 7046 15964 7098
rect 16026 7046 16038 7098
rect 16100 7046 16102 7098
rect 15940 7044 15964 7046
rect 16020 7044 16044 7046
rect 16100 7044 16124 7046
rect 15884 7024 16180 7044
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15764 5710 15792 6598
rect 15884 6012 16180 6032
rect 15940 6010 15964 6012
rect 16020 6010 16044 6012
rect 16100 6010 16124 6012
rect 15962 5958 15964 6010
rect 16026 5958 16038 6010
rect 16100 5958 16102 6010
rect 15940 5956 15964 5958
rect 16020 5956 16044 5958
rect 16100 5956 16124 5958
rect 15884 5936 16180 5956
rect 16028 5772 16080 5778
rect 16224 5760 16252 6598
rect 16080 5732 16252 5760
rect 16028 5714 16080 5720
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 16316 5166 16344 8774
rect 16592 8566 16620 8774
rect 16684 8566 16712 8774
rect 16580 8560 16632 8566
rect 16580 8502 16632 8508
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16488 7880 16540 7886
rect 16486 7848 16488 7857
rect 16540 7848 16542 7857
rect 16486 7783 16542 7792
rect 16776 7206 16804 11494
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16868 10198 16896 11290
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16856 9648 16908 9654
rect 16854 9616 16856 9625
rect 16908 9616 16910 9625
rect 16854 9551 16910 9560
rect 17052 9518 17080 12650
rect 17144 12374 17172 12679
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 17222 12336 17278 12345
rect 17328 12322 17356 13194
rect 17512 12782 17540 13262
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17328 12294 17448 12322
rect 17222 12271 17278 12280
rect 17236 12238 17264 12271
rect 17420 12238 17448 12294
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 17144 11762 17172 12106
rect 17224 11892 17276 11898
rect 17224 11834 17276 11840
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17236 11558 17264 11834
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17420 11150 17448 12174
rect 17512 11665 17540 12718
rect 17604 12714 17632 14554
rect 17788 13870 17816 14962
rect 17972 14618 18000 18158
rect 18248 18086 18276 18278
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18052 16720 18104 16726
rect 18050 16688 18052 16697
rect 18104 16688 18106 16697
rect 18050 16623 18106 16632
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18064 14793 18092 14894
rect 18050 14784 18106 14793
rect 18050 14719 18106 14728
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17498 11656 17554 11665
rect 17498 11591 17554 11600
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17512 10810 17540 11591
rect 17604 11354 17632 12242
rect 17696 11762 17724 12582
rect 17788 12238 17816 12922
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17788 11694 17816 12038
rect 17880 11898 17908 14350
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17972 11830 18000 12106
rect 18064 11898 18092 14418
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 18064 11286 18092 11834
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17144 9908 17172 10542
rect 18064 10538 18092 11086
rect 17224 10532 17276 10538
rect 17224 10474 17276 10480
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 17236 10062 17264 10474
rect 17500 10464 17552 10470
rect 18064 10441 18092 10474
rect 17500 10406 17552 10412
rect 18050 10432 18106 10441
rect 17406 10160 17462 10169
rect 17406 10095 17408 10104
rect 17460 10095 17462 10104
rect 17408 10066 17460 10072
rect 17224 10056 17276 10062
rect 17276 10004 17356 10010
rect 17224 9998 17356 10004
rect 17236 9982 17356 9998
rect 17224 9920 17276 9926
rect 17144 9880 17224 9908
rect 17224 9862 17276 9868
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 17328 9450 17356 9982
rect 17512 9450 17540 10406
rect 18050 10367 18106 10376
rect 18156 9450 18184 15098
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17500 9444 17552 9450
rect 17500 9386 17552 9392
rect 17592 9444 17644 9450
rect 17592 9386 17644 9392
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16960 9042 16988 9318
rect 17512 9178 17540 9386
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 17604 8566 17632 9386
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 17592 8560 17644 8566
rect 17592 8502 17644 8508
rect 16856 8288 16908 8294
rect 16856 8230 16908 8236
rect 16868 8090 16896 8230
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16960 7750 16988 8502
rect 17972 8498 18000 9046
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8634 18092 8774
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18248 8498 18276 18022
rect 18432 15162 18460 19306
rect 18708 18034 18736 21490
rect 18800 21146 18828 21966
rect 18984 21894 19012 23800
rect 19628 22098 19656 23800
rect 20168 22160 20220 22166
rect 20168 22102 20220 22108
rect 19064 22092 19116 22098
rect 19064 22034 19116 22040
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19616 22092 19668 22098
rect 19616 22034 19668 22040
rect 20076 22092 20128 22098
rect 20076 22034 20128 22040
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18880 21344 18932 21350
rect 18880 21286 18932 21292
rect 18788 21140 18840 21146
rect 18788 21082 18840 21088
rect 18892 21010 18920 21286
rect 19076 21146 19104 22034
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19154 21584 19210 21593
rect 19260 21554 19288 21966
rect 19154 21519 19210 21528
rect 19248 21548 19300 21554
rect 19168 21418 19196 21519
rect 19248 21490 19300 21496
rect 19156 21412 19208 21418
rect 19156 21354 19208 21360
rect 19168 21146 19196 21354
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18892 20466 18920 20946
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 18984 20466 19012 20742
rect 19260 20602 19288 21490
rect 19352 20602 19380 22034
rect 19444 21078 19472 22034
rect 19616 21788 19912 21808
rect 19672 21786 19696 21788
rect 19752 21786 19776 21788
rect 19832 21786 19856 21788
rect 19694 21734 19696 21786
rect 19758 21734 19770 21786
rect 19832 21734 19834 21786
rect 19672 21732 19696 21734
rect 19752 21732 19776 21734
rect 19832 21732 19856 21734
rect 19616 21712 19912 21732
rect 20088 21622 20116 22034
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 20180 21486 20208 22102
rect 20272 22098 20300 23800
rect 20916 22098 20944 23800
rect 20260 22092 20312 22098
rect 20260 22034 20312 22040
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20904 22092 20956 22098
rect 20904 22034 20956 22040
rect 21088 22092 21140 22098
rect 21088 22034 21140 22040
rect 21456 22092 21508 22098
rect 21456 22034 21508 22040
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 19432 21072 19484 21078
rect 19432 21014 19484 21020
rect 20444 21004 20496 21010
rect 20444 20946 20496 20952
rect 19616 20700 19912 20720
rect 19672 20698 19696 20700
rect 19752 20698 19776 20700
rect 19832 20698 19856 20700
rect 19694 20646 19696 20698
rect 19758 20646 19770 20698
rect 19832 20646 19834 20698
rect 19672 20644 19696 20646
rect 19752 20644 19776 20646
rect 19832 20644 19856 20646
rect 19616 20624 19912 20644
rect 19248 20596 19300 20602
rect 19248 20538 19300 20544
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18972 20460 19024 20466
rect 18972 20402 19024 20408
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18800 20074 18828 20334
rect 18984 20262 19012 20402
rect 18972 20256 19024 20262
rect 18972 20198 19024 20204
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 18800 20046 19012 20074
rect 19076 20058 19104 20198
rect 18984 19854 19012 20046
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18984 19310 19012 19790
rect 19260 19417 19288 19994
rect 19246 19408 19302 19417
rect 19246 19343 19302 19352
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19168 18766 19196 19246
rect 19156 18760 19208 18766
rect 19156 18702 19208 18708
rect 19168 18154 19196 18702
rect 19260 18698 19288 19343
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 18616 18006 18736 18034
rect 18512 15972 18564 15978
rect 18512 15914 18564 15920
rect 18420 15156 18472 15162
rect 18340 15116 18420 15144
rect 18340 13920 18368 15116
rect 18420 15098 18472 15104
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18432 14521 18460 14758
rect 18418 14512 18474 14521
rect 18418 14447 18474 14456
rect 18340 13892 18460 13920
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18340 13530 18368 13738
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18328 13388 18380 13394
rect 18328 13330 18380 13336
rect 18340 13297 18368 13330
rect 18326 13288 18382 13297
rect 18326 13223 18382 13232
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18340 8838 18368 9998
rect 18432 9674 18460 13892
rect 18524 12306 18552 15914
rect 18616 14074 18644 18006
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18512 12300 18564 12306
rect 18512 12242 18564 12248
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 10062 18552 10406
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18432 9646 18552 9674
rect 18616 9654 18644 13466
rect 18708 13462 18736 17818
rect 19064 17740 19116 17746
rect 19064 17682 19116 17688
rect 19076 17338 19104 17682
rect 19352 17678 19380 19110
rect 19444 18222 19472 19110
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19536 18034 19564 20198
rect 20088 19990 20116 20198
rect 20076 19984 20128 19990
rect 20076 19926 20128 19932
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19616 19612 19912 19632
rect 19672 19610 19696 19612
rect 19752 19610 19776 19612
rect 19832 19610 19856 19612
rect 19694 19558 19696 19610
rect 19758 19558 19770 19610
rect 19832 19558 19834 19610
rect 19672 19556 19696 19558
rect 19752 19556 19776 19558
rect 19832 19556 19856 19558
rect 19616 19536 19912 19556
rect 19616 18524 19912 18544
rect 19672 18522 19696 18524
rect 19752 18522 19776 18524
rect 19832 18522 19856 18524
rect 19694 18470 19696 18522
rect 19758 18470 19770 18522
rect 19832 18470 19834 18522
rect 19672 18468 19696 18470
rect 19752 18468 19776 18470
rect 19832 18468 19856 18470
rect 19616 18448 19912 18468
rect 19708 18216 19760 18222
rect 19708 18158 19760 18164
rect 19444 18006 19564 18034
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 19352 17270 19380 17478
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 18880 16652 18932 16658
rect 18880 16594 18932 16600
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18892 16250 18920 16594
rect 18972 16584 19024 16590
rect 18972 16526 19024 16532
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18880 15904 18932 15910
rect 18984 15892 19012 16526
rect 18932 15864 19012 15892
rect 18880 15846 18932 15852
rect 18892 15502 18920 15846
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18880 15360 18932 15366
rect 18800 15320 18880 15348
rect 18696 13456 18748 13462
rect 18696 13398 18748 13404
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18708 11286 18736 13262
rect 18696 11280 18748 11286
rect 18696 11222 18748 11228
rect 18696 10464 18748 10470
rect 18694 10432 18696 10441
rect 18748 10432 18750 10441
rect 18694 10367 18750 10376
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18432 9382 18460 9522
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18328 8832 18380 8838
rect 18328 8774 18380 8780
rect 18340 8566 18368 8774
rect 18328 8560 18380 8566
rect 18328 8502 18380 8508
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17314 7984 17370 7993
rect 17224 7948 17276 7954
rect 17314 7919 17316 7928
rect 17224 7890 17276 7896
rect 17368 7919 17370 7928
rect 17316 7890 17368 7896
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 17236 7410 17264 7890
rect 17604 7886 17632 8298
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7546 17632 7822
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 17144 6730 17172 7346
rect 17406 7304 17462 7313
rect 17406 7239 17462 7248
rect 17420 7206 17448 7239
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16960 6254 16988 6598
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16960 5234 16988 6190
rect 17144 6186 17172 6666
rect 17328 6458 17356 7142
rect 17604 6866 17632 7346
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17972 6458 18000 8434
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 18156 7857 18184 8366
rect 18340 8090 18368 8502
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18142 7848 18198 7857
rect 18142 7783 18144 7792
rect 18196 7783 18198 7792
rect 18144 7754 18196 7760
rect 18156 7723 18184 7754
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 18236 6180 18288 6186
rect 18236 6122 18288 6128
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 8420 4924 8716 4944
rect 8476 4922 8500 4924
rect 8556 4922 8580 4924
rect 8636 4922 8660 4924
rect 8498 4870 8500 4922
rect 8562 4870 8574 4922
rect 8636 4870 8638 4922
rect 8476 4868 8500 4870
rect 8556 4868 8580 4870
rect 8636 4868 8660 4870
rect 8420 4848 8716 4868
rect 15884 4924 16180 4944
rect 15940 4922 15964 4924
rect 16020 4922 16044 4924
rect 16100 4922 16124 4924
rect 15962 4870 15964 4922
rect 16026 4870 16038 4922
rect 16100 4870 16102 4922
rect 15940 4868 15964 4870
rect 16020 4868 16044 4870
rect 16100 4868 16124 4870
rect 15884 4848 16180 4868
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 4688 4380 4984 4400
rect 4744 4378 4768 4380
rect 4824 4378 4848 4380
rect 4904 4378 4928 4380
rect 4766 4326 4768 4378
rect 4830 4326 4842 4378
rect 4904 4326 4906 4378
rect 4744 4324 4768 4326
rect 4824 4324 4848 4326
rect 4904 4324 4928 4326
rect 4688 4304 4984 4324
rect 12152 4380 12448 4400
rect 12208 4378 12232 4380
rect 12288 4378 12312 4380
rect 12368 4378 12392 4380
rect 12230 4326 12232 4378
rect 12294 4326 12306 4378
rect 12368 4326 12370 4378
rect 12208 4324 12232 4326
rect 12288 4324 12312 4326
rect 12368 4324 12392 4326
rect 12152 4304 12448 4324
rect 16132 4282 16160 4626
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16684 4078 16712 4422
rect 16960 4146 16988 5170
rect 17236 5166 17264 5850
rect 18052 5840 18104 5846
rect 18052 5782 18104 5788
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17684 5704 17736 5710
rect 17684 5646 17736 5652
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17696 4826 17724 5646
rect 17880 5370 17908 5714
rect 17960 5636 18012 5642
rect 17960 5578 18012 5584
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17880 4758 17908 5306
rect 17972 5030 18000 5578
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17868 4752 17920 4758
rect 17868 4694 17920 4700
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17236 4078 17264 4626
rect 18064 4622 18092 5782
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 5234 18184 5510
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 17776 4616 17828 4622
rect 17776 4558 17828 4564
rect 18052 4616 18104 4622
rect 18052 4558 18104 4564
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17788 4010 17816 4558
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 8420 3836 8716 3856
rect 8476 3834 8500 3836
rect 8556 3834 8580 3836
rect 8636 3834 8660 3836
rect 8498 3782 8500 3834
rect 8562 3782 8574 3834
rect 8636 3782 8638 3834
rect 8476 3780 8500 3782
rect 8556 3780 8580 3782
rect 8636 3780 8660 3782
rect 8420 3760 8716 3780
rect 15884 3836 16180 3856
rect 15940 3834 15964 3836
rect 16020 3834 16044 3836
rect 16100 3834 16124 3836
rect 15962 3782 15964 3834
rect 16026 3782 16038 3834
rect 16100 3782 16102 3834
rect 15940 3780 15964 3782
rect 16020 3780 16044 3782
rect 16100 3780 16124 3782
rect 15884 3760 16180 3780
rect 4068 3664 4120 3670
rect 4068 3606 4120 3612
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3712 3194 3740 3334
rect 4688 3292 4984 3312
rect 4744 3290 4768 3292
rect 4824 3290 4848 3292
rect 4904 3290 4928 3292
rect 4766 3238 4768 3290
rect 4830 3238 4842 3290
rect 4904 3238 4906 3290
rect 4744 3236 4768 3238
rect 4824 3236 4848 3238
rect 4904 3236 4928 3238
rect 4688 3216 4984 3236
rect 12152 3292 12448 3312
rect 12208 3290 12232 3292
rect 12288 3290 12312 3292
rect 12368 3290 12392 3292
rect 12230 3238 12232 3290
rect 12294 3238 12306 3290
rect 12368 3238 12370 3290
rect 12208 3236 12232 3238
rect 12288 3236 12312 3238
rect 12368 3236 12392 3238
rect 12152 3216 12448 3236
rect 16500 3194 16528 3878
rect 17788 3602 17816 3946
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 1400 3120 1452 3126
rect 1398 3088 1400 3097
rect 1452 3088 1454 3097
rect 1398 3023 1454 3032
rect 3712 2922 3740 3130
rect 17236 2990 17264 3334
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 3700 2916 3752 2922
rect 3700 2858 3752 2864
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2516 2582 2544 2790
rect 6104 2582 6132 2926
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 8420 2748 8716 2768
rect 8476 2746 8500 2748
rect 8556 2746 8580 2748
rect 8636 2746 8660 2748
rect 8498 2694 8500 2746
rect 8562 2694 8574 2746
rect 8636 2694 8638 2746
rect 8476 2692 8500 2694
rect 8556 2692 8580 2694
rect 8636 2692 8660 2694
rect 8420 2672 8716 2692
rect 10704 2650 10732 2790
rect 15884 2748 16180 2768
rect 15940 2746 15964 2748
rect 16020 2746 16044 2748
rect 16100 2746 16124 2748
rect 15962 2694 15964 2746
rect 16026 2694 16038 2746
rect 16100 2694 16102 2746
rect 15940 2692 15964 2694
rect 16020 2692 16044 2694
rect 16100 2692 16124 2694
rect 15884 2672 16180 2692
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 2504 2576 2556 2582
rect 2504 2518 2556 2524
rect 6092 2576 6144 2582
rect 6092 2518 6144 2524
rect 16960 2514 16988 2926
rect 17788 2514 17816 3538
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 17972 2854 18000 3062
rect 18248 2922 18276 6122
rect 18524 5914 18552 9646
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18708 9466 18736 10367
rect 18800 10266 18828 15320
rect 18880 15302 18932 15308
rect 18984 14906 19012 15642
rect 19076 15570 19104 16594
rect 19260 15609 19288 16934
rect 19444 16726 19472 18006
rect 19720 17882 19748 18158
rect 19708 17876 19760 17882
rect 19708 17818 19760 17824
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19536 16969 19564 17750
rect 19616 17436 19912 17456
rect 19672 17434 19696 17436
rect 19752 17434 19776 17436
rect 19832 17434 19856 17436
rect 19694 17382 19696 17434
rect 19758 17382 19770 17434
rect 19832 17382 19834 17434
rect 19672 17380 19696 17382
rect 19752 17380 19776 17382
rect 19832 17380 19856 17382
rect 19616 17360 19912 17380
rect 19996 17338 20024 19858
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 20088 19514 20116 19790
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20076 18964 20128 18970
rect 20076 18906 20128 18912
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19522 16960 19578 16969
rect 19522 16895 19578 16904
rect 19628 16810 19656 17138
rect 19892 16992 19944 16998
rect 19892 16934 19944 16940
rect 19536 16782 19656 16810
rect 19904 16794 19932 16934
rect 19800 16788 19852 16794
rect 19432 16720 19484 16726
rect 19432 16662 19484 16668
rect 19432 16584 19484 16590
rect 19430 16552 19432 16561
rect 19484 16552 19486 16561
rect 19340 16516 19392 16522
rect 19430 16487 19486 16496
rect 19340 16458 19392 16464
rect 19352 16046 19380 16458
rect 19536 16114 19564 16782
rect 19800 16730 19852 16736
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19812 16697 19840 16730
rect 19798 16688 19854 16697
rect 19798 16623 19854 16632
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19616 16348 19912 16368
rect 19672 16346 19696 16348
rect 19752 16346 19776 16348
rect 19832 16346 19856 16348
rect 19694 16294 19696 16346
rect 19758 16294 19770 16346
rect 19832 16294 19834 16346
rect 19672 16292 19696 16294
rect 19752 16292 19776 16294
rect 19832 16292 19856 16294
rect 19616 16272 19912 16292
rect 19996 16250 20024 16594
rect 19984 16244 20036 16250
rect 20088 16232 20116 18906
rect 20180 18222 20208 19654
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 20088 16204 20208 16232
rect 19984 16186 20036 16192
rect 19616 16176 19668 16182
rect 19800 16176 19852 16182
rect 19668 16124 19800 16130
rect 19616 16118 19852 16124
rect 19524 16108 19576 16114
rect 19628 16102 19840 16118
rect 20076 16108 20128 16114
rect 19524 16050 19576 16056
rect 20076 16050 20128 16056
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 20088 15910 20116 16050
rect 19800 15904 19852 15910
rect 19800 15846 19852 15852
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19812 15706 19840 15846
rect 19800 15700 19852 15706
rect 19800 15642 19852 15648
rect 19246 15600 19302 15609
rect 19064 15564 19116 15570
rect 19246 15535 19302 15544
rect 19984 15564 20036 15570
rect 19064 15506 19116 15512
rect 19984 15506 20036 15512
rect 18975 14878 19012 14906
rect 18880 14816 18932 14822
rect 18878 14784 18880 14793
rect 18932 14784 18934 14793
rect 18975 14770 19003 14878
rect 18975 14742 19012 14770
rect 18878 14719 18934 14728
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18892 12782 18920 13126
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18984 11506 19012 14742
rect 19076 12345 19104 15506
rect 19340 15496 19392 15502
rect 19392 15456 19564 15484
rect 19340 15438 19392 15444
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 19168 14385 19196 15098
rect 19536 15076 19564 15456
rect 19616 15260 19912 15280
rect 19672 15258 19696 15260
rect 19752 15258 19776 15260
rect 19832 15258 19856 15260
rect 19694 15206 19696 15258
rect 19758 15206 19770 15258
rect 19832 15206 19834 15258
rect 19672 15204 19696 15206
rect 19752 15204 19776 15206
rect 19832 15204 19856 15206
rect 19616 15184 19912 15204
rect 19536 15048 19656 15076
rect 19248 14884 19300 14890
rect 19248 14826 19300 14832
rect 19154 14376 19210 14385
rect 19260 14346 19288 14826
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19154 14311 19210 14320
rect 19248 14340 19300 14346
rect 19248 14282 19300 14288
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19168 13938 19196 14214
rect 19260 14074 19288 14282
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19248 13864 19300 13870
rect 19248 13806 19300 13812
rect 19260 12918 19288 13806
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 19062 12336 19118 12345
rect 19062 12271 19118 12280
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19076 11626 19104 12174
rect 19168 11694 19196 12582
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19064 11620 19116 11626
rect 19064 11562 19116 11568
rect 18984 11478 19104 11506
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18616 9438 18736 9466
rect 18616 8294 18644 9438
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18708 8498 18736 9318
rect 18800 8634 18828 9522
rect 18892 9160 18920 10406
rect 18984 9625 19012 10542
rect 19076 9654 19104 11478
rect 19156 11280 19208 11286
rect 19156 11222 19208 11228
rect 19168 10606 19196 11222
rect 19260 11218 19288 12582
rect 19352 11626 19380 14554
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19444 14006 19472 14418
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19536 13852 19564 14758
rect 19628 14385 19656 15048
rect 19890 15056 19946 15065
rect 19996 15042 20024 15506
rect 19946 15014 20024 15042
rect 19890 14991 19946 15000
rect 19904 14958 19932 14991
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 19892 14816 19944 14822
rect 19812 14776 19892 14804
rect 19812 14414 19840 14776
rect 19892 14758 19944 14764
rect 19996 14618 20024 14826
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 19800 14408 19852 14414
rect 19614 14376 19670 14385
rect 19800 14350 19852 14356
rect 19614 14311 19670 14320
rect 19616 14172 19912 14192
rect 19672 14170 19696 14172
rect 19752 14170 19776 14172
rect 19832 14170 19856 14172
rect 19694 14118 19696 14170
rect 19758 14118 19770 14170
rect 19832 14118 19834 14170
rect 19672 14116 19696 14118
rect 19752 14116 19776 14118
rect 19832 14116 19856 14118
rect 19616 14096 19912 14116
rect 19444 13824 19564 13852
rect 19444 12889 19472 13824
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19430 12880 19486 12889
rect 19536 12850 19564 13126
rect 19616 13084 19912 13104
rect 19672 13082 19696 13084
rect 19752 13082 19776 13084
rect 19832 13082 19856 13084
rect 19694 13030 19696 13082
rect 19758 13030 19770 13082
rect 19832 13030 19834 13082
rect 19672 13028 19696 13030
rect 19752 13028 19776 13030
rect 19832 13028 19856 13030
rect 19616 13008 19912 13028
rect 19430 12815 19486 12824
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19444 12442 19472 12650
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19628 12442 19656 12582
rect 19996 12442 20024 14418
rect 20180 14090 20208 16204
rect 20272 15745 20300 20198
rect 20352 19236 20404 19242
rect 20352 19178 20404 19184
rect 20364 18630 20392 19178
rect 20456 18970 20484 20946
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20640 19718 20668 19858
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 17134 20392 18566
rect 20456 18086 20484 18770
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20456 17202 20484 18022
rect 20548 17202 20576 19246
rect 20640 18329 20668 19654
rect 20626 18320 20682 18329
rect 20626 18255 20682 18264
rect 20732 17882 20760 19722
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20732 17202 20760 17818
rect 20824 17320 20852 22034
rect 21100 21350 21128 22034
rect 21088 21344 21140 21350
rect 21088 21286 21140 21292
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21376 21010 21404 21286
rect 21468 21146 21496 22034
rect 21560 22030 21588 23800
rect 21836 22273 21864 24239
rect 22190 23800 22246 24600
rect 22834 23800 22890 24600
rect 23478 23800 23534 24600
rect 24122 23800 24178 24600
rect 22098 23624 22154 23633
rect 22098 23559 22154 23568
rect 22006 22944 22062 22953
rect 22006 22879 22062 22888
rect 21822 22264 21878 22273
rect 21822 22199 21878 22208
rect 21638 22128 21694 22137
rect 21638 22063 21640 22072
rect 21692 22063 21694 22072
rect 21824 22092 21876 22098
rect 21640 22034 21692 22040
rect 21824 22034 21876 22040
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21456 21140 21508 21146
rect 21456 21082 21508 21088
rect 21560 21026 21588 21286
rect 21180 21004 21232 21010
rect 21364 21004 21416 21010
rect 21180 20946 21232 20952
rect 21284 20964 21364 20992
rect 21192 20874 21220 20946
rect 21180 20868 21232 20874
rect 21180 20810 21232 20816
rect 20904 20392 20956 20398
rect 20904 20334 20956 20340
rect 20916 20262 20944 20334
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 20916 18873 20944 20198
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20902 18864 20958 18873
rect 20902 18799 20958 18808
rect 21008 18766 21036 19790
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 21008 18154 21036 18702
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 21008 17678 21036 18090
rect 21100 17898 21128 19858
rect 21192 19242 21220 20198
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21100 17870 21220 17898
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21100 17338 21128 17682
rect 21088 17332 21140 17338
rect 20824 17292 21036 17320
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20444 17060 20496 17066
rect 20444 17002 20496 17008
rect 20456 16114 20484 17002
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20258 15736 20314 15745
rect 20258 15671 20314 15680
rect 20260 15632 20312 15638
rect 20260 15574 20312 15580
rect 20272 14618 20300 15574
rect 20456 14822 20484 16050
rect 20548 15638 20576 16594
rect 20732 16590 20760 17138
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20916 16250 20944 16526
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20732 15638 20760 15982
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20720 15632 20772 15638
rect 20720 15574 20772 15580
rect 20628 15360 20680 15366
rect 20548 15308 20628 15314
rect 20548 15302 20680 15308
rect 20548 15286 20668 15302
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20180 14062 20484 14090
rect 20260 14000 20312 14006
rect 20260 13942 20312 13948
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19432 11688 19484 11694
rect 19430 11656 19432 11665
rect 19484 11656 19486 11665
rect 19340 11620 19392 11626
rect 19430 11591 19486 11600
rect 19340 11562 19392 11568
rect 19430 11248 19486 11257
rect 19248 11212 19300 11218
rect 19430 11183 19486 11192
rect 19248 11154 19300 11160
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19352 10713 19380 11086
rect 19444 10810 19472 11183
rect 19432 10804 19484 10810
rect 19536 10792 19564 12038
rect 19616 11996 19912 12016
rect 19672 11994 19696 11996
rect 19752 11994 19776 11996
rect 19832 11994 19856 11996
rect 19694 11942 19696 11994
rect 19758 11942 19770 11994
rect 19832 11942 19834 11994
rect 19672 11940 19696 11942
rect 19752 11940 19776 11942
rect 19832 11940 19856 11942
rect 19616 11920 19912 11940
rect 19996 11558 20024 12038
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19996 11150 20024 11494
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19616 10908 19912 10928
rect 19672 10906 19696 10908
rect 19752 10906 19776 10908
rect 19832 10906 19856 10908
rect 19694 10854 19696 10906
rect 19758 10854 19770 10906
rect 19832 10854 19834 10906
rect 19672 10852 19696 10854
rect 19752 10852 19776 10854
rect 19832 10852 19856 10854
rect 19616 10832 19912 10852
rect 19996 10792 20024 10950
rect 19536 10764 19656 10792
rect 19432 10746 19484 10752
rect 19628 10713 19656 10764
rect 19720 10764 20024 10792
rect 19338 10704 19394 10713
rect 19614 10704 19670 10713
rect 19338 10639 19394 10648
rect 19432 10668 19484 10674
rect 19484 10628 19564 10656
rect 19614 10639 19670 10648
rect 19432 10610 19484 10616
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19430 10568 19486 10577
rect 19168 10169 19196 10542
rect 19430 10503 19486 10512
rect 19340 10464 19392 10470
rect 19444 10452 19472 10503
rect 19392 10424 19472 10452
rect 19340 10406 19392 10412
rect 19338 10296 19394 10305
rect 19338 10231 19394 10240
rect 19154 10160 19210 10169
rect 19154 10095 19210 10104
rect 19064 9648 19116 9654
rect 18970 9616 19026 9625
rect 19064 9590 19116 9596
rect 18970 9551 19026 9560
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 18892 9132 19012 9160
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18616 7750 18644 8230
rect 18892 7886 18920 8978
rect 18880 7880 18932 7886
rect 18800 7840 18880 7868
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 18800 7546 18828 7840
rect 18880 7822 18932 7828
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18984 7426 19012 9132
rect 19076 8090 19104 9318
rect 19168 8514 19196 10095
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9625 19288 9862
rect 19352 9722 19380 10231
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19246 9616 19302 9625
rect 19444 9586 19472 10134
rect 19536 10044 19564 10628
rect 19720 10554 19748 10764
rect 19798 10704 19854 10713
rect 19798 10639 19800 10648
rect 19852 10639 19854 10648
rect 19800 10610 19852 10616
rect 19628 10526 19748 10554
rect 19628 10198 19656 10526
rect 19708 10464 19760 10470
rect 19706 10432 19708 10441
rect 19812 10452 19840 10610
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19892 10464 19944 10470
rect 19760 10432 19762 10441
rect 19812 10424 19892 10452
rect 19892 10406 19944 10412
rect 19706 10367 19762 10376
rect 19996 10266 20024 10542
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19616 10192 19668 10198
rect 19616 10134 19668 10140
rect 19616 10056 19668 10062
rect 19536 10016 19616 10044
rect 19246 9551 19302 9560
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19352 9110 19380 9386
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19168 8486 19288 8514
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19168 7954 19196 8366
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19260 7818 19288 8486
rect 19248 7812 19300 7818
rect 19248 7754 19300 7760
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 18892 7398 19012 7426
rect 18788 6860 18840 6866
rect 18788 6802 18840 6808
rect 18800 6186 18828 6802
rect 18892 6390 18920 7398
rect 19168 6934 19196 7686
rect 19246 7440 19302 7449
rect 19246 7375 19302 7384
rect 19156 6928 19208 6934
rect 19156 6870 19208 6876
rect 19168 6458 19196 6870
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 18880 6384 18932 6390
rect 18880 6326 18932 6332
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18524 5574 18552 5850
rect 18892 5710 18920 6326
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18984 5914 19012 6054
rect 18972 5908 19024 5914
rect 18972 5850 19024 5856
rect 19168 5778 19196 6258
rect 19156 5772 19208 5778
rect 19156 5714 19208 5720
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18788 5160 18840 5166
rect 18788 5102 18840 5108
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18616 4826 18644 4966
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18696 4684 18748 4690
rect 18696 4626 18748 4632
rect 18340 4214 18368 4626
rect 18328 4208 18380 4214
rect 18328 4150 18380 4156
rect 18340 3670 18368 4150
rect 18708 4010 18736 4626
rect 18800 4282 18828 5102
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18696 4004 18748 4010
rect 18696 3946 18748 3952
rect 18708 3738 18736 3946
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18236 2916 18288 2922
rect 18236 2858 18288 2864
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18340 2582 18368 2790
rect 18524 2650 18552 3538
rect 19076 3058 19104 4490
rect 19168 3602 19196 4558
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19260 2922 19288 7375
rect 19352 7154 19380 9046
rect 19444 8090 19472 9318
rect 19536 8906 19564 10016
rect 19616 9998 19668 10004
rect 19616 9820 19912 9840
rect 19672 9818 19696 9820
rect 19752 9818 19776 9820
rect 19832 9818 19856 9820
rect 19694 9766 19696 9818
rect 19758 9766 19770 9818
rect 19832 9766 19834 9818
rect 19672 9764 19696 9766
rect 19752 9764 19776 9766
rect 19832 9764 19856 9766
rect 19616 9744 19912 9764
rect 19996 9586 20024 10202
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 20088 9518 20116 13874
rect 20166 13832 20222 13841
rect 20166 13767 20168 13776
rect 20220 13767 20222 13776
rect 20168 13738 20220 13744
rect 20166 13560 20222 13569
rect 20166 13495 20222 13504
rect 20180 12986 20208 13495
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20180 11286 20208 11630
rect 20168 11280 20220 11286
rect 20168 11222 20220 11228
rect 20166 11112 20222 11121
rect 20166 11047 20222 11056
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 20088 9178 20116 9454
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19892 8900 19944 8906
rect 19944 8860 20024 8888
rect 19892 8842 19944 8848
rect 19616 8732 19912 8752
rect 19672 8730 19696 8732
rect 19752 8730 19776 8732
rect 19832 8730 19856 8732
rect 19694 8678 19696 8730
rect 19758 8678 19770 8730
rect 19832 8678 19834 8730
rect 19672 8676 19696 8678
rect 19752 8676 19776 8678
rect 19832 8676 19856 8678
rect 19616 8656 19912 8676
rect 19996 8430 20024 8860
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19708 7880 19760 7886
rect 19706 7848 19708 7857
rect 19760 7848 19762 7857
rect 19706 7783 19762 7792
rect 19616 7644 19912 7664
rect 19672 7642 19696 7644
rect 19752 7642 19776 7644
rect 19832 7642 19856 7644
rect 19694 7590 19696 7642
rect 19758 7590 19770 7642
rect 19832 7590 19834 7642
rect 19672 7588 19696 7590
rect 19752 7588 19776 7590
rect 19832 7588 19856 7590
rect 19616 7568 19912 7588
rect 19996 7342 20024 8366
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 20088 7750 20116 7822
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 20180 7449 20208 11047
rect 20272 10985 20300 13942
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20258 10976 20314 10985
rect 20258 10911 20314 10920
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20272 9110 20300 9318
rect 20260 9104 20312 9110
rect 20260 9046 20312 9052
rect 20364 8945 20392 13806
rect 20456 13802 20484 14062
rect 20444 13796 20496 13802
rect 20444 13738 20496 13744
rect 20456 13297 20484 13738
rect 20442 13288 20498 13297
rect 20442 13223 20498 13232
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20456 12102 20484 13126
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20456 11762 20484 11834
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20548 11665 20576 15286
rect 20732 15178 20760 15574
rect 20732 15162 20852 15178
rect 20628 15156 20680 15162
rect 20732 15156 20864 15162
rect 20732 15150 20812 15156
rect 20628 15098 20680 15104
rect 20812 15098 20864 15104
rect 20640 12102 20668 15098
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20732 14618 20760 14894
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 13870 20944 14214
rect 20720 13864 20772 13870
rect 20904 13864 20956 13870
rect 20720 13806 20772 13812
rect 20810 13832 20866 13841
rect 20732 12918 20760 13806
rect 20904 13806 20956 13812
rect 20810 13767 20866 13776
rect 20824 13394 20852 13767
rect 20902 13424 20958 13433
rect 20812 13388 20864 13394
rect 20902 13359 20958 13368
rect 20812 13330 20864 13336
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20720 12912 20772 12918
rect 20720 12854 20772 12860
rect 20732 12306 20760 12854
rect 20720 12300 20772 12306
rect 20720 12242 20772 12248
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20534 11656 20590 11665
rect 20534 11591 20590 11600
rect 20640 11286 20668 12038
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20442 11112 20498 11121
rect 20442 11047 20498 11056
rect 20350 8936 20406 8945
rect 20260 8900 20312 8906
rect 20350 8871 20406 8880
rect 20260 8842 20312 8848
rect 20166 7440 20222 7449
rect 20166 7375 20222 7384
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19616 7268 19668 7274
rect 19536 7228 19616 7256
rect 19352 7126 19472 7154
rect 19338 7032 19394 7041
rect 19338 6967 19394 6976
rect 19352 6866 19380 6967
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19444 6746 19472 7126
rect 19352 6718 19472 6746
rect 19352 3398 19380 6718
rect 19432 6248 19484 6254
rect 19536 6236 19564 7228
rect 19616 7210 19668 7216
rect 20076 7268 20128 7274
rect 20076 7210 20128 7216
rect 20088 6905 20116 7210
rect 20074 6896 20130 6905
rect 20074 6831 20130 6840
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19616 6556 19912 6576
rect 19672 6554 19696 6556
rect 19752 6554 19776 6556
rect 19832 6554 19856 6556
rect 19694 6502 19696 6554
rect 19758 6502 19770 6554
rect 19832 6502 19834 6554
rect 19672 6500 19696 6502
rect 19752 6500 19776 6502
rect 19832 6500 19856 6502
rect 19616 6480 19912 6500
rect 19996 6361 20024 6666
rect 19982 6352 20038 6361
rect 19982 6287 20038 6296
rect 19484 6208 19564 6236
rect 19432 6190 19484 6196
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19536 4622 19564 5646
rect 19616 5468 19912 5488
rect 19672 5466 19696 5468
rect 19752 5466 19776 5468
rect 19832 5466 19856 5468
rect 19694 5414 19696 5466
rect 19758 5414 19770 5466
rect 19832 5414 19834 5466
rect 19672 5412 19696 5414
rect 19752 5412 19776 5414
rect 19832 5412 19856 5414
rect 19616 5392 19912 5412
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 20166 4992 20222 5001
rect 19524 4616 19576 4622
rect 19524 4558 19576 4564
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19352 3194 19380 3334
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19444 3058 19472 4082
rect 19536 4078 19564 4558
rect 19616 4380 19912 4400
rect 19672 4378 19696 4380
rect 19752 4378 19776 4380
rect 19832 4378 19856 4380
rect 19694 4326 19696 4378
rect 19758 4326 19770 4378
rect 19832 4326 19834 4378
rect 19672 4324 19696 4326
rect 19752 4324 19776 4326
rect 19832 4324 19856 4326
rect 19616 4304 19912 4324
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19536 3602 19564 4014
rect 19892 3664 19944 3670
rect 19890 3632 19892 3641
rect 19944 3632 19946 3641
rect 19524 3596 19576 3602
rect 19890 3567 19946 3576
rect 19524 3538 19576 3544
rect 19616 3292 19912 3312
rect 19672 3290 19696 3292
rect 19752 3290 19776 3292
rect 19832 3290 19856 3292
rect 19694 3238 19696 3290
rect 19758 3238 19770 3290
rect 19832 3238 19834 3290
rect 19672 3236 19696 3238
rect 19752 3236 19776 3238
rect 19832 3236 19856 3238
rect 19616 3216 19912 3236
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 19260 2774 19288 2858
rect 19168 2746 19288 2774
rect 19168 2650 19196 2746
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 19996 2514 20024 4966
rect 20166 4927 20222 4936
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 20088 3942 20116 4694
rect 20180 4146 20208 4927
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20088 2854 20116 3878
rect 20272 3754 20300 8842
rect 20456 7970 20484 11047
rect 20548 10044 20576 11154
rect 20628 10056 20680 10062
rect 20548 10016 20628 10044
rect 20628 9998 20680 10004
rect 20640 9518 20668 9998
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20640 8974 20668 9454
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20364 7942 20484 7970
rect 20364 6882 20392 7942
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20456 7750 20484 7822
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20548 7546 20576 8774
rect 20640 8430 20668 8910
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20628 8288 20680 8294
rect 20628 8230 20680 8236
rect 20640 7886 20668 8230
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20732 7392 20760 11834
rect 20824 10130 20852 13126
rect 20916 11762 20944 13359
rect 21008 11898 21036 17292
rect 21088 17274 21140 17280
rect 21192 15570 21220 17870
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21180 14476 21232 14482
rect 21180 14418 21232 14424
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21100 13326 21128 14350
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21192 13172 21220 14418
rect 21100 13144 21220 13172
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20904 11756 20956 11762
rect 20904 11698 20956 11704
rect 20916 10470 20944 11698
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20916 9926 20944 10066
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20916 9042 20944 9862
rect 21008 9450 21036 10950
rect 20996 9444 21048 9450
rect 20996 9386 21048 9392
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20812 7880 20864 7886
rect 20810 7848 20812 7857
rect 20864 7848 20866 7857
rect 20810 7783 20866 7792
rect 20916 7562 20944 8298
rect 20916 7546 21036 7562
rect 20916 7540 21048 7546
rect 20916 7534 20996 7540
rect 20996 7482 21048 7488
rect 20732 7364 20852 7392
rect 20442 7304 20498 7313
rect 20442 7239 20444 7248
rect 20496 7239 20498 7248
rect 20720 7268 20772 7274
rect 20444 7210 20496 7216
rect 20720 7210 20772 7216
rect 20628 6928 20680 6934
rect 20364 6854 20576 6882
rect 20628 6870 20680 6876
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 20364 5914 20392 6734
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20456 6458 20484 6666
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20364 4078 20392 5510
rect 20548 4434 20576 6854
rect 20640 6730 20668 6870
rect 20628 6724 20680 6730
rect 20628 6666 20680 6672
rect 20732 6390 20760 7210
rect 20824 6798 20852 7364
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20824 6390 20852 6598
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20812 6384 20864 6390
rect 20812 6326 20864 6332
rect 20720 6180 20772 6186
rect 20720 6122 20772 6128
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20640 4554 20668 6054
rect 20732 5642 20760 6122
rect 20916 6118 20944 6938
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20824 5930 20852 6054
rect 21008 5930 21036 7142
rect 20824 5902 21036 5930
rect 21100 5846 21128 13144
rect 21178 12744 21234 12753
rect 21178 12679 21234 12688
rect 21192 11257 21220 12679
rect 21178 11248 21234 11257
rect 21178 11183 21234 11192
rect 21284 9874 21312 20964
rect 21364 20946 21416 20952
rect 21468 20998 21588 21026
rect 21468 20058 21496 20998
rect 21652 20602 21680 21422
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21744 20754 21772 20946
rect 21836 20874 21864 22034
rect 21928 20874 21956 22034
rect 22020 22030 22048 22879
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 22112 21894 22140 23559
rect 22204 21962 22232 23800
rect 22284 22228 22336 22234
rect 22284 22170 22336 22176
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22296 21434 22324 22170
rect 22848 21690 22876 23800
rect 23110 22264 23166 22273
rect 23110 22199 23166 22208
rect 23124 22098 23152 22199
rect 23112 22092 23164 22098
rect 23112 22034 23164 22040
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 23492 21622 23520 23800
rect 23480 21616 23532 21622
rect 23110 21584 23166 21593
rect 23480 21558 23532 21564
rect 23110 21519 23112 21528
rect 23164 21519 23166 21528
rect 23112 21490 23164 21496
rect 22112 21406 22324 21434
rect 22112 21146 22140 21406
rect 22192 21344 22244 21350
rect 22192 21286 22244 21292
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 22008 21072 22060 21078
rect 22008 21014 22060 21020
rect 21824 20868 21876 20874
rect 21824 20810 21876 20816
rect 21916 20868 21968 20874
rect 21916 20810 21968 20816
rect 21744 20726 21864 20754
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 21548 20528 21600 20534
rect 21548 20470 21600 20476
rect 21560 20346 21588 20470
rect 21640 20392 21692 20398
rect 21560 20340 21640 20346
rect 21560 20334 21692 20340
rect 21560 20318 21680 20334
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21376 18902 21404 19110
rect 21364 18896 21416 18902
rect 21364 18838 21416 18844
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21376 17134 21404 18090
rect 21456 17740 21508 17746
rect 21456 17682 21508 17688
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21468 16658 21496 17682
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21468 16046 21496 16390
rect 21456 16040 21508 16046
rect 21456 15982 21508 15988
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21376 13841 21404 14758
rect 21468 14521 21496 15302
rect 21454 14512 21510 14521
rect 21454 14447 21510 14456
rect 21362 13832 21418 13841
rect 21468 13802 21496 14447
rect 21362 13767 21418 13776
rect 21456 13796 21508 13802
rect 21456 13738 21508 13744
rect 21364 12708 21416 12714
rect 21468 12696 21496 13738
rect 21416 12668 21496 12696
rect 21364 12650 21416 12656
rect 21468 12374 21496 12668
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21192 9846 21312 9874
rect 21192 8906 21220 9846
rect 21376 9674 21404 12038
rect 21456 11280 21508 11286
rect 21456 11222 21508 11228
rect 21468 10674 21496 11222
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21468 10266 21496 10610
rect 21456 10260 21508 10266
rect 21456 10202 21508 10208
rect 21376 9646 21496 9674
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21272 8288 21324 8294
rect 21178 8256 21234 8265
rect 21272 8230 21324 8236
rect 21178 8191 21234 8200
rect 21192 6798 21220 8191
rect 21284 7886 21312 8230
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 21088 5840 21140 5846
rect 21088 5782 21140 5788
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20456 4406 20576 4434
rect 20456 4214 20484 4406
rect 20534 4312 20590 4321
rect 20534 4247 20590 4256
rect 20444 4208 20496 4214
rect 20444 4150 20496 4156
rect 20548 4146 20576 4247
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20352 4072 20404 4078
rect 20352 4014 20404 4020
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20272 3738 20392 3754
rect 20272 3732 20404 3738
rect 20272 3726 20352 3732
rect 20352 3674 20404 3680
rect 20260 3664 20312 3670
rect 20260 3606 20312 3612
rect 20168 3188 20220 3194
rect 20272 3176 20300 3606
rect 20640 3602 20668 4014
rect 20732 3738 20760 4966
rect 20824 3942 20852 5102
rect 21008 4622 21036 5170
rect 21088 5024 21140 5030
rect 21088 4966 21140 4972
rect 20996 4616 21048 4622
rect 20996 4558 21048 4564
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20220 3148 20300 3176
rect 20444 3188 20496 3194
rect 20168 3130 20220 3136
rect 20444 3130 20496 3136
rect 20258 3088 20314 3097
rect 20258 3023 20314 3032
rect 20272 2990 20300 3023
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20456 2922 20484 3130
rect 20824 2990 20852 3538
rect 20812 2984 20864 2990
rect 20534 2952 20590 2961
rect 20444 2916 20496 2922
rect 20812 2926 20864 2932
rect 20534 2887 20590 2896
rect 20444 2858 20496 2864
rect 20076 2848 20128 2854
rect 20076 2790 20128 2796
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20364 2378 20392 2450
rect 20548 2446 20576 2887
rect 20720 2508 20772 2514
rect 20824 2496 20852 2926
rect 20916 2514 20944 3674
rect 21008 2990 21036 4422
rect 21100 3670 21128 4966
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21088 3664 21140 3670
rect 21088 3606 21140 3612
rect 21192 3194 21220 3878
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 20772 2468 20852 2496
rect 20904 2508 20956 2514
rect 20720 2450 20772 2456
rect 20904 2450 20956 2456
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 6092 2372 6144 2378
rect 6092 2314 6144 2320
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 18420 2372 18472 2378
rect 18420 2314 18472 2320
rect 20352 2372 20404 2378
rect 20352 2314 20404 2320
rect 2056 800 2084 2314
rect 4688 2204 4984 2224
rect 4744 2202 4768 2204
rect 4824 2202 4848 2204
rect 4904 2202 4928 2204
rect 4766 2150 4768 2202
rect 4830 2150 4842 2202
rect 4904 2150 4906 2202
rect 4744 2148 4768 2150
rect 4824 2148 4848 2150
rect 4904 2148 4928 2150
rect 4688 2128 4984 2148
rect 6104 800 6132 2314
rect 10244 800 10272 2314
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 12152 2204 12448 2224
rect 12208 2202 12232 2204
rect 12288 2202 12312 2204
rect 12368 2202 12392 2204
rect 12230 2150 12232 2202
rect 12294 2150 12306 2202
rect 12368 2150 12370 2202
rect 12208 2148 12232 2150
rect 12288 2148 12312 2150
rect 12368 2148 12392 2150
rect 12152 2128 12448 2148
rect 14292 800 14320 2246
rect 18432 800 18460 2314
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19444 2106 19472 2246
rect 19616 2204 19912 2224
rect 19672 2202 19696 2204
rect 19752 2202 19776 2204
rect 19832 2202 19856 2204
rect 19694 2150 19696 2202
rect 19758 2150 19770 2202
rect 19832 2150 19834 2202
rect 19672 2148 19696 2150
rect 19752 2148 19776 2150
rect 19832 2148 19856 2150
rect 19616 2128 19912 2148
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 20364 2038 20392 2314
rect 21284 2310 21312 6054
rect 21362 5672 21418 5681
rect 21468 5658 21496 9646
rect 21560 9382 21588 20318
rect 21640 19372 21692 19378
rect 21640 19314 21692 19320
rect 21652 14482 21680 19314
rect 21732 19304 21784 19310
rect 21732 19246 21784 19252
rect 21744 18902 21772 19246
rect 21732 18896 21784 18902
rect 21732 18838 21784 18844
rect 21836 17218 21864 20726
rect 22020 20602 22048 21014
rect 22100 21004 22152 21010
rect 22204 20992 22232 21286
rect 24136 21146 24164 23800
rect 24124 21140 24176 21146
rect 24124 21082 24176 21088
rect 22152 20964 22232 20992
rect 22284 21004 22336 21010
rect 22100 20946 22152 20952
rect 22284 20946 22336 20952
rect 22112 20874 22140 20946
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 22192 20392 22244 20398
rect 22192 20334 22244 20340
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 21916 19304 21968 19310
rect 21968 19264 22048 19292
rect 21916 19246 21968 19252
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21744 17190 21864 17218
rect 21640 14476 21692 14482
rect 21640 14418 21692 14424
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 21652 12782 21680 13670
rect 21640 12776 21692 12782
rect 21640 12718 21692 12724
rect 21744 12102 21772 17190
rect 21824 17128 21876 17134
rect 21824 17070 21876 17076
rect 21836 16250 21864 17070
rect 21928 17066 21956 19110
rect 22020 18086 22048 19264
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 21916 17060 21968 17066
rect 21916 17002 21968 17008
rect 22020 16726 22048 18022
rect 22112 17746 22140 20198
rect 22100 17740 22152 17746
rect 22100 17682 22152 17688
rect 22204 17338 22232 20334
rect 22296 19514 22324 20946
rect 23480 20936 23532 20942
rect 22742 20904 22798 20913
rect 23480 20878 23532 20884
rect 22742 20839 22744 20848
rect 22796 20839 22798 20848
rect 22744 20810 22796 20816
rect 23020 20800 23072 20806
rect 23020 20742 23072 20748
rect 22836 20324 22888 20330
rect 22836 20266 22888 20272
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22388 19310 22416 19858
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22376 19304 22428 19310
rect 22376 19246 22428 19252
rect 22388 18970 22416 19246
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 22008 16720 22060 16726
rect 21914 16688 21970 16697
rect 22008 16662 22060 16668
rect 21914 16623 21970 16632
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21824 13796 21876 13802
rect 21824 13738 21876 13744
rect 21836 13190 21864 13738
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 21928 13002 21956 16623
rect 22112 14958 22140 17206
rect 22480 17202 22508 18362
rect 22572 18086 22600 19654
rect 22848 19378 22876 20266
rect 23032 20233 23060 20742
rect 23018 20224 23074 20233
rect 23018 20159 23074 20168
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 23112 19780 23164 19786
rect 23112 19722 23164 19728
rect 23124 19553 23152 19722
rect 23110 19544 23166 19553
rect 23110 19479 23166 19488
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22848 18290 22876 19314
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 23032 18902 23060 19110
rect 23020 18896 23072 18902
rect 23020 18838 23072 18844
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22560 18080 22612 18086
rect 22560 18022 22612 18028
rect 22572 17814 22600 18022
rect 22560 17808 22612 17814
rect 22560 17750 22612 17756
rect 22664 17610 22692 18158
rect 22652 17604 22704 17610
rect 22652 17546 22704 17552
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22468 17196 22520 17202
rect 22468 17138 22520 17144
rect 22572 17134 22600 17478
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22192 16992 22244 16998
rect 22192 16934 22244 16940
rect 22204 16046 22232 16934
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 22192 16040 22244 16046
rect 22192 15982 22244 15988
rect 22204 15094 22232 15982
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 22296 15026 22324 15574
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22388 14618 22416 16050
rect 22756 15978 22784 17138
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22744 15972 22796 15978
rect 22744 15914 22796 15920
rect 22756 15706 22784 15914
rect 22744 15700 22796 15706
rect 22744 15642 22796 15648
rect 22848 15638 22876 16390
rect 22836 15632 22888 15638
rect 22836 15574 22888 15580
rect 22560 15360 22612 15366
rect 22560 15302 22612 15308
rect 22468 14816 22520 14822
rect 22468 14758 22520 14764
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22100 14544 22152 14550
rect 22100 14486 22152 14492
rect 22112 13954 22140 14486
rect 22204 14074 22232 14554
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22284 14000 22336 14006
rect 22112 13926 22232 13954
rect 22284 13942 22336 13948
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 21836 12974 21956 13002
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21836 11914 21864 12974
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21928 12374 21956 12786
rect 21916 12368 21968 12374
rect 21916 12310 21968 12316
rect 21744 11886 21864 11914
rect 22020 11898 22048 13330
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22008 11892 22060 11898
rect 21744 9674 21772 11886
rect 22008 11834 22060 11840
rect 21916 11008 21968 11014
rect 21916 10950 21968 10956
rect 21928 10577 21956 10950
rect 21914 10568 21970 10577
rect 21914 10503 21970 10512
rect 21824 9920 21876 9926
rect 21876 9880 21956 9908
rect 21824 9862 21876 9868
rect 21652 9654 21772 9674
rect 21640 9648 21772 9654
rect 21692 9646 21772 9648
rect 21928 9674 21956 9880
rect 21928 9646 22048 9674
rect 21640 9590 21692 9596
rect 21640 9444 21692 9450
rect 21640 9386 21692 9392
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21560 7206 21588 8570
rect 21652 7750 21680 9386
rect 21815 9036 21867 9042
rect 21744 8996 21815 9024
rect 21744 8634 21772 8996
rect 21815 8978 21867 8984
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21732 8016 21784 8022
rect 21732 7958 21784 7964
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21744 7546 21772 7958
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 21732 7540 21784 7546
rect 21732 7482 21784 7488
rect 21640 7472 21692 7478
rect 21640 7414 21692 7420
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 21652 6934 21680 7414
rect 21836 7290 21864 7890
rect 21744 7262 21864 7290
rect 21744 7002 21772 7262
rect 21732 6996 21784 7002
rect 21732 6938 21784 6944
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21560 5914 21588 6802
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21652 5778 21680 6598
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21916 6180 21968 6186
rect 22020 6168 22048 9646
rect 22112 9518 22140 12786
rect 22204 11898 22232 13926
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22112 8294 22140 9318
rect 22204 9178 22232 10610
rect 22192 9172 22244 9178
rect 22192 9114 22244 9120
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 22100 7336 22152 7342
rect 22098 7304 22100 7313
rect 22152 7304 22154 7313
rect 22098 7239 22154 7248
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 21968 6140 22048 6168
rect 21916 6122 21968 6128
rect 21640 5772 21692 5778
rect 21640 5714 21692 5720
rect 21468 5630 21680 5658
rect 21362 5607 21418 5616
rect 21376 4758 21404 5607
rect 21456 5568 21508 5574
rect 21456 5510 21508 5516
rect 21364 4752 21416 4758
rect 21364 4694 21416 4700
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21376 4282 21404 4558
rect 21364 4276 21416 4282
rect 21364 4218 21416 4224
rect 21376 3097 21404 4218
rect 21362 3088 21418 3097
rect 21362 3023 21364 3032
rect 21416 3023 21418 3032
rect 21364 2994 21416 3000
rect 21468 2514 21496 5510
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21560 4554 21588 5170
rect 21548 4548 21600 4554
rect 21548 4490 21600 4496
rect 21560 4010 21588 4490
rect 21652 4078 21680 5630
rect 21744 5030 21772 6122
rect 22204 5574 22232 7210
rect 22296 6254 22324 13942
rect 22480 13802 22508 14758
rect 22572 14482 22600 15302
rect 22940 15026 22968 16390
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 22650 14512 22706 14521
rect 22560 14476 22612 14482
rect 22650 14447 22652 14456
rect 22560 14418 22612 14424
rect 22704 14447 22706 14456
rect 22652 14418 22704 14424
rect 22572 13938 22600 14418
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22468 13796 22520 13802
rect 22468 13738 22520 13744
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22388 12753 22416 13330
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22374 12744 22430 12753
rect 22374 12679 22430 12688
rect 22376 12640 22428 12646
rect 22376 12582 22428 12588
rect 22388 10810 22416 12582
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22480 10674 22508 13262
rect 22560 12980 22612 12986
rect 22560 12922 22612 12928
rect 22572 11694 22600 12922
rect 22652 12708 22704 12714
rect 22652 12650 22704 12656
rect 22664 12186 22692 12650
rect 22756 12306 22784 14214
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22848 12306 22876 13262
rect 22744 12300 22796 12306
rect 22744 12242 22796 12248
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 22664 12158 22784 12186
rect 22560 11688 22612 11694
rect 22560 11630 22612 11636
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22664 11354 22692 11494
rect 22652 11348 22704 11354
rect 22652 11290 22704 11296
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22468 10532 22520 10538
rect 22468 10474 22520 10480
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22388 9722 22416 10406
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22480 9178 22508 10474
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22480 8838 22508 9114
rect 22572 9042 22600 11086
rect 22756 11014 22784 12158
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22652 10532 22704 10538
rect 22652 10474 22704 10480
rect 22560 9036 22612 9042
rect 22560 8978 22612 8984
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22376 8424 22428 8430
rect 22376 8366 22428 8372
rect 22388 7886 22416 8366
rect 22468 8288 22520 8294
rect 22468 8230 22520 8236
rect 22560 8288 22612 8294
rect 22560 8230 22612 8236
rect 22480 7954 22508 8230
rect 22572 8090 22600 8230
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22572 7546 22600 8026
rect 22664 7818 22692 10474
rect 22836 10056 22888 10062
rect 22836 9998 22888 10004
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22756 8634 22784 9522
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22388 5302 22416 7346
rect 22848 6746 22876 9998
rect 22928 7880 22980 7886
rect 23032 7834 23060 18838
rect 23112 16652 23164 16658
rect 23112 16594 23164 16600
rect 23124 16250 23152 16594
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23216 10742 23244 19858
rect 23492 12918 23520 20878
rect 23572 19372 23624 19378
rect 23572 19314 23624 19320
rect 23584 17649 23612 19314
rect 23570 17640 23626 17649
rect 23570 17575 23626 17584
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23204 10736 23256 10742
rect 23204 10678 23256 10684
rect 22980 7828 23060 7834
rect 22928 7822 23060 7828
rect 22756 6718 22876 6746
rect 22940 7806 23060 7822
rect 22756 6662 22784 6718
rect 22744 6656 22796 6662
rect 22744 6598 22796 6604
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22468 5840 22520 5846
rect 22468 5782 22520 5788
rect 22376 5296 22428 5302
rect 22376 5238 22428 5244
rect 22192 5160 22244 5166
rect 22192 5102 22244 5108
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 21640 4072 21692 4078
rect 21640 4014 21692 4020
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 21744 3602 21772 3878
rect 22112 3602 22140 4966
rect 22204 4282 22232 5102
rect 22192 4276 22244 4282
rect 22192 4218 22244 4224
rect 22296 4146 22324 5102
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 22388 4758 22416 5034
rect 22480 5030 22508 5782
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22376 4752 22428 4758
rect 22376 4694 22428 4700
rect 22480 4214 22508 4966
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22468 4208 22520 4214
rect 22468 4150 22520 4156
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22572 4078 22600 4626
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22572 3738 22600 4014
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 21732 3596 21784 3602
rect 21732 3538 21784 3544
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 21744 2310 21772 3538
rect 22008 2916 22060 2922
rect 22008 2858 22060 2864
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 21732 2304 21784 2310
rect 21928 2281 21956 2790
rect 22020 2582 22048 2858
rect 22664 2650 22692 6394
rect 22744 6180 22796 6186
rect 22744 6122 22796 6128
rect 22756 5234 22784 6122
rect 22848 5778 22876 6598
rect 22836 5772 22888 5778
rect 22836 5714 22888 5720
rect 22744 5228 22796 5234
rect 22744 5170 22796 5176
rect 22848 4690 22876 5714
rect 22836 4684 22888 4690
rect 22756 4644 22836 4672
rect 22756 3670 22784 4644
rect 22836 4626 22888 4632
rect 22744 3664 22796 3670
rect 22744 3606 22796 3612
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 2990 22876 3334
rect 22836 2984 22888 2990
rect 22836 2926 22888 2932
rect 22940 2774 22968 7806
rect 23112 6384 23164 6390
rect 23112 6326 23164 6332
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 23032 3738 23060 6054
rect 23124 4690 23152 6326
rect 23112 4684 23164 4690
rect 23112 4626 23164 4632
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 22848 2746 22968 2774
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22008 2576 22060 2582
rect 22008 2518 22060 2524
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 21732 2246 21784 2252
rect 21914 2272 21970 2281
rect 21914 2207 21970 2216
rect 20352 2032 20404 2038
rect 20352 1974 20404 1980
rect 22020 921 22048 2382
rect 22204 2106 22232 2450
rect 22192 2100 22244 2106
rect 22192 2042 22244 2048
rect 22006 912 22062 921
rect 22006 847 22062 856
rect 22480 800 22508 2586
rect 22848 2446 22876 2746
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 23032 1601 23060 2790
rect 23216 2582 23244 10678
rect 23296 10124 23348 10130
rect 23296 10066 23348 10072
rect 23308 9382 23336 10066
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23296 9376 23348 9382
rect 23296 9318 23348 9324
rect 23308 7585 23336 9318
rect 23294 7576 23350 7585
rect 23294 7511 23350 7520
rect 23308 7041 23336 7511
rect 23294 7032 23350 7041
rect 23294 6967 23350 6976
rect 23308 3942 23336 6967
rect 23400 5098 23428 9590
rect 23388 5092 23440 5098
rect 23388 5034 23440 5040
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 23204 2576 23256 2582
rect 23204 2518 23256 2524
rect 23492 2038 23520 12854
rect 23480 2032 23532 2038
rect 23480 1974 23532 1980
rect 23018 1592 23074 1601
rect 23018 1527 23074 1536
rect 23572 1420 23624 1426
rect 23572 1362 23624 1368
rect 2042 0 2098 800
rect 6090 0 6146 800
rect 10230 0 10286 800
rect 14278 0 14334 800
rect 18418 0 18474 800
rect 22466 0 22522 800
rect 23584 377 23612 1362
rect 23570 368 23626 377
rect 23570 303 23626 312
<< via2 >>
rect 21822 24248 21878 24304
rect 1582 21428 1584 21448
rect 1584 21428 1636 21448
rect 1636 21428 1638 21448
rect 1582 21392 1638 21428
rect 2502 21564 2504 21584
rect 2504 21564 2556 21584
rect 2556 21564 2558 21584
rect 2502 21528 2558 21564
rect 3698 21936 3754 21992
rect 1674 20868 1730 20904
rect 1674 20848 1676 20868
rect 1676 20848 1728 20868
rect 1728 20848 1730 20868
rect 4688 21786 4744 21788
rect 4768 21786 4824 21788
rect 4848 21786 4904 21788
rect 4928 21786 4984 21788
rect 4688 21734 4714 21786
rect 4714 21734 4744 21786
rect 4768 21734 4778 21786
rect 4778 21734 4824 21786
rect 4848 21734 4894 21786
rect 4894 21734 4904 21786
rect 4928 21734 4958 21786
rect 4958 21734 4984 21786
rect 4688 21732 4744 21734
rect 4768 21732 4824 21734
rect 4848 21732 4904 21734
rect 4928 21732 4984 21734
rect 4688 20698 4744 20700
rect 4768 20698 4824 20700
rect 4848 20698 4904 20700
rect 4928 20698 4984 20700
rect 4688 20646 4714 20698
rect 4714 20646 4744 20698
rect 4768 20646 4778 20698
rect 4778 20646 4824 20698
rect 4848 20646 4894 20698
rect 4894 20646 4904 20698
rect 4928 20646 4958 20698
rect 4958 20646 4984 20698
rect 4688 20644 4744 20646
rect 4768 20644 4824 20646
rect 4848 20644 4904 20646
rect 4928 20644 4984 20646
rect 4688 19610 4744 19612
rect 4768 19610 4824 19612
rect 4848 19610 4904 19612
rect 4928 19610 4984 19612
rect 4688 19558 4714 19610
rect 4714 19558 4744 19610
rect 4768 19558 4778 19610
rect 4778 19558 4824 19610
rect 4848 19558 4894 19610
rect 4894 19558 4904 19610
rect 4928 19558 4958 19610
rect 4958 19558 4984 19610
rect 4688 19556 4744 19558
rect 4768 19556 4824 19558
rect 4848 19556 4904 19558
rect 4928 19556 4984 19558
rect 4688 18522 4744 18524
rect 4768 18522 4824 18524
rect 4848 18522 4904 18524
rect 4928 18522 4984 18524
rect 4688 18470 4714 18522
rect 4714 18470 4744 18522
rect 4768 18470 4778 18522
rect 4778 18470 4824 18522
rect 4848 18470 4894 18522
rect 4894 18470 4904 18522
rect 4928 18470 4958 18522
rect 4958 18470 4984 18522
rect 4688 18468 4744 18470
rect 4768 18468 4824 18470
rect 4848 18468 4904 18470
rect 4928 18468 4984 18470
rect 4688 17434 4744 17436
rect 4768 17434 4824 17436
rect 4848 17434 4904 17436
rect 4928 17434 4984 17436
rect 4688 17382 4714 17434
rect 4714 17382 4744 17434
rect 4768 17382 4778 17434
rect 4778 17382 4824 17434
rect 4848 17382 4894 17434
rect 4894 17382 4904 17434
rect 4928 17382 4958 17434
rect 4958 17382 4984 17434
rect 4688 17380 4744 17382
rect 4768 17380 4824 17382
rect 4848 17380 4904 17382
rect 4928 17380 4984 17382
rect 1490 15272 1546 15328
rect 1398 9152 1454 9208
rect 4688 16346 4744 16348
rect 4768 16346 4824 16348
rect 4848 16346 4904 16348
rect 4928 16346 4984 16348
rect 4688 16294 4714 16346
rect 4714 16294 4744 16346
rect 4768 16294 4778 16346
rect 4778 16294 4824 16346
rect 4848 16294 4894 16346
rect 4894 16294 4904 16346
rect 4928 16294 4958 16346
rect 4958 16294 4984 16346
rect 4688 16292 4744 16294
rect 4768 16292 4824 16294
rect 4848 16292 4904 16294
rect 4928 16292 4984 16294
rect 4688 15258 4744 15260
rect 4768 15258 4824 15260
rect 4848 15258 4904 15260
rect 4928 15258 4984 15260
rect 4688 15206 4714 15258
rect 4714 15206 4744 15258
rect 4768 15206 4778 15258
rect 4778 15206 4824 15258
rect 4848 15206 4894 15258
rect 4894 15206 4904 15258
rect 4928 15206 4958 15258
rect 4958 15206 4984 15258
rect 4688 15204 4744 15206
rect 4768 15204 4824 15206
rect 4848 15204 4904 15206
rect 4928 15204 4984 15206
rect 4688 14170 4744 14172
rect 4768 14170 4824 14172
rect 4848 14170 4904 14172
rect 4928 14170 4984 14172
rect 4688 14118 4714 14170
rect 4714 14118 4744 14170
rect 4768 14118 4778 14170
rect 4778 14118 4824 14170
rect 4848 14118 4894 14170
rect 4894 14118 4904 14170
rect 4928 14118 4958 14170
rect 4958 14118 4984 14170
rect 4688 14116 4744 14118
rect 4768 14116 4824 14118
rect 4848 14116 4904 14118
rect 4928 14116 4984 14118
rect 7562 21392 7618 21448
rect 8420 22330 8476 22332
rect 8500 22330 8556 22332
rect 8580 22330 8636 22332
rect 8660 22330 8716 22332
rect 8420 22278 8446 22330
rect 8446 22278 8476 22330
rect 8500 22278 8510 22330
rect 8510 22278 8556 22330
rect 8580 22278 8626 22330
rect 8626 22278 8636 22330
rect 8660 22278 8690 22330
rect 8690 22278 8716 22330
rect 8420 22276 8476 22278
rect 8500 22276 8556 22278
rect 8580 22276 8636 22278
rect 8660 22276 8716 22278
rect 8758 21972 8760 21992
rect 8760 21972 8812 21992
rect 8812 21972 8814 21992
rect 8758 21936 8814 21972
rect 8574 21548 8630 21584
rect 8574 21528 8576 21548
rect 8576 21528 8628 21548
rect 8628 21528 8630 21548
rect 8390 21428 8392 21448
rect 8392 21428 8444 21448
rect 8444 21428 8446 21448
rect 8390 21392 8446 21428
rect 8420 21242 8476 21244
rect 8500 21242 8556 21244
rect 8580 21242 8636 21244
rect 8660 21242 8716 21244
rect 8420 21190 8446 21242
rect 8446 21190 8476 21242
rect 8500 21190 8510 21242
rect 8510 21190 8556 21242
rect 8580 21190 8626 21242
rect 8626 21190 8636 21242
rect 8660 21190 8690 21242
rect 8690 21190 8716 21242
rect 8420 21188 8476 21190
rect 8500 21188 8556 21190
rect 8580 21188 8636 21190
rect 8660 21188 8716 21190
rect 8482 20848 8538 20904
rect 8420 20154 8476 20156
rect 8500 20154 8556 20156
rect 8580 20154 8636 20156
rect 8660 20154 8716 20156
rect 8420 20102 8446 20154
rect 8446 20102 8476 20154
rect 8500 20102 8510 20154
rect 8510 20102 8556 20154
rect 8580 20102 8626 20154
rect 8626 20102 8636 20154
rect 8660 20102 8690 20154
rect 8690 20102 8716 20154
rect 8420 20100 8476 20102
rect 8500 20100 8556 20102
rect 8580 20100 8636 20102
rect 8660 20100 8716 20102
rect 8420 19066 8476 19068
rect 8500 19066 8556 19068
rect 8580 19066 8636 19068
rect 8660 19066 8716 19068
rect 8420 19014 8446 19066
rect 8446 19014 8476 19066
rect 8500 19014 8510 19066
rect 8510 19014 8556 19066
rect 8580 19014 8626 19066
rect 8626 19014 8636 19066
rect 8660 19014 8690 19066
rect 8690 19014 8716 19066
rect 8420 19012 8476 19014
rect 8500 19012 8556 19014
rect 8580 19012 8636 19014
rect 8660 19012 8716 19014
rect 8420 17978 8476 17980
rect 8500 17978 8556 17980
rect 8580 17978 8636 17980
rect 8660 17978 8716 17980
rect 8420 17926 8446 17978
rect 8446 17926 8476 17978
rect 8500 17926 8510 17978
rect 8510 17926 8556 17978
rect 8580 17926 8626 17978
rect 8626 17926 8636 17978
rect 8660 17926 8690 17978
rect 8690 17926 8716 17978
rect 8420 17924 8476 17926
rect 8500 17924 8556 17926
rect 8580 17924 8636 17926
rect 8660 17924 8716 17926
rect 8420 16890 8476 16892
rect 8500 16890 8556 16892
rect 8580 16890 8636 16892
rect 8660 16890 8716 16892
rect 8420 16838 8446 16890
rect 8446 16838 8476 16890
rect 8500 16838 8510 16890
rect 8510 16838 8556 16890
rect 8580 16838 8626 16890
rect 8626 16838 8636 16890
rect 8660 16838 8690 16890
rect 8690 16838 8716 16890
rect 8420 16836 8476 16838
rect 8500 16836 8556 16838
rect 8580 16836 8636 16838
rect 8660 16836 8716 16838
rect 8420 15802 8476 15804
rect 8500 15802 8556 15804
rect 8580 15802 8636 15804
rect 8660 15802 8716 15804
rect 8420 15750 8446 15802
rect 8446 15750 8476 15802
rect 8500 15750 8510 15802
rect 8510 15750 8556 15802
rect 8580 15750 8626 15802
rect 8626 15750 8636 15802
rect 8660 15750 8690 15802
rect 8690 15750 8716 15802
rect 8420 15748 8476 15750
rect 8500 15748 8556 15750
rect 8580 15748 8636 15750
rect 8660 15748 8716 15750
rect 10046 22072 10102 22128
rect 10414 21256 10470 21312
rect 10690 21428 10692 21448
rect 10692 21428 10744 21448
rect 10744 21428 10746 21448
rect 10690 21392 10746 21428
rect 11702 22072 11758 22128
rect 10966 21548 11022 21584
rect 10966 21528 10968 21548
rect 10968 21528 11020 21548
rect 11020 21528 11022 21548
rect 11242 21936 11298 21992
rect 11242 21392 11298 21448
rect 10690 19372 10746 19408
rect 10690 19352 10692 19372
rect 10692 19352 10744 19372
rect 10744 19352 10746 19372
rect 9862 15156 9918 15192
rect 9862 15136 9864 15156
rect 9864 15136 9916 15156
rect 9916 15136 9918 15156
rect 11150 15136 11206 15192
rect 8420 14714 8476 14716
rect 8500 14714 8556 14716
rect 8580 14714 8636 14716
rect 8660 14714 8716 14716
rect 8420 14662 8446 14714
rect 8446 14662 8476 14714
rect 8500 14662 8510 14714
rect 8510 14662 8556 14714
rect 8580 14662 8626 14714
rect 8626 14662 8636 14714
rect 8660 14662 8690 14714
rect 8690 14662 8716 14714
rect 8420 14660 8476 14662
rect 8500 14660 8556 14662
rect 8580 14660 8636 14662
rect 8660 14660 8716 14662
rect 4688 13082 4744 13084
rect 4768 13082 4824 13084
rect 4848 13082 4904 13084
rect 4928 13082 4984 13084
rect 4688 13030 4714 13082
rect 4714 13030 4744 13082
rect 4768 13030 4778 13082
rect 4778 13030 4824 13082
rect 4848 13030 4894 13082
rect 4894 13030 4904 13082
rect 4928 13030 4958 13082
rect 4958 13030 4984 13082
rect 4688 13028 4744 13030
rect 4768 13028 4824 13030
rect 4848 13028 4904 13030
rect 4928 13028 4984 13030
rect 8420 13626 8476 13628
rect 8500 13626 8556 13628
rect 8580 13626 8636 13628
rect 8660 13626 8716 13628
rect 8420 13574 8446 13626
rect 8446 13574 8476 13626
rect 8500 13574 8510 13626
rect 8510 13574 8556 13626
rect 8580 13574 8626 13626
rect 8626 13574 8636 13626
rect 8660 13574 8690 13626
rect 8690 13574 8716 13626
rect 8420 13572 8476 13574
rect 8500 13572 8556 13574
rect 8580 13572 8636 13574
rect 8660 13572 8716 13574
rect 4688 11994 4744 11996
rect 4768 11994 4824 11996
rect 4848 11994 4904 11996
rect 4928 11994 4984 11996
rect 4688 11942 4714 11994
rect 4714 11942 4744 11994
rect 4768 11942 4778 11994
rect 4778 11942 4824 11994
rect 4848 11942 4894 11994
rect 4894 11942 4904 11994
rect 4928 11942 4958 11994
rect 4958 11942 4984 11994
rect 4688 11940 4744 11942
rect 4768 11940 4824 11942
rect 4848 11940 4904 11942
rect 4928 11940 4984 11942
rect 8420 12538 8476 12540
rect 8500 12538 8556 12540
rect 8580 12538 8636 12540
rect 8660 12538 8716 12540
rect 8420 12486 8446 12538
rect 8446 12486 8476 12538
rect 8500 12486 8510 12538
rect 8510 12486 8556 12538
rect 8580 12486 8626 12538
rect 8626 12486 8636 12538
rect 8660 12486 8690 12538
rect 8690 12486 8716 12538
rect 8420 12484 8476 12486
rect 8500 12484 8556 12486
rect 8580 12484 8636 12486
rect 8660 12484 8716 12486
rect 4688 10906 4744 10908
rect 4768 10906 4824 10908
rect 4848 10906 4904 10908
rect 4928 10906 4984 10908
rect 4688 10854 4714 10906
rect 4714 10854 4744 10906
rect 4768 10854 4778 10906
rect 4778 10854 4824 10906
rect 4848 10854 4894 10906
rect 4894 10854 4904 10906
rect 4928 10854 4958 10906
rect 4958 10854 4984 10906
rect 4688 10852 4744 10854
rect 4768 10852 4824 10854
rect 4848 10852 4904 10854
rect 4928 10852 4984 10854
rect 8420 11450 8476 11452
rect 8500 11450 8556 11452
rect 8580 11450 8636 11452
rect 8660 11450 8716 11452
rect 8420 11398 8446 11450
rect 8446 11398 8476 11450
rect 8500 11398 8510 11450
rect 8510 11398 8556 11450
rect 8580 11398 8626 11450
rect 8626 11398 8636 11450
rect 8660 11398 8690 11450
rect 8690 11398 8716 11450
rect 8420 11396 8476 11398
rect 8500 11396 8556 11398
rect 8580 11396 8636 11398
rect 8660 11396 8716 11398
rect 4688 9818 4744 9820
rect 4768 9818 4824 9820
rect 4848 9818 4904 9820
rect 4928 9818 4984 9820
rect 4688 9766 4714 9818
rect 4714 9766 4744 9818
rect 4768 9766 4778 9818
rect 4778 9766 4824 9818
rect 4848 9766 4894 9818
rect 4894 9766 4904 9818
rect 4928 9766 4958 9818
rect 4958 9766 4984 9818
rect 4688 9764 4744 9766
rect 4768 9764 4824 9766
rect 4848 9764 4904 9766
rect 4928 9764 4984 9766
rect 8420 10362 8476 10364
rect 8500 10362 8556 10364
rect 8580 10362 8636 10364
rect 8660 10362 8716 10364
rect 8420 10310 8446 10362
rect 8446 10310 8476 10362
rect 8500 10310 8510 10362
rect 8510 10310 8556 10362
rect 8580 10310 8626 10362
rect 8626 10310 8636 10362
rect 8660 10310 8690 10362
rect 8690 10310 8716 10362
rect 8420 10308 8476 10310
rect 8500 10308 8556 10310
rect 8580 10308 8636 10310
rect 8660 10308 8716 10310
rect 10966 14456 11022 14512
rect 10782 13912 10838 13968
rect 9678 13368 9734 13424
rect 10506 12144 10562 12200
rect 11702 21548 11758 21584
rect 11702 21528 11704 21548
rect 11704 21528 11756 21548
rect 11756 21528 11758 21548
rect 12152 21786 12208 21788
rect 12232 21786 12288 21788
rect 12312 21786 12368 21788
rect 12392 21786 12448 21788
rect 12152 21734 12178 21786
rect 12178 21734 12208 21786
rect 12232 21734 12242 21786
rect 12242 21734 12288 21786
rect 12312 21734 12358 21786
rect 12358 21734 12368 21786
rect 12392 21734 12422 21786
rect 12422 21734 12448 21786
rect 12152 21732 12208 21734
rect 12232 21732 12288 21734
rect 12312 21732 12368 21734
rect 12392 21732 12448 21734
rect 12346 21528 12402 21584
rect 12346 21004 12402 21040
rect 12346 20984 12348 21004
rect 12348 20984 12400 21004
rect 12400 20984 12402 21004
rect 12152 20698 12208 20700
rect 12232 20698 12288 20700
rect 12312 20698 12368 20700
rect 12392 20698 12448 20700
rect 12152 20646 12178 20698
rect 12178 20646 12208 20698
rect 12232 20646 12242 20698
rect 12242 20646 12288 20698
rect 12312 20646 12358 20698
rect 12358 20646 12368 20698
rect 12392 20646 12422 20698
rect 12422 20646 12448 20698
rect 12152 20644 12208 20646
rect 12232 20644 12288 20646
rect 12312 20644 12368 20646
rect 12392 20644 12448 20646
rect 12152 19610 12208 19612
rect 12232 19610 12288 19612
rect 12312 19610 12368 19612
rect 12392 19610 12448 19612
rect 12152 19558 12178 19610
rect 12178 19558 12208 19610
rect 12232 19558 12242 19610
rect 12242 19558 12288 19610
rect 12312 19558 12358 19610
rect 12358 19558 12368 19610
rect 12392 19558 12422 19610
rect 12422 19558 12448 19610
rect 12152 19556 12208 19558
rect 12232 19556 12288 19558
rect 12312 19556 12368 19558
rect 12392 19556 12448 19558
rect 11702 19216 11758 19272
rect 12152 18522 12208 18524
rect 12232 18522 12288 18524
rect 12312 18522 12368 18524
rect 12392 18522 12448 18524
rect 12152 18470 12178 18522
rect 12178 18470 12208 18522
rect 12232 18470 12242 18522
rect 12242 18470 12288 18522
rect 12312 18470 12358 18522
rect 12358 18470 12368 18522
rect 12392 18470 12422 18522
rect 12422 18470 12448 18522
rect 12152 18468 12208 18470
rect 12232 18468 12288 18470
rect 12312 18468 12368 18470
rect 12392 18468 12448 18470
rect 12152 17434 12208 17436
rect 12232 17434 12288 17436
rect 12312 17434 12368 17436
rect 12392 17434 12448 17436
rect 12152 17382 12178 17434
rect 12178 17382 12208 17434
rect 12232 17382 12242 17434
rect 12242 17382 12288 17434
rect 12312 17382 12358 17434
rect 12358 17382 12368 17434
rect 12392 17382 12422 17434
rect 12422 17382 12448 17434
rect 12152 17380 12208 17382
rect 12232 17380 12288 17382
rect 12312 17380 12368 17382
rect 12392 17380 12448 17382
rect 12152 16346 12208 16348
rect 12232 16346 12288 16348
rect 12312 16346 12368 16348
rect 12392 16346 12448 16348
rect 12152 16294 12178 16346
rect 12178 16294 12208 16346
rect 12232 16294 12242 16346
rect 12242 16294 12288 16346
rect 12312 16294 12358 16346
rect 12358 16294 12368 16346
rect 12392 16294 12422 16346
rect 12422 16294 12448 16346
rect 12152 16292 12208 16294
rect 12232 16292 12288 16294
rect 12312 16292 12368 16294
rect 12392 16292 12448 16294
rect 12152 15258 12208 15260
rect 12232 15258 12288 15260
rect 12312 15258 12368 15260
rect 12392 15258 12448 15260
rect 12152 15206 12178 15258
rect 12178 15206 12208 15258
rect 12232 15206 12242 15258
rect 12242 15206 12288 15258
rect 12312 15206 12358 15258
rect 12358 15206 12368 15258
rect 12392 15206 12422 15258
rect 12422 15206 12448 15258
rect 12152 15204 12208 15206
rect 12232 15204 12288 15206
rect 12312 15204 12368 15206
rect 12392 15204 12448 15206
rect 12806 21936 12862 21992
rect 13542 21528 13598 21584
rect 13358 20984 13414 21040
rect 15884 22330 15940 22332
rect 15964 22330 16020 22332
rect 16044 22330 16100 22332
rect 16124 22330 16180 22332
rect 15884 22278 15910 22330
rect 15910 22278 15940 22330
rect 15964 22278 15974 22330
rect 15974 22278 16020 22330
rect 16044 22278 16090 22330
rect 16090 22278 16100 22330
rect 16124 22278 16154 22330
rect 16154 22278 16180 22330
rect 15884 22276 15940 22278
rect 15964 22276 16020 22278
rect 16044 22276 16100 22278
rect 16124 22276 16180 22278
rect 12152 14170 12208 14172
rect 12232 14170 12288 14172
rect 12312 14170 12368 14172
rect 12392 14170 12448 14172
rect 12152 14118 12178 14170
rect 12178 14118 12208 14170
rect 12232 14118 12242 14170
rect 12242 14118 12288 14170
rect 12312 14118 12358 14170
rect 12358 14118 12368 14170
rect 12392 14118 12422 14170
rect 12422 14118 12448 14170
rect 12152 14116 12208 14118
rect 12232 14116 12288 14118
rect 12312 14116 12368 14118
rect 12392 14116 12448 14118
rect 13082 13932 13138 13968
rect 13082 13912 13084 13932
rect 13084 13912 13136 13932
rect 13136 13912 13138 13932
rect 12152 13082 12208 13084
rect 12232 13082 12288 13084
rect 12312 13082 12368 13084
rect 12392 13082 12448 13084
rect 12152 13030 12178 13082
rect 12178 13030 12208 13082
rect 12232 13030 12242 13082
rect 12242 13030 12288 13082
rect 12312 13030 12358 13082
rect 12358 13030 12368 13082
rect 12392 13030 12422 13082
rect 12422 13030 12448 13082
rect 12152 13028 12208 13030
rect 12232 13028 12288 13030
rect 12312 13028 12368 13030
rect 12392 13028 12448 13030
rect 12254 12144 12310 12200
rect 12152 11994 12208 11996
rect 12232 11994 12288 11996
rect 12312 11994 12368 11996
rect 12392 11994 12448 11996
rect 12152 11942 12178 11994
rect 12178 11942 12208 11994
rect 12232 11942 12242 11994
rect 12242 11942 12288 11994
rect 12312 11942 12358 11994
rect 12358 11942 12368 11994
rect 12392 11942 12422 11994
rect 12422 11942 12448 11994
rect 12152 11940 12208 11942
rect 12232 11940 12288 11942
rect 12312 11940 12368 11942
rect 12392 11940 12448 11942
rect 14186 20984 14242 21040
rect 14462 21256 14518 21312
rect 15884 21242 15940 21244
rect 15964 21242 16020 21244
rect 16044 21242 16100 21244
rect 16124 21242 16180 21244
rect 15884 21190 15910 21242
rect 15910 21190 15940 21242
rect 15964 21190 15974 21242
rect 15974 21190 16020 21242
rect 16044 21190 16090 21242
rect 16090 21190 16100 21242
rect 16124 21190 16154 21242
rect 16154 21190 16180 21242
rect 15884 21188 15940 21190
rect 15964 21188 16020 21190
rect 16044 21188 16100 21190
rect 16124 21188 16180 21190
rect 15884 20154 15940 20156
rect 15964 20154 16020 20156
rect 16044 20154 16100 20156
rect 16124 20154 16180 20156
rect 15884 20102 15910 20154
rect 15910 20102 15940 20154
rect 15964 20102 15974 20154
rect 15974 20102 16020 20154
rect 16044 20102 16090 20154
rect 16090 20102 16100 20154
rect 16124 20102 16154 20154
rect 16154 20102 16180 20154
rect 15884 20100 15940 20102
rect 15964 20100 16020 20102
rect 16044 20100 16100 20102
rect 16124 20100 16180 20102
rect 17314 20984 17370 21040
rect 18050 21392 18106 21448
rect 15474 19216 15530 19272
rect 15884 19066 15940 19068
rect 15964 19066 16020 19068
rect 16044 19066 16100 19068
rect 16124 19066 16180 19068
rect 15884 19014 15910 19066
rect 15910 19014 15940 19066
rect 15964 19014 15974 19066
rect 15974 19014 16020 19066
rect 16044 19014 16090 19066
rect 16090 19014 16100 19066
rect 16124 19014 16154 19066
rect 16154 19014 16180 19066
rect 15884 19012 15940 19014
rect 15964 19012 16020 19014
rect 16044 19012 16100 19014
rect 16124 19012 16180 19014
rect 15474 16652 15530 16688
rect 15474 16632 15476 16652
rect 15476 16632 15528 16652
rect 15528 16632 15530 16652
rect 15198 13232 15254 13288
rect 12152 10906 12208 10908
rect 12232 10906 12288 10908
rect 12312 10906 12368 10908
rect 12392 10906 12448 10908
rect 12152 10854 12178 10906
rect 12178 10854 12208 10906
rect 12232 10854 12242 10906
rect 12242 10854 12288 10906
rect 12312 10854 12358 10906
rect 12358 10854 12368 10906
rect 12392 10854 12422 10906
rect 12422 10854 12448 10906
rect 12152 10852 12208 10854
rect 12232 10852 12288 10854
rect 12312 10852 12368 10854
rect 12392 10852 12448 10854
rect 8420 9274 8476 9276
rect 8500 9274 8556 9276
rect 8580 9274 8636 9276
rect 8660 9274 8716 9276
rect 8420 9222 8446 9274
rect 8446 9222 8476 9274
rect 8500 9222 8510 9274
rect 8510 9222 8556 9274
rect 8580 9222 8626 9274
rect 8626 9222 8636 9274
rect 8660 9222 8690 9274
rect 8690 9222 8716 9274
rect 8420 9220 8476 9222
rect 8500 9220 8556 9222
rect 8580 9220 8636 9222
rect 8660 9220 8716 9222
rect 12152 9818 12208 9820
rect 12232 9818 12288 9820
rect 12312 9818 12368 9820
rect 12392 9818 12448 9820
rect 12152 9766 12178 9818
rect 12178 9766 12208 9818
rect 12232 9766 12242 9818
rect 12242 9766 12288 9818
rect 12312 9766 12358 9818
rect 12358 9766 12368 9818
rect 12392 9766 12422 9818
rect 12422 9766 12448 9818
rect 12152 9764 12208 9766
rect 12232 9764 12288 9766
rect 12312 9764 12368 9766
rect 12392 9764 12448 9766
rect 4688 8730 4744 8732
rect 4768 8730 4824 8732
rect 4848 8730 4904 8732
rect 4928 8730 4984 8732
rect 4688 8678 4714 8730
rect 4714 8678 4744 8730
rect 4768 8678 4778 8730
rect 4778 8678 4824 8730
rect 4848 8678 4894 8730
rect 4894 8678 4904 8730
rect 4928 8678 4958 8730
rect 4958 8678 4984 8730
rect 4688 8676 4744 8678
rect 4768 8676 4824 8678
rect 4848 8676 4904 8678
rect 4928 8676 4984 8678
rect 8420 8186 8476 8188
rect 8500 8186 8556 8188
rect 8580 8186 8636 8188
rect 8660 8186 8716 8188
rect 8420 8134 8446 8186
rect 8446 8134 8476 8186
rect 8500 8134 8510 8186
rect 8510 8134 8556 8186
rect 8580 8134 8626 8186
rect 8626 8134 8636 8186
rect 8660 8134 8690 8186
rect 8690 8134 8716 8186
rect 8420 8132 8476 8134
rect 8500 8132 8556 8134
rect 8580 8132 8636 8134
rect 8660 8132 8716 8134
rect 4688 7642 4744 7644
rect 4768 7642 4824 7644
rect 4848 7642 4904 7644
rect 4928 7642 4984 7644
rect 4688 7590 4714 7642
rect 4714 7590 4744 7642
rect 4768 7590 4778 7642
rect 4778 7590 4824 7642
rect 4848 7590 4894 7642
rect 4894 7590 4904 7642
rect 4928 7590 4958 7642
rect 4958 7590 4984 7642
rect 4688 7588 4744 7590
rect 4768 7588 4824 7590
rect 4848 7588 4904 7590
rect 4928 7588 4984 7590
rect 12152 8730 12208 8732
rect 12232 8730 12288 8732
rect 12312 8730 12368 8732
rect 12392 8730 12448 8732
rect 12152 8678 12178 8730
rect 12178 8678 12208 8730
rect 12232 8678 12242 8730
rect 12242 8678 12288 8730
rect 12312 8678 12358 8730
rect 12358 8678 12368 8730
rect 12392 8678 12422 8730
rect 12422 8678 12448 8730
rect 12152 8676 12208 8678
rect 12232 8676 12288 8678
rect 12312 8676 12368 8678
rect 12392 8676 12448 8678
rect 8420 7098 8476 7100
rect 8500 7098 8556 7100
rect 8580 7098 8636 7100
rect 8660 7098 8716 7100
rect 8420 7046 8446 7098
rect 8446 7046 8476 7098
rect 8500 7046 8510 7098
rect 8510 7046 8556 7098
rect 8580 7046 8626 7098
rect 8626 7046 8636 7098
rect 8660 7046 8690 7098
rect 8690 7046 8716 7098
rect 8420 7044 8476 7046
rect 8500 7044 8556 7046
rect 8580 7044 8636 7046
rect 8660 7044 8716 7046
rect 4688 6554 4744 6556
rect 4768 6554 4824 6556
rect 4848 6554 4904 6556
rect 4928 6554 4984 6556
rect 4688 6502 4714 6554
rect 4714 6502 4744 6554
rect 4768 6502 4778 6554
rect 4778 6502 4824 6554
rect 4848 6502 4894 6554
rect 4894 6502 4904 6554
rect 4928 6502 4958 6554
rect 4958 6502 4984 6554
rect 4688 6500 4744 6502
rect 4768 6500 4824 6502
rect 4848 6500 4904 6502
rect 4928 6500 4984 6502
rect 12152 7642 12208 7644
rect 12232 7642 12288 7644
rect 12312 7642 12368 7644
rect 12392 7642 12448 7644
rect 12152 7590 12178 7642
rect 12178 7590 12208 7642
rect 12232 7590 12242 7642
rect 12242 7590 12288 7642
rect 12312 7590 12358 7642
rect 12358 7590 12368 7642
rect 12392 7590 12422 7642
rect 12422 7590 12448 7642
rect 12152 7588 12208 7590
rect 12232 7588 12288 7590
rect 12312 7588 12368 7590
rect 12392 7588 12448 7590
rect 15014 12280 15070 12336
rect 11886 7248 11942 7304
rect 8420 6010 8476 6012
rect 8500 6010 8556 6012
rect 8580 6010 8636 6012
rect 8660 6010 8716 6012
rect 8420 5958 8446 6010
rect 8446 5958 8476 6010
rect 8500 5958 8510 6010
rect 8510 5958 8556 6010
rect 8580 5958 8626 6010
rect 8626 5958 8636 6010
rect 8660 5958 8690 6010
rect 8690 5958 8716 6010
rect 8420 5956 8476 5958
rect 8500 5956 8556 5958
rect 8580 5956 8636 5958
rect 8660 5956 8716 5958
rect 12152 6554 12208 6556
rect 12232 6554 12288 6556
rect 12312 6554 12368 6556
rect 12392 6554 12448 6556
rect 12152 6502 12178 6554
rect 12178 6502 12208 6554
rect 12232 6502 12242 6554
rect 12242 6502 12288 6554
rect 12312 6502 12358 6554
rect 12358 6502 12368 6554
rect 12392 6502 12422 6554
rect 12422 6502 12448 6554
rect 12152 6500 12208 6502
rect 12232 6500 12288 6502
rect 12312 6500 12368 6502
rect 12392 6500 12448 6502
rect 14554 7828 14556 7848
rect 14556 7828 14608 7848
rect 14608 7828 14610 7848
rect 14554 7792 14610 7828
rect 4688 5466 4744 5468
rect 4768 5466 4824 5468
rect 4848 5466 4904 5468
rect 4928 5466 4984 5468
rect 4688 5414 4714 5466
rect 4714 5414 4744 5466
rect 4768 5414 4778 5466
rect 4778 5414 4824 5466
rect 4848 5414 4894 5466
rect 4894 5414 4904 5466
rect 4928 5414 4958 5466
rect 4958 5414 4984 5466
rect 4688 5412 4744 5414
rect 4768 5412 4824 5414
rect 4848 5412 4904 5414
rect 4928 5412 4984 5414
rect 12152 5466 12208 5468
rect 12232 5466 12288 5468
rect 12312 5466 12368 5468
rect 12392 5466 12448 5468
rect 12152 5414 12178 5466
rect 12178 5414 12208 5466
rect 12232 5414 12242 5466
rect 12242 5414 12288 5466
rect 12312 5414 12358 5466
rect 12358 5414 12368 5466
rect 12392 5414 12422 5466
rect 12422 5414 12448 5466
rect 12152 5412 12208 5414
rect 12232 5412 12288 5414
rect 12312 5412 12368 5414
rect 12392 5412 12448 5414
rect 15884 17978 15940 17980
rect 15964 17978 16020 17980
rect 16044 17978 16100 17980
rect 16124 17978 16180 17980
rect 15884 17926 15910 17978
rect 15910 17926 15940 17978
rect 15964 17926 15974 17978
rect 15974 17926 16020 17978
rect 16044 17926 16090 17978
rect 16090 17926 16100 17978
rect 16124 17926 16154 17978
rect 16154 17926 16180 17978
rect 15884 17924 15940 17926
rect 15964 17924 16020 17926
rect 16044 17924 16100 17926
rect 16124 17924 16180 17926
rect 15884 16890 15940 16892
rect 15964 16890 16020 16892
rect 16044 16890 16100 16892
rect 16124 16890 16180 16892
rect 15884 16838 15910 16890
rect 15910 16838 15940 16890
rect 15964 16838 15974 16890
rect 15974 16838 16020 16890
rect 16044 16838 16090 16890
rect 16090 16838 16100 16890
rect 16124 16838 16154 16890
rect 16154 16838 16180 16890
rect 15884 16836 15940 16838
rect 15964 16836 16020 16838
rect 16044 16836 16100 16838
rect 16124 16836 16180 16838
rect 15884 15802 15940 15804
rect 15964 15802 16020 15804
rect 16044 15802 16100 15804
rect 16124 15802 16180 15804
rect 15884 15750 15910 15802
rect 15910 15750 15940 15802
rect 15964 15750 15974 15802
rect 15974 15750 16020 15802
rect 16044 15750 16090 15802
rect 16090 15750 16100 15802
rect 16124 15750 16154 15802
rect 16154 15750 16180 15802
rect 15884 15748 15940 15750
rect 15964 15748 16020 15750
rect 16044 15748 16100 15750
rect 16124 15748 16180 15750
rect 15884 14714 15940 14716
rect 15964 14714 16020 14716
rect 16044 14714 16100 14716
rect 16124 14714 16180 14716
rect 15884 14662 15910 14714
rect 15910 14662 15940 14714
rect 15964 14662 15974 14714
rect 15974 14662 16020 14714
rect 16044 14662 16090 14714
rect 16090 14662 16100 14714
rect 16124 14662 16154 14714
rect 16154 14662 16180 14714
rect 15884 14660 15940 14662
rect 15964 14660 16020 14662
rect 16044 14660 16100 14662
rect 16124 14660 16180 14662
rect 15884 13626 15940 13628
rect 15964 13626 16020 13628
rect 16044 13626 16100 13628
rect 16124 13626 16180 13628
rect 15884 13574 15910 13626
rect 15910 13574 15940 13626
rect 15964 13574 15974 13626
rect 15974 13574 16020 13626
rect 16044 13574 16090 13626
rect 16090 13574 16100 13626
rect 16124 13574 16154 13626
rect 16154 13574 16180 13626
rect 15884 13572 15940 13574
rect 15964 13572 16020 13574
rect 16044 13572 16100 13574
rect 16124 13572 16180 13574
rect 15934 12724 15936 12744
rect 15936 12724 15988 12744
rect 15988 12724 15990 12744
rect 15934 12688 15990 12724
rect 15884 12538 15940 12540
rect 15964 12538 16020 12540
rect 16044 12538 16100 12540
rect 16124 12538 16180 12540
rect 15884 12486 15910 12538
rect 15910 12486 15940 12538
rect 15964 12486 15974 12538
rect 15974 12486 16020 12538
rect 16044 12486 16090 12538
rect 16090 12486 16100 12538
rect 16124 12486 16154 12538
rect 16154 12486 16180 12538
rect 15884 12484 15940 12486
rect 15964 12484 16020 12486
rect 16044 12484 16100 12486
rect 16124 12484 16180 12486
rect 15290 7948 15346 7984
rect 15290 7928 15292 7948
rect 15292 7928 15344 7948
rect 15344 7928 15346 7948
rect 15884 11450 15940 11452
rect 15964 11450 16020 11452
rect 16044 11450 16100 11452
rect 16124 11450 16180 11452
rect 15884 11398 15910 11450
rect 15910 11398 15940 11450
rect 15964 11398 15974 11450
rect 15974 11398 16020 11450
rect 16044 11398 16090 11450
rect 16090 11398 16100 11450
rect 16124 11398 16154 11450
rect 16154 11398 16180 11450
rect 15884 11396 15940 11398
rect 15964 11396 16020 11398
rect 16044 11396 16100 11398
rect 16124 11396 16180 11398
rect 16670 14320 16726 14376
rect 17774 15020 17830 15056
rect 17774 15000 17776 15020
rect 17776 15000 17828 15020
rect 17828 15000 17830 15020
rect 17406 14864 17462 14920
rect 15884 10362 15940 10364
rect 15964 10362 16020 10364
rect 16044 10362 16100 10364
rect 16124 10362 16180 10364
rect 15884 10310 15910 10362
rect 15910 10310 15940 10362
rect 15964 10310 15974 10362
rect 15974 10310 16020 10362
rect 16044 10310 16090 10362
rect 16090 10310 16100 10362
rect 16124 10310 16154 10362
rect 16154 10310 16180 10362
rect 15884 10308 15940 10310
rect 15964 10308 16020 10310
rect 16044 10308 16100 10310
rect 16124 10308 16180 10310
rect 17130 12688 17186 12744
rect 16486 10376 16542 10432
rect 15884 9274 15940 9276
rect 15964 9274 16020 9276
rect 16044 9274 16100 9276
rect 16124 9274 16180 9276
rect 15884 9222 15910 9274
rect 15910 9222 15940 9274
rect 15964 9222 15974 9274
rect 15974 9222 16020 9274
rect 16044 9222 16090 9274
rect 16090 9222 16100 9274
rect 16124 9222 16154 9274
rect 16154 9222 16180 9274
rect 15884 9220 15940 9222
rect 15964 9220 16020 9222
rect 16044 9220 16100 9222
rect 16124 9220 16180 9222
rect 15884 8186 15940 8188
rect 15964 8186 16020 8188
rect 16044 8186 16100 8188
rect 16124 8186 16180 8188
rect 15884 8134 15910 8186
rect 15910 8134 15940 8186
rect 15964 8134 15974 8186
rect 15974 8134 16020 8186
rect 16044 8134 16090 8186
rect 16090 8134 16100 8186
rect 16124 8134 16154 8186
rect 16154 8134 16180 8186
rect 15884 8132 15940 8134
rect 15964 8132 16020 8134
rect 16044 8132 16100 8134
rect 16124 8132 16180 8134
rect 15842 7404 15898 7440
rect 15842 7384 15844 7404
rect 15844 7384 15896 7404
rect 15896 7384 15898 7404
rect 15884 7098 15940 7100
rect 15964 7098 16020 7100
rect 16044 7098 16100 7100
rect 16124 7098 16180 7100
rect 15884 7046 15910 7098
rect 15910 7046 15940 7098
rect 15964 7046 15974 7098
rect 15974 7046 16020 7098
rect 16044 7046 16090 7098
rect 16090 7046 16100 7098
rect 16124 7046 16154 7098
rect 16154 7046 16180 7098
rect 15884 7044 15940 7046
rect 15964 7044 16020 7046
rect 16044 7044 16100 7046
rect 16124 7044 16180 7046
rect 15884 6010 15940 6012
rect 15964 6010 16020 6012
rect 16044 6010 16100 6012
rect 16124 6010 16180 6012
rect 15884 5958 15910 6010
rect 15910 5958 15940 6010
rect 15964 5958 15974 6010
rect 15974 5958 16020 6010
rect 16044 5958 16090 6010
rect 16090 5958 16100 6010
rect 16124 5958 16154 6010
rect 16154 5958 16180 6010
rect 15884 5956 15940 5958
rect 15964 5956 16020 5958
rect 16044 5956 16100 5958
rect 16124 5956 16180 5958
rect 16486 7828 16488 7848
rect 16488 7828 16540 7848
rect 16540 7828 16542 7848
rect 16486 7792 16542 7828
rect 16854 9596 16856 9616
rect 16856 9596 16908 9616
rect 16908 9596 16910 9616
rect 16854 9560 16910 9596
rect 17222 12280 17278 12336
rect 18050 16668 18052 16688
rect 18052 16668 18104 16688
rect 18104 16668 18106 16688
rect 18050 16632 18106 16668
rect 18050 14728 18106 14784
rect 17498 11600 17554 11656
rect 17406 10124 17462 10160
rect 17406 10104 17408 10124
rect 17408 10104 17460 10124
rect 17460 10104 17462 10124
rect 18050 10376 18106 10432
rect 19154 21528 19210 21584
rect 19616 21786 19672 21788
rect 19696 21786 19752 21788
rect 19776 21786 19832 21788
rect 19856 21786 19912 21788
rect 19616 21734 19642 21786
rect 19642 21734 19672 21786
rect 19696 21734 19706 21786
rect 19706 21734 19752 21786
rect 19776 21734 19822 21786
rect 19822 21734 19832 21786
rect 19856 21734 19886 21786
rect 19886 21734 19912 21786
rect 19616 21732 19672 21734
rect 19696 21732 19752 21734
rect 19776 21732 19832 21734
rect 19856 21732 19912 21734
rect 19616 20698 19672 20700
rect 19696 20698 19752 20700
rect 19776 20698 19832 20700
rect 19856 20698 19912 20700
rect 19616 20646 19642 20698
rect 19642 20646 19672 20698
rect 19696 20646 19706 20698
rect 19706 20646 19752 20698
rect 19776 20646 19822 20698
rect 19822 20646 19832 20698
rect 19856 20646 19886 20698
rect 19886 20646 19912 20698
rect 19616 20644 19672 20646
rect 19696 20644 19752 20646
rect 19776 20644 19832 20646
rect 19856 20644 19912 20646
rect 19246 19352 19302 19408
rect 18418 14456 18474 14512
rect 18326 13232 18382 13288
rect 19616 19610 19672 19612
rect 19696 19610 19752 19612
rect 19776 19610 19832 19612
rect 19856 19610 19912 19612
rect 19616 19558 19642 19610
rect 19642 19558 19672 19610
rect 19696 19558 19706 19610
rect 19706 19558 19752 19610
rect 19776 19558 19822 19610
rect 19822 19558 19832 19610
rect 19856 19558 19886 19610
rect 19886 19558 19912 19610
rect 19616 19556 19672 19558
rect 19696 19556 19752 19558
rect 19776 19556 19832 19558
rect 19856 19556 19912 19558
rect 19616 18522 19672 18524
rect 19696 18522 19752 18524
rect 19776 18522 19832 18524
rect 19856 18522 19912 18524
rect 19616 18470 19642 18522
rect 19642 18470 19672 18522
rect 19696 18470 19706 18522
rect 19706 18470 19752 18522
rect 19776 18470 19822 18522
rect 19822 18470 19832 18522
rect 19856 18470 19886 18522
rect 19886 18470 19912 18522
rect 19616 18468 19672 18470
rect 19696 18468 19752 18470
rect 19776 18468 19832 18470
rect 19856 18468 19912 18470
rect 18694 10412 18696 10432
rect 18696 10412 18748 10432
rect 18748 10412 18750 10432
rect 18694 10376 18750 10412
rect 17314 7948 17370 7984
rect 17314 7928 17316 7948
rect 17316 7928 17368 7948
rect 17368 7928 17370 7948
rect 17406 7248 17462 7304
rect 18142 7812 18198 7848
rect 18142 7792 18144 7812
rect 18144 7792 18196 7812
rect 18196 7792 18198 7812
rect 8420 4922 8476 4924
rect 8500 4922 8556 4924
rect 8580 4922 8636 4924
rect 8660 4922 8716 4924
rect 8420 4870 8446 4922
rect 8446 4870 8476 4922
rect 8500 4870 8510 4922
rect 8510 4870 8556 4922
rect 8580 4870 8626 4922
rect 8626 4870 8636 4922
rect 8660 4870 8690 4922
rect 8690 4870 8716 4922
rect 8420 4868 8476 4870
rect 8500 4868 8556 4870
rect 8580 4868 8636 4870
rect 8660 4868 8716 4870
rect 15884 4922 15940 4924
rect 15964 4922 16020 4924
rect 16044 4922 16100 4924
rect 16124 4922 16180 4924
rect 15884 4870 15910 4922
rect 15910 4870 15940 4922
rect 15964 4870 15974 4922
rect 15974 4870 16020 4922
rect 16044 4870 16090 4922
rect 16090 4870 16100 4922
rect 16124 4870 16154 4922
rect 16154 4870 16180 4922
rect 15884 4868 15940 4870
rect 15964 4868 16020 4870
rect 16044 4868 16100 4870
rect 16124 4868 16180 4870
rect 4688 4378 4744 4380
rect 4768 4378 4824 4380
rect 4848 4378 4904 4380
rect 4928 4378 4984 4380
rect 4688 4326 4714 4378
rect 4714 4326 4744 4378
rect 4768 4326 4778 4378
rect 4778 4326 4824 4378
rect 4848 4326 4894 4378
rect 4894 4326 4904 4378
rect 4928 4326 4958 4378
rect 4958 4326 4984 4378
rect 4688 4324 4744 4326
rect 4768 4324 4824 4326
rect 4848 4324 4904 4326
rect 4928 4324 4984 4326
rect 12152 4378 12208 4380
rect 12232 4378 12288 4380
rect 12312 4378 12368 4380
rect 12392 4378 12448 4380
rect 12152 4326 12178 4378
rect 12178 4326 12208 4378
rect 12232 4326 12242 4378
rect 12242 4326 12288 4378
rect 12312 4326 12358 4378
rect 12358 4326 12368 4378
rect 12392 4326 12422 4378
rect 12422 4326 12448 4378
rect 12152 4324 12208 4326
rect 12232 4324 12288 4326
rect 12312 4324 12368 4326
rect 12392 4324 12448 4326
rect 8420 3834 8476 3836
rect 8500 3834 8556 3836
rect 8580 3834 8636 3836
rect 8660 3834 8716 3836
rect 8420 3782 8446 3834
rect 8446 3782 8476 3834
rect 8500 3782 8510 3834
rect 8510 3782 8556 3834
rect 8580 3782 8626 3834
rect 8626 3782 8636 3834
rect 8660 3782 8690 3834
rect 8690 3782 8716 3834
rect 8420 3780 8476 3782
rect 8500 3780 8556 3782
rect 8580 3780 8636 3782
rect 8660 3780 8716 3782
rect 15884 3834 15940 3836
rect 15964 3834 16020 3836
rect 16044 3834 16100 3836
rect 16124 3834 16180 3836
rect 15884 3782 15910 3834
rect 15910 3782 15940 3834
rect 15964 3782 15974 3834
rect 15974 3782 16020 3834
rect 16044 3782 16090 3834
rect 16090 3782 16100 3834
rect 16124 3782 16154 3834
rect 16154 3782 16180 3834
rect 15884 3780 15940 3782
rect 15964 3780 16020 3782
rect 16044 3780 16100 3782
rect 16124 3780 16180 3782
rect 4688 3290 4744 3292
rect 4768 3290 4824 3292
rect 4848 3290 4904 3292
rect 4928 3290 4984 3292
rect 4688 3238 4714 3290
rect 4714 3238 4744 3290
rect 4768 3238 4778 3290
rect 4778 3238 4824 3290
rect 4848 3238 4894 3290
rect 4894 3238 4904 3290
rect 4928 3238 4958 3290
rect 4958 3238 4984 3290
rect 4688 3236 4744 3238
rect 4768 3236 4824 3238
rect 4848 3236 4904 3238
rect 4928 3236 4984 3238
rect 12152 3290 12208 3292
rect 12232 3290 12288 3292
rect 12312 3290 12368 3292
rect 12392 3290 12448 3292
rect 12152 3238 12178 3290
rect 12178 3238 12208 3290
rect 12232 3238 12242 3290
rect 12242 3238 12288 3290
rect 12312 3238 12358 3290
rect 12358 3238 12368 3290
rect 12392 3238 12422 3290
rect 12422 3238 12448 3290
rect 12152 3236 12208 3238
rect 12232 3236 12288 3238
rect 12312 3236 12368 3238
rect 12392 3236 12448 3238
rect 1398 3068 1400 3088
rect 1400 3068 1452 3088
rect 1452 3068 1454 3088
rect 1398 3032 1454 3068
rect 8420 2746 8476 2748
rect 8500 2746 8556 2748
rect 8580 2746 8636 2748
rect 8660 2746 8716 2748
rect 8420 2694 8446 2746
rect 8446 2694 8476 2746
rect 8500 2694 8510 2746
rect 8510 2694 8556 2746
rect 8580 2694 8626 2746
rect 8626 2694 8636 2746
rect 8660 2694 8690 2746
rect 8690 2694 8716 2746
rect 8420 2692 8476 2694
rect 8500 2692 8556 2694
rect 8580 2692 8636 2694
rect 8660 2692 8716 2694
rect 15884 2746 15940 2748
rect 15964 2746 16020 2748
rect 16044 2746 16100 2748
rect 16124 2746 16180 2748
rect 15884 2694 15910 2746
rect 15910 2694 15940 2746
rect 15964 2694 15974 2746
rect 15974 2694 16020 2746
rect 16044 2694 16090 2746
rect 16090 2694 16100 2746
rect 16124 2694 16154 2746
rect 16154 2694 16180 2746
rect 15884 2692 15940 2694
rect 15964 2692 16020 2694
rect 16044 2692 16100 2694
rect 16124 2692 16180 2694
rect 19616 17434 19672 17436
rect 19696 17434 19752 17436
rect 19776 17434 19832 17436
rect 19856 17434 19912 17436
rect 19616 17382 19642 17434
rect 19642 17382 19672 17434
rect 19696 17382 19706 17434
rect 19706 17382 19752 17434
rect 19776 17382 19822 17434
rect 19822 17382 19832 17434
rect 19856 17382 19886 17434
rect 19886 17382 19912 17434
rect 19616 17380 19672 17382
rect 19696 17380 19752 17382
rect 19776 17380 19832 17382
rect 19856 17380 19912 17382
rect 19522 16904 19578 16960
rect 19430 16532 19432 16552
rect 19432 16532 19484 16552
rect 19484 16532 19486 16552
rect 19430 16496 19486 16532
rect 19798 16632 19854 16688
rect 19616 16346 19672 16348
rect 19696 16346 19752 16348
rect 19776 16346 19832 16348
rect 19856 16346 19912 16348
rect 19616 16294 19642 16346
rect 19642 16294 19672 16346
rect 19696 16294 19706 16346
rect 19706 16294 19752 16346
rect 19776 16294 19822 16346
rect 19822 16294 19832 16346
rect 19856 16294 19886 16346
rect 19886 16294 19912 16346
rect 19616 16292 19672 16294
rect 19696 16292 19752 16294
rect 19776 16292 19832 16294
rect 19856 16292 19912 16294
rect 19246 15544 19302 15600
rect 18878 14764 18880 14784
rect 18880 14764 18932 14784
rect 18932 14764 18934 14784
rect 18878 14728 18934 14764
rect 19616 15258 19672 15260
rect 19696 15258 19752 15260
rect 19776 15258 19832 15260
rect 19856 15258 19912 15260
rect 19616 15206 19642 15258
rect 19642 15206 19672 15258
rect 19696 15206 19706 15258
rect 19706 15206 19752 15258
rect 19776 15206 19822 15258
rect 19822 15206 19832 15258
rect 19856 15206 19886 15258
rect 19886 15206 19912 15258
rect 19616 15204 19672 15206
rect 19696 15204 19752 15206
rect 19776 15204 19832 15206
rect 19856 15204 19912 15206
rect 19154 14320 19210 14376
rect 19062 12280 19118 12336
rect 19890 15000 19946 15056
rect 19614 14320 19670 14376
rect 19616 14170 19672 14172
rect 19696 14170 19752 14172
rect 19776 14170 19832 14172
rect 19856 14170 19912 14172
rect 19616 14118 19642 14170
rect 19642 14118 19672 14170
rect 19696 14118 19706 14170
rect 19706 14118 19752 14170
rect 19776 14118 19822 14170
rect 19822 14118 19832 14170
rect 19856 14118 19886 14170
rect 19886 14118 19912 14170
rect 19616 14116 19672 14118
rect 19696 14116 19752 14118
rect 19776 14116 19832 14118
rect 19856 14116 19912 14118
rect 19430 12824 19486 12880
rect 19616 13082 19672 13084
rect 19696 13082 19752 13084
rect 19776 13082 19832 13084
rect 19856 13082 19912 13084
rect 19616 13030 19642 13082
rect 19642 13030 19672 13082
rect 19696 13030 19706 13082
rect 19706 13030 19752 13082
rect 19776 13030 19822 13082
rect 19822 13030 19832 13082
rect 19856 13030 19886 13082
rect 19886 13030 19912 13082
rect 19616 13028 19672 13030
rect 19696 13028 19752 13030
rect 19776 13028 19832 13030
rect 19856 13028 19912 13030
rect 20626 18264 20682 18320
rect 22098 23568 22154 23624
rect 22006 22888 22062 22944
rect 21822 22208 21878 22264
rect 21638 22092 21694 22128
rect 21638 22072 21640 22092
rect 21640 22072 21692 22092
rect 21692 22072 21694 22092
rect 20902 18808 20958 18864
rect 20258 15680 20314 15736
rect 19430 11636 19432 11656
rect 19432 11636 19484 11656
rect 19484 11636 19486 11656
rect 19430 11600 19486 11636
rect 19430 11192 19486 11248
rect 19616 11994 19672 11996
rect 19696 11994 19752 11996
rect 19776 11994 19832 11996
rect 19856 11994 19912 11996
rect 19616 11942 19642 11994
rect 19642 11942 19672 11994
rect 19696 11942 19706 11994
rect 19706 11942 19752 11994
rect 19776 11942 19822 11994
rect 19822 11942 19832 11994
rect 19856 11942 19886 11994
rect 19886 11942 19912 11994
rect 19616 11940 19672 11942
rect 19696 11940 19752 11942
rect 19776 11940 19832 11942
rect 19856 11940 19912 11942
rect 19616 10906 19672 10908
rect 19696 10906 19752 10908
rect 19776 10906 19832 10908
rect 19856 10906 19912 10908
rect 19616 10854 19642 10906
rect 19642 10854 19672 10906
rect 19696 10854 19706 10906
rect 19706 10854 19752 10906
rect 19776 10854 19822 10906
rect 19822 10854 19832 10906
rect 19856 10854 19886 10906
rect 19886 10854 19912 10906
rect 19616 10852 19672 10854
rect 19696 10852 19752 10854
rect 19776 10852 19832 10854
rect 19856 10852 19912 10854
rect 19338 10648 19394 10704
rect 19614 10648 19670 10704
rect 19430 10512 19486 10568
rect 19338 10240 19394 10296
rect 19154 10104 19210 10160
rect 18970 9560 19026 9616
rect 19246 9560 19302 9616
rect 19798 10668 19854 10704
rect 19798 10648 19800 10668
rect 19800 10648 19852 10668
rect 19852 10648 19854 10668
rect 19706 10412 19708 10432
rect 19708 10412 19760 10432
rect 19760 10412 19762 10432
rect 19706 10376 19762 10412
rect 19246 7384 19302 7440
rect 19616 9818 19672 9820
rect 19696 9818 19752 9820
rect 19776 9818 19832 9820
rect 19856 9818 19912 9820
rect 19616 9766 19642 9818
rect 19642 9766 19672 9818
rect 19696 9766 19706 9818
rect 19706 9766 19752 9818
rect 19776 9766 19822 9818
rect 19822 9766 19832 9818
rect 19856 9766 19886 9818
rect 19886 9766 19912 9818
rect 19616 9764 19672 9766
rect 19696 9764 19752 9766
rect 19776 9764 19832 9766
rect 19856 9764 19912 9766
rect 20166 13796 20222 13832
rect 20166 13776 20168 13796
rect 20168 13776 20220 13796
rect 20220 13776 20222 13796
rect 20166 13504 20222 13560
rect 20166 11056 20222 11112
rect 19616 8730 19672 8732
rect 19696 8730 19752 8732
rect 19776 8730 19832 8732
rect 19856 8730 19912 8732
rect 19616 8678 19642 8730
rect 19642 8678 19672 8730
rect 19696 8678 19706 8730
rect 19706 8678 19752 8730
rect 19776 8678 19822 8730
rect 19822 8678 19832 8730
rect 19856 8678 19886 8730
rect 19886 8678 19912 8730
rect 19616 8676 19672 8678
rect 19696 8676 19752 8678
rect 19776 8676 19832 8678
rect 19856 8676 19912 8678
rect 19706 7828 19708 7848
rect 19708 7828 19760 7848
rect 19760 7828 19762 7848
rect 19706 7792 19762 7828
rect 19616 7642 19672 7644
rect 19696 7642 19752 7644
rect 19776 7642 19832 7644
rect 19856 7642 19912 7644
rect 19616 7590 19642 7642
rect 19642 7590 19672 7642
rect 19696 7590 19706 7642
rect 19706 7590 19752 7642
rect 19776 7590 19822 7642
rect 19822 7590 19832 7642
rect 19856 7590 19886 7642
rect 19886 7590 19912 7642
rect 19616 7588 19672 7590
rect 19696 7588 19752 7590
rect 19776 7588 19832 7590
rect 19856 7588 19912 7590
rect 20258 10920 20314 10976
rect 20442 13232 20498 13288
rect 20810 13776 20866 13832
rect 20902 13368 20958 13424
rect 20534 11600 20590 11656
rect 20442 11056 20498 11112
rect 20350 8880 20406 8936
rect 20166 7384 20222 7440
rect 19338 6976 19394 7032
rect 20074 6840 20130 6896
rect 19616 6554 19672 6556
rect 19696 6554 19752 6556
rect 19776 6554 19832 6556
rect 19856 6554 19912 6556
rect 19616 6502 19642 6554
rect 19642 6502 19672 6554
rect 19696 6502 19706 6554
rect 19706 6502 19752 6554
rect 19776 6502 19822 6554
rect 19822 6502 19832 6554
rect 19856 6502 19886 6554
rect 19886 6502 19912 6554
rect 19616 6500 19672 6502
rect 19696 6500 19752 6502
rect 19776 6500 19832 6502
rect 19856 6500 19912 6502
rect 19982 6296 20038 6352
rect 19616 5466 19672 5468
rect 19696 5466 19752 5468
rect 19776 5466 19832 5468
rect 19856 5466 19912 5468
rect 19616 5414 19642 5466
rect 19642 5414 19672 5466
rect 19696 5414 19706 5466
rect 19706 5414 19752 5466
rect 19776 5414 19822 5466
rect 19822 5414 19832 5466
rect 19856 5414 19886 5466
rect 19886 5414 19912 5466
rect 19616 5412 19672 5414
rect 19696 5412 19752 5414
rect 19776 5412 19832 5414
rect 19856 5412 19912 5414
rect 19616 4378 19672 4380
rect 19696 4378 19752 4380
rect 19776 4378 19832 4380
rect 19856 4378 19912 4380
rect 19616 4326 19642 4378
rect 19642 4326 19672 4378
rect 19696 4326 19706 4378
rect 19706 4326 19752 4378
rect 19776 4326 19822 4378
rect 19822 4326 19832 4378
rect 19856 4326 19886 4378
rect 19886 4326 19912 4378
rect 19616 4324 19672 4326
rect 19696 4324 19752 4326
rect 19776 4324 19832 4326
rect 19856 4324 19912 4326
rect 19890 3612 19892 3632
rect 19892 3612 19944 3632
rect 19944 3612 19946 3632
rect 19890 3576 19946 3612
rect 19616 3290 19672 3292
rect 19696 3290 19752 3292
rect 19776 3290 19832 3292
rect 19856 3290 19912 3292
rect 19616 3238 19642 3290
rect 19642 3238 19672 3290
rect 19696 3238 19706 3290
rect 19706 3238 19752 3290
rect 19776 3238 19822 3290
rect 19822 3238 19832 3290
rect 19856 3238 19886 3290
rect 19886 3238 19912 3290
rect 19616 3236 19672 3238
rect 19696 3236 19752 3238
rect 19776 3236 19832 3238
rect 19856 3236 19912 3238
rect 20166 4936 20222 4992
rect 20810 7828 20812 7848
rect 20812 7828 20864 7848
rect 20864 7828 20866 7848
rect 20810 7792 20866 7828
rect 20442 7268 20498 7304
rect 20442 7248 20444 7268
rect 20444 7248 20496 7268
rect 20496 7248 20498 7268
rect 21178 12688 21234 12744
rect 21178 11192 21234 11248
rect 23110 22208 23166 22264
rect 23110 21548 23166 21584
rect 23110 21528 23112 21548
rect 23112 21528 23164 21548
rect 23164 21528 23166 21548
rect 21454 14456 21510 14512
rect 21362 13776 21418 13832
rect 21178 8200 21234 8256
rect 20534 4256 20590 4312
rect 20258 3032 20314 3088
rect 20534 2896 20590 2952
rect 4688 2202 4744 2204
rect 4768 2202 4824 2204
rect 4848 2202 4904 2204
rect 4928 2202 4984 2204
rect 4688 2150 4714 2202
rect 4714 2150 4744 2202
rect 4768 2150 4778 2202
rect 4778 2150 4824 2202
rect 4848 2150 4894 2202
rect 4894 2150 4904 2202
rect 4928 2150 4958 2202
rect 4958 2150 4984 2202
rect 4688 2148 4744 2150
rect 4768 2148 4824 2150
rect 4848 2148 4904 2150
rect 4928 2148 4984 2150
rect 12152 2202 12208 2204
rect 12232 2202 12288 2204
rect 12312 2202 12368 2204
rect 12392 2202 12448 2204
rect 12152 2150 12178 2202
rect 12178 2150 12208 2202
rect 12232 2150 12242 2202
rect 12242 2150 12288 2202
rect 12312 2150 12358 2202
rect 12358 2150 12368 2202
rect 12392 2150 12422 2202
rect 12422 2150 12448 2202
rect 12152 2148 12208 2150
rect 12232 2148 12288 2150
rect 12312 2148 12368 2150
rect 12392 2148 12448 2150
rect 19616 2202 19672 2204
rect 19696 2202 19752 2204
rect 19776 2202 19832 2204
rect 19856 2202 19912 2204
rect 19616 2150 19642 2202
rect 19642 2150 19672 2202
rect 19696 2150 19706 2202
rect 19706 2150 19752 2202
rect 19776 2150 19822 2202
rect 19822 2150 19832 2202
rect 19856 2150 19886 2202
rect 19886 2150 19912 2202
rect 19616 2148 19672 2150
rect 19696 2148 19752 2150
rect 19776 2148 19832 2150
rect 19856 2148 19912 2150
rect 21362 5616 21418 5672
rect 22742 20868 22798 20904
rect 22742 20848 22744 20868
rect 22744 20848 22796 20868
rect 22796 20848 22798 20868
rect 21914 16632 21970 16688
rect 23018 20168 23074 20224
rect 23110 19488 23166 19544
rect 21914 10512 21970 10568
rect 22098 7284 22100 7304
rect 22100 7284 22152 7304
rect 22152 7284 22154 7304
rect 22098 7248 22154 7284
rect 21362 3052 21418 3088
rect 21362 3032 21364 3052
rect 21364 3032 21416 3052
rect 21416 3032 21418 3052
rect 22650 14476 22706 14512
rect 22650 14456 22652 14476
rect 22652 14456 22704 14476
rect 22704 14456 22706 14476
rect 22374 12688 22430 12744
rect 23570 17584 23626 17640
rect 21914 2216 21970 2272
rect 22006 856 22062 912
rect 23294 7520 23350 7576
rect 23294 6976 23350 7032
rect 23018 1536 23074 1592
rect 23570 312 23626 368
<< metal3 >>
rect 21817 24306 21883 24309
rect 23800 24306 24600 24336
rect 21817 24304 24600 24306
rect 21817 24248 21822 24304
rect 21878 24248 24600 24304
rect 21817 24246 24600 24248
rect 21817 24243 21883 24246
rect 23800 24216 24600 24246
rect 22093 23626 22159 23629
rect 23800 23626 24600 23656
rect 22093 23624 24600 23626
rect 22093 23568 22098 23624
rect 22154 23568 24600 23624
rect 22093 23566 24600 23568
rect 22093 23563 22159 23566
rect 23800 23536 24600 23566
rect 22001 22946 22067 22949
rect 23800 22946 24600 22976
rect 22001 22944 24600 22946
rect 22001 22888 22006 22944
rect 22062 22888 24600 22944
rect 22001 22886 24600 22888
rect 22001 22883 22067 22886
rect 23800 22856 24600 22886
rect 8408 22336 8728 22337
rect 8408 22272 8416 22336
rect 8480 22272 8496 22336
rect 8560 22272 8576 22336
rect 8640 22272 8656 22336
rect 8720 22272 8728 22336
rect 8408 22271 8728 22272
rect 15872 22336 16192 22337
rect 15872 22272 15880 22336
rect 15944 22272 15960 22336
rect 16024 22272 16040 22336
rect 16104 22272 16120 22336
rect 16184 22272 16192 22336
rect 15872 22271 16192 22272
rect 21817 22266 21883 22269
rect 21774 22264 21883 22266
rect 21774 22208 21822 22264
rect 21878 22208 21883 22264
rect 21774 22203 21883 22208
rect 23105 22266 23171 22269
rect 23800 22266 24600 22296
rect 23105 22264 24600 22266
rect 23105 22208 23110 22264
rect 23166 22208 24600 22264
rect 23105 22206 24600 22208
rect 23105 22203 23171 22206
rect 10041 22130 10107 22133
rect 11697 22130 11763 22133
rect 10041 22128 11763 22130
rect 10041 22072 10046 22128
rect 10102 22072 11702 22128
rect 11758 22072 11763 22128
rect 10041 22070 11763 22072
rect 10041 22067 10107 22070
rect 11697 22067 11763 22070
rect 21633 22130 21699 22133
rect 21774 22130 21834 22203
rect 23800 22176 24600 22206
rect 21633 22128 21834 22130
rect 21633 22072 21638 22128
rect 21694 22072 21834 22128
rect 21633 22070 21834 22072
rect 21633 22067 21699 22070
rect 3693 21994 3759 21997
rect 8753 21994 8819 21997
rect 3693 21992 8819 21994
rect 3693 21936 3698 21992
rect 3754 21936 8758 21992
rect 8814 21936 8819 21992
rect 3693 21934 8819 21936
rect 3693 21931 3759 21934
rect 8753 21931 8819 21934
rect 11237 21994 11303 21997
rect 12801 21994 12867 21997
rect 11237 21992 12867 21994
rect 11237 21936 11242 21992
rect 11298 21936 12806 21992
rect 12862 21936 12867 21992
rect 11237 21934 12867 21936
rect 11237 21931 11303 21934
rect 12801 21931 12867 21934
rect 4676 21792 4996 21793
rect 4676 21728 4684 21792
rect 4748 21728 4764 21792
rect 4828 21728 4844 21792
rect 4908 21728 4924 21792
rect 4988 21728 4996 21792
rect 4676 21727 4996 21728
rect 12140 21792 12460 21793
rect 12140 21728 12148 21792
rect 12212 21728 12228 21792
rect 12292 21728 12308 21792
rect 12372 21728 12388 21792
rect 12452 21728 12460 21792
rect 12140 21727 12460 21728
rect 19604 21792 19924 21793
rect 19604 21728 19612 21792
rect 19676 21728 19692 21792
rect 19756 21728 19772 21792
rect 19836 21728 19852 21792
rect 19916 21728 19924 21792
rect 19604 21727 19924 21728
rect 2497 21586 2563 21589
rect 8569 21586 8635 21589
rect 2497 21584 8635 21586
rect 2497 21528 2502 21584
rect 2558 21528 8574 21584
rect 8630 21528 8635 21584
rect 2497 21526 8635 21528
rect 2497 21523 2563 21526
rect 8569 21523 8635 21526
rect 10961 21586 11027 21589
rect 11697 21586 11763 21589
rect 10961 21584 11763 21586
rect 10961 21528 10966 21584
rect 11022 21528 11702 21584
rect 11758 21528 11763 21584
rect 10961 21526 11763 21528
rect 10961 21523 11027 21526
rect 11697 21523 11763 21526
rect 12341 21586 12407 21589
rect 13537 21586 13603 21589
rect 19149 21586 19215 21589
rect 12341 21584 19215 21586
rect 12341 21528 12346 21584
rect 12402 21528 13542 21584
rect 13598 21528 19154 21584
rect 19210 21528 19215 21584
rect 12341 21526 19215 21528
rect 12341 21523 12407 21526
rect 13537 21523 13603 21526
rect 19149 21523 19215 21526
rect 23105 21586 23171 21589
rect 23800 21586 24600 21616
rect 23105 21584 24600 21586
rect 23105 21528 23110 21584
rect 23166 21528 24600 21584
rect 23105 21526 24600 21528
rect 23105 21523 23171 21526
rect 23800 21496 24600 21526
rect 0 21450 800 21480
rect 1577 21450 1643 21453
rect 0 21448 1643 21450
rect 0 21392 1582 21448
rect 1638 21392 1643 21448
rect 0 21390 1643 21392
rect 0 21360 800 21390
rect 1577 21387 1643 21390
rect 7557 21450 7623 21453
rect 8385 21450 8451 21453
rect 7557 21448 8451 21450
rect 7557 21392 7562 21448
rect 7618 21392 8390 21448
rect 8446 21392 8451 21448
rect 7557 21390 8451 21392
rect 7557 21387 7623 21390
rect 8385 21387 8451 21390
rect 10685 21450 10751 21453
rect 11237 21450 11303 21453
rect 18045 21450 18111 21453
rect 10685 21448 18111 21450
rect 10685 21392 10690 21448
rect 10746 21392 11242 21448
rect 11298 21392 18050 21448
rect 18106 21392 18111 21448
rect 10685 21390 18111 21392
rect 10685 21387 10751 21390
rect 11237 21387 11303 21390
rect 18045 21387 18111 21390
rect 10409 21314 10475 21317
rect 14457 21314 14523 21317
rect 10409 21312 14523 21314
rect 10409 21256 10414 21312
rect 10470 21256 14462 21312
rect 14518 21256 14523 21312
rect 10409 21254 14523 21256
rect 10409 21251 10475 21254
rect 14457 21251 14523 21254
rect 8408 21248 8728 21249
rect 8408 21184 8416 21248
rect 8480 21184 8496 21248
rect 8560 21184 8576 21248
rect 8640 21184 8656 21248
rect 8720 21184 8728 21248
rect 8408 21183 8728 21184
rect 15872 21248 16192 21249
rect 15872 21184 15880 21248
rect 15944 21184 15960 21248
rect 16024 21184 16040 21248
rect 16104 21184 16120 21248
rect 16184 21184 16192 21248
rect 15872 21183 16192 21184
rect 12341 21042 12407 21045
rect 13353 21042 13419 21045
rect 12341 21040 13419 21042
rect 12341 20984 12346 21040
rect 12402 20984 13358 21040
rect 13414 20984 13419 21040
rect 12341 20982 13419 20984
rect 12341 20979 12407 20982
rect 13353 20979 13419 20982
rect 14181 21042 14247 21045
rect 17309 21042 17375 21045
rect 14181 21040 17375 21042
rect 14181 20984 14186 21040
rect 14242 20984 17314 21040
rect 17370 20984 17375 21040
rect 14181 20982 17375 20984
rect 14181 20979 14247 20982
rect 17309 20979 17375 20982
rect 1669 20906 1735 20909
rect 8477 20906 8543 20909
rect 1669 20904 8543 20906
rect 1669 20848 1674 20904
rect 1730 20848 8482 20904
rect 8538 20848 8543 20904
rect 1669 20846 8543 20848
rect 1669 20843 1735 20846
rect 8477 20843 8543 20846
rect 22737 20906 22803 20909
rect 23800 20906 24600 20936
rect 22737 20904 24600 20906
rect 22737 20848 22742 20904
rect 22798 20848 24600 20904
rect 22737 20846 24600 20848
rect 22737 20843 22803 20846
rect 23800 20816 24600 20846
rect 4676 20704 4996 20705
rect 4676 20640 4684 20704
rect 4748 20640 4764 20704
rect 4828 20640 4844 20704
rect 4908 20640 4924 20704
rect 4988 20640 4996 20704
rect 4676 20639 4996 20640
rect 12140 20704 12460 20705
rect 12140 20640 12148 20704
rect 12212 20640 12228 20704
rect 12292 20640 12308 20704
rect 12372 20640 12388 20704
rect 12452 20640 12460 20704
rect 12140 20639 12460 20640
rect 19604 20704 19924 20705
rect 19604 20640 19612 20704
rect 19676 20640 19692 20704
rect 19756 20640 19772 20704
rect 19836 20640 19852 20704
rect 19916 20640 19924 20704
rect 19604 20639 19924 20640
rect 23013 20226 23079 20229
rect 23800 20226 24600 20256
rect 23013 20224 24600 20226
rect 23013 20168 23018 20224
rect 23074 20168 24600 20224
rect 23013 20166 24600 20168
rect 23013 20163 23079 20166
rect 8408 20160 8728 20161
rect 8408 20096 8416 20160
rect 8480 20096 8496 20160
rect 8560 20096 8576 20160
rect 8640 20096 8656 20160
rect 8720 20096 8728 20160
rect 8408 20095 8728 20096
rect 15872 20160 16192 20161
rect 15872 20096 15880 20160
rect 15944 20096 15960 20160
rect 16024 20096 16040 20160
rect 16104 20096 16120 20160
rect 16184 20096 16192 20160
rect 23800 20136 24600 20166
rect 15872 20095 16192 20096
rect 4676 19616 4996 19617
rect 4676 19552 4684 19616
rect 4748 19552 4764 19616
rect 4828 19552 4844 19616
rect 4908 19552 4924 19616
rect 4988 19552 4996 19616
rect 4676 19551 4996 19552
rect 12140 19616 12460 19617
rect 12140 19552 12148 19616
rect 12212 19552 12228 19616
rect 12292 19552 12308 19616
rect 12372 19552 12388 19616
rect 12452 19552 12460 19616
rect 12140 19551 12460 19552
rect 19604 19616 19924 19617
rect 19604 19552 19612 19616
rect 19676 19552 19692 19616
rect 19756 19552 19772 19616
rect 19836 19552 19852 19616
rect 19916 19552 19924 19616
rect 19604 19551 19924 19552
rect 23105 19546 23171 19549
rect 23800 19546 24600 19576
rect 23105 19544 24600 19546
rect 23105 19488 23110 19544
rect 23166 19488 24600 19544
rect 23105 19486 24600 19488
rect 23105 19483 23171 19486
rect 23800 19456 24600 19486
rect 10685 19410 10751 19413
rect 19241 19410 19307 19413
rect 10685 19408 19307 19410
rect 10685 19352 10690 19408
rect 10746 19352 19246 19408
rect 19302 19352 19307 19408
rect 10685 19350 19307 19352
rect 10685 19347 10751 19350
rect 19241 19347 19307 19350
rect 11697 19274 11763 19277
rect 15469 19274 15535 19277
rect 11697 19272 15535 19274
rect 11697 19216 11702 19272
rect 11758 19216 15474 19272
rect 15530 19216 15535 19272
rect 11697 19214 15535 19216
rect 11697 19211 11763 19214
rect 15469 19211 15535 19214
rect 8408 19072 8728 19073
rect 8408 19008 8416 19072
rect 8480 19008 8496 19072
rect 8560 19008 8576 19072
rect 8640 19008 8656 19072
rect 8720 19008 8728 19072
rect 8408 19007 8728 19008
rect 15872 19072 16192 19073
rect 15872 19008 15880 19072
rect 15944 19008 15960 19072
rect 16024 19008 16040 19072
rect 16104 19008 16120 19072
rect 16184 19008 16192 19072
rect 15872 19007 16192 19008
rect 20897 18866 20963 18869
rect 23800 18866 24600 18896
rect 20897 18864 24600 18866
rect 20897 18808 20902 18864
rect 20958 18808 24600 18864
rect 20897 18806 24600 18808
rect 20897 18803 20963 18806
rect 23800 18776 24600 18806
rect 4676 18528 4996 18529
rect 4676 18464 4684 18528
rect 4748 18464 4764 18528
rect 4828 18464 4844 18528
rect 4908 18464 4924 18528
rect 4988 18464 4996 18528
rect 4676 18463 4996 18464
rect 12140 18528 12460 18529
rect 12140 18464 12148 18528
rect 12212 18464 12228 18528
rect 12292 18464 12308 18528
rect 12372 18464 12388 18528
rect 12452 18464 12460 18528
rect 12140 18463 12460 18464
rect 19604 18528 19924 18529
rect 19604 18464 19612 18528
rect 19676 18464 19692 18528
rect 19756 18464 19772 18528
rect 19836 18464 19852 18528
rect 19916 18464 19924 18528
rect 19604 18463 19924 18464
rect 20621 18322 20687 18325
rect 23800 18322 24600 18352
rect 20621 18320 24600 18322
rect 20621 18264 20626 18320
rect 20682 18264 24600 18320
rect 20621 18262 24600 18264
rect 20621 18259 20687 18262
rect 23800 18232 24600 18262
rect 8408 17984 8728 17985
rect 8408 17920 8416 17984
rect 8480 17920 8496 17984
rect 8560 17920 8576 17984
rect 8640 17920 8656 17984
rect 8720 17920 8728 17984
rect 8408 17919 8728 17920
rect 15872 17984 16192 17985
rect 15872 17920 15880 17984
rect 15944 17920 15960 17984
rect 16024 17920 16040 17984
rect 16104 17920 16120 17984
rect 16184 17920 16192 17984
rect 15872 17919 16192 17920
rect 23565 17642 23631 17645
rect 23800 17642 24600 17672
rect 23565 17640 24600 17642
rect 23565 17584 23570 17640
rect 23626 17584 24600 17640
rect 23565 17582 24600 17584
rect 23565 17579 23631 17582
rect 23800 17552 24600 17582
rect 4676 17440 4996 17441
rect 4676 17376 4684 17440
rect 4748 17376 4764 17440
rect 4828 17376 4844 17440
rect 4908 17376 4924 17440
rect 4988 17376 4996 17440
rect 4676 17375 4996 17376
rect 12140 17440 12460 17441
rect 12140 17376 12148 17440
rect 12212 17376 12228 17440
rect 12292 17376 12308 17440
rect 12372 17376 12388 17440
rect 12452 17376 12460 17440
rect 12140 17375 12460 17376
rect 19604 17440 19924 17441
rect 19604 17376 19612 17440
rect 19676 17376 19692 17440
rect 19756 17376 19772 17440
rect 19836 17376 19852 17440
rect 19916 17376 19924 17440
rect 19604 17375 19924 17376
rect 19517 16962 19583 16965
rect 23800 16962 24600 16992
rect 19517 16960 24600 16962
rect 19517 16904 19522 16960
rect 19578 16904 24600 16960
rect 19517 16902 24600 16904
rect 19517 16899 19583 16902
rect 8408 16896 8728 16897
rect 8408 16832 8416 16896
rect 8480 16832 8496 16896
rect 8560 16832 8576 16896
rect 8640 16832 8656 16896
rect 8720 16832 8728 16896
rect 8408 16831 8728 16832
rect 15872 16896 16192 16897
rect 15872 16832 15880 16896
rect 15944 16832 15960 16896
rect 16024 16832 16040 16896
rect 16104 16832 16120 16896
rect 16184 16832 16192 16896
rect 23800 16872 24600 16902
rect 15872 16831 16192 16832
rect 15469 16690 15535 16693
rect 18045 16690 18111 16693
rect 15469 16688 18111 16690
rect 15469 16632 15474 16688
rect 15530 16632 18050 16688
rect 18106 16632 18111 16688
rect 15469 16630 18111 16632
rect 15469 16627 15535 16630
rect 18045 16627 18111 16630
rect 19793 16690 19859 16693
rect 21909 16690 21975 16693
rect 19793 16688 21975 16690
rect 19793 16632 19798 16688
rect 19854 16632 21914 16688
rect 21970 16632 21975 16688
rect 19793 16630 21975 16632
rect 19793 16627 19859 16630
rect 21909 16627 21975 16630
rect 19425 16554 19491 16557
rect 19425 16552 22110 16554
rect 19425 16496 19430 16552
rect 19486 16496 22110 16552
rect 19425 16494 22110 16496
rect 19425 16491 19491 16494
rect 4676 16352 4996 16353
rect 4676 16288 4684 16352
rect 4748 16288 4764 16352
rect 4828 16288 4844 16352
rect 4908 16288 4924 16352
rect 4988 16288 4996 16352
rect 4676 16287 4996 16288
rect 12140 16352 12460 16353
rect 12140 16288 12148 16352
rect 12212 16288 12228 16352
rect 12292 16288 12308 16352
rect 12372 16288 12388 16352
rect 12452 16288 12460 16352
rect 12140 16287 12460 16288
rect 19604 16352 19924 16353
rect 19604 16288 19612 16352
rect 19676 16288 19692 16352
rect 19756 16288 19772 16352
rect 19836 16288 19852 16352
rect 19916 16288 19924 16352
rect 19604 16287 19924 16288
rect 22050 16282 22110 16494
rect 23800 16282 24600 16312
rect 22050 16222 24600 16282
rect 23800 16192 24600 16222
rect 8408 15808 8728 15809
rect 8408 15744 8416 15808
rect 8480 15744 8496 15808
rect 8560 15744 8576 15808
rect 8640 15744 8656 15808
rect 8720 15744 8728 15808
rect 8408 15743 8728 15744
rect 15872 15808 16192 15809
rect 15872 15744 15880 15808
rect 15944 15744 15960 15808
rect 16024 15744 16040 15808
rect 16104 15744 16120 15808
rect 16184 15744 16192 15808
rect 15872 15743 16192 15744
rect 20110 15676 20116 15740
rect 20180 15738 20186 15740
rect 20253 15738 20319 15741
rect 20180 15736 20319 15738
rect 20180 15680 20258 15736
rect 20314 15680 20319 15736
rect 20180 15678 20319 15680
rect 20180 15676 20186 15678
rect 20253 15675 20319 15678
rect 19241 15602 19307 15605
rect 23800 15602 24600 15632
rect 19241 15600 24600 15602
rect 19241 15544 19246 15600
rect 19302 15544 24600 15600
rect 19241 15542 24600 15544
rect 19241 15539 19307 15542
rect 23800 15512 24600 15542
rect 0 15330 800 15360
rect 1485 15330 1551 15333
rect 0 15328 1551 15330
rect 0 15272 1490 15328
rect 1546 15272 1551 15328
rect 0 15270 1551 15272
rect 0 15240 800 15270
rect 1485 15267 1551 15270
rect 4676 15264 4996 15265
rect 4676 15200 4684 15264
rect 4748 15200 4764 15264
rect 4828 15200 4844 15264
rect 4908 15200 4924 15264
rect 4988 15200 4996 15264
rect 4676 15199 4996 15200
rect 12140 15264 12460 15265
rect 12140 15200 12148 15264
rect 12212 15200 12228 15264
rect 12292 15200 12308 15264
rect 12372 15200 12388 15264
rect 12452 15200 12460 15264
rect 12140 15199 12460 15200
rect 19604 15264 19924 15265
rect 19604 15200 19612 15264
rect 19676 15200 19692 15264
rect 19756 15200 19772 15264
rect 19836 15200 19852 15264
rect 19916 15200 19924 15264
rect 19604 15199 19924 15200
rect 9857 15194 9923 15197
rect 11145 15194 11211 15197
rect 9857 15192 11211 15194
rect 9857 15136 9862 15192
rect 9918 15136 11150 15192
rect 11206 15136 11211 15192
rect 9857 15134 11211 15136
rect 9857 15131 9923 15134
rect 11145 15131 11211 15134
rect 17769 15058 17835 15061
rect 19885 15058 19951 15061
rect 17769 15056 19951 15058
rect 17769 15000 17774 15056
rect 17830 15000 19890 15056
rect 19946 15000 19951 15056
rect 17769 14998 19951 15000
rect 17769 14995 17835 14998
rect 19885 14995 19951 14998
rect 17401 14922 17467 14925
rect 23800 14922 24600 14952
rect 17401 14920 24600 14922
rect 17401 14864 17406 14920
rect 17462 14864 24600 14920
rect 17401 14862 24600 14864
rect 17401 14859 17467 14862
rect 23800 14832 24600 14862
rect 18045 14786 18111 14789
rect 18873 14786 18939 14789
rect 18045 14784 18939 14786
rect 18045 14728 18050 14784
rect 18106 14728 18878 14784
rect 18934 14728 18939 14784
rect 18045 14726 18939 14728
rect 18045 14723 18111 14726
rect 18873 14723 18939 14726
rect 8408 14720 8728 14721
rect 8408 14656 8416 14720
rect 8480 14656 8496 14720
rect 8560 14656 8576 14720
rect 8640 14656 8656 14720
rect 8720 14656 8728 14720
rect 8408 14655 8728 14656
rect 15872 14720 16192 14721
rect 15872 14656 15880 14720
rect 15944 14656 15960 14720
rect 16024 14656 16040 14720
rect 16104 14656 16120 14720
rect 16184 14656 16192 14720
rect 15872 14655 16192 14656
rect 10961 14514 11027 14517
rect 18413 14514 18479 14517
rect 10961 14512 18479 14514
rect 10961 14456 10966 14512
rect 11022 14456 18418 14512
rect 18474 14456 18479 14512
rect 10961 14454 18479 14456
rect 10961 14451 11027 14454
rect 18413 14451 18479 14454
rect 21449 14514 21515 14517
rect 22645 14514 22711 14517
rect 21449 14512 22711 14514
rect 21449 14456 21454 14512
rect 21510 14456 22650 14512
rect 22706 14456 22711 14512
rect 21449 14454 22711 14456
rect 21449 14451 21515 14454
rect 22645 14451 22711 14454
rect 16665 14378 16731 14381
rect 19149 14378 19215 14381
rect 16665 14376 19215 14378
rect 16665 14320 16670 14376
rect 16726 14320 19154 14376
rect 19210 14320 19215 14376
rect 16665 14318 19215 14320
rect 16665 14315 16731 14318
rect 19149 14315 19215 14318
rect 19609 14378 19675 14381
rect 19609 14376 22110 14378
rect 19609 14320 19614 14376
rect 19670 14320 22110 14376
rect 19609 14318 22110 14320
rect 19609 14315 19675 14318
rect 22050 14242 22110 14318
rect 23800 14242 24600 14272
rect 22050 14182 24600 14242
rect 4676 14176 4996 14177
rect 4676 14112 4684 14176
rect 4748 14112 4764 14176
rect 4828 14112 4844 14176
rect 4908 14112 4924 14176
rect 4988 14112 4996 14176
rect 4676 14111 4996 14112
rect 12140 14176 12460 14177
rect 12140 14112 12148 14176
rect 12212 14112 12228 14176
rect 12292 14112 12308 14176
rect 12372 14112 12388 14176
rect 12452 14112 12460 14176
rect 12140 14111 12460 14112
rect 19604 14176 19924 14177
rect 19604 14112 19612 14176
rect 19676 14112 19692 14176
rect 19756 14112 19772 14176
rect 19836 14112 19852 14176
rect 19916 14112 19924 14176
rect 23800 14152 24600 14182
rect 19604 14111 19924 14112
rect 10777 13970 10843 13973
rect 13077 13970 13143 13973
rect 10777 13968 13143 13970
rect 10777 13912 10782 13968
rect 10838 13912 13082 13968
rect 13138 13912 13143 13968
rect 10777 13910 13143 13912
rect 10777 13907 10843 13910
rect 13077 13907 13143 13910
rect 20161 13834 20227 13837
rect 20805 13834 20871 13837
rect 21357 13834 21423 13837
rect 20161 13832 21423 13834
rect 20161 13776 20166 13832
rect 20222 13776 20810 13832
rect 20866 13776 21362 13832
rect 21418 13776 21423 13832
rect 20161 13774 21423 13776
rect 20161 13771 20227 13774
rect 20805 13771 20871 13774
rect 21357 13771 21423 13774
rect 8408 13632 8728 13633
rect 8408 13568 8416 13632
rect 8480 13568 8496 13632
rect 8560 13568 8576 13632
rect 8640 13568 8656 13632
rect 8720 13568 8728 13632
rect 8408 13567 8728 13568
rect 15872 13632 16192 13633
rect 15872 13568 15880 13632
rect 15944 13568 15960 13632
rect 16024 13568 16040 13632
rect 16104 13568 16120 13632
rect 16184 13568 16192 13632
rect 15872 13567 16192 13568
rect 20161 13562 20227 13565
rect 23800 13562 24600 13592
rect 20161 13560 24600 13562
rect 20161 13504 20166 13560
rect 20222 13504 24600 13560
rect 20161 13502 24600 13504
rect 20161 13499 20227 13502
rect 23800 13472 24600 13502
rect 9673 13426 9739 13429
rect 20897 13426 20963 13429
rect 9673 13424 20963 13426
rect 9673 13368 9678 13424
rect 9734 13368 20902 13424
rect 20958 13368 20963 13424
rect 9673 13366 20963 13368
rect 9673 13363 9739 13366
rect 20897 13363 20963 13366
rect 15193 13290 15259 13293
rect 18321 13290 18387 13293
rect 15193 13288 18387 13290
rect 15193 13232 15198 13288
rect 15254 13232 18326 13288
rect 18382 13232 18387 13288
rect 15193 13230 18387 13232
rect 15193 13227 15259 13230
rect 18321 13227 18387 13230
rect 20437 13292 20503 13293
rect 20437 13288 20484 13292
rect 20548 13290 20554 13292
rect 20437 13232 20442 13288
rect 20437 13228 20484 13232
rect 20548 13230 20594 13290
rect 20548 13228 20554 13230
rect 20437 13227 20503 13228
rect 4676 13088 4996 13089
rect 4676 13024 4684 13088
rect 4748 13024 4764 13088
rect 4828 13024 4844 13088
rect 4908 13024 4924 13088
rect 4988 13024 4996 13088
rect 4676 13023 4996 13024
rect 12140 13088 12460 13089
rect 12140 13024 12148 13088
rect 12212 13024 12228 13088
rect 12292 13024 12308 13088
rect 12372 13024 12388 13088
rect 12452 13024 12460 13088
rect 12140 13023 12460 13024
rect 19604 13088 19924 13089
rect 19604 13024 19612 13088
rect 19676 13024 19692 13088
rect 19756 13024 19772 13088
rect 19836 13024 19852 13088
rect 19916 13024 19924 13088
rect 19604 13023 19924 13024
rect 19425 12882 19491 12885
rect 23800 12882 24600 12912
rect 19425 12880 24600 12882
rect 19425 12824 19430 12880
rect 19486 12824 24600 12880
rect 19425 12822 24600 12824
rect 19425 12819 19491 12822
rect 23800 12792 24600 12822
rect 15929 12746 15995 12749
rect 17125 12746 17191 12749
rect 15929 12744 17191 12746
rect 15929 12688 15934 12744
rect 15990 12688 17130 12744
rect 17186 12688 17191 12744
rect 15929 12686 17191 12688
rect 15929 12683 15995 12686
rect 17125 12683 17191 12686
rect 21173 12746 21239 12749
rect 22369 12746 22435 12749
rect 21173 12744 22435 12746
rect 21173 12688 21178 12744
rect 21234 12688 22374 12744
rect 22430 12688 22435 12744
rect 21173 12686 22435 12688
rect 21173 12683 21239 12686
rect 22369 12683 22435 12686
rect 8408 12544 8728 12545
rect 8408 12480 8416 12544
rect 8480 12480 8496 12544
rect 8560 12480 8576 12544
rect 8640 12480 8656 12544
rect 8720 12480 8728 12544
rect 8408 12479 8728 12480
rect 15872 12544 16192 12545
rect 15872 12480 15880 12544
rect 15944 12480 15960 12544
rect 16024 12480 16040 12544
rect 16104 12480 16120 12544
rect 16184 12480 16192 12544
rect 15872 12479 16192 12480
rect 15009 12338 15075 12341
rect 17217 12338 17283 12341
rect 15009 12336 17283 12338
rect 15009 12280 15014 12336
rect 15070 12280 17222 12336
rect 17278 12280 17283 12336
rect 15009 12278 17283 12280
rect 15009 12275 15075 12278
rect 17217 12275 17283 12278
rect 19057 12338 19123 12341
rect 23800 12338 24600 12368
rect 19057 12336 24600 12338
rect 19057 12280 19062 12336
rect 19118 12280 24600 12336
rect 19057 12278 24600 12280
rect 19057 12275 19123 12278
rect 23800 12248 24600 12278
rect 10501 12202 10567 12205
rect 12249 12202 12315 12205
rect 10501 12200 12315 12202
rect 10501 12144 10506 12200
rect 10562 12144 12254 12200
rect 12310 12144 12315 12200
rect 10501 12142 12315 12144
rect 10501 12139 10567 12142
rect 12249 12139 12315 12142
rect 4676 12000 4996 12001
rect 4676 11936 4684 12000
rect 4748 11936 4764 12000
rect 4828 11936 4844 12000
rect 4908 11936 4924 12000
rect 4988 11936 4996 12000
rect 4676 11935 4996 11936
rect 12140 12000 12460 12001
rect 12140 11936 12148 12000
rect 12212 11936 12228 12000
rect 12292 11936 12308 12000
rect 12372 11936 12388 12000
rect 12452 11936 12460 12000
rect 12140 11935 12460 11936
rect 19604 12000 19924 12001
rect 19604 11936 19612 12000
rect 19676 11936 19692 12000
rect 19756 11936 19772 12000
rect 19836 11936 19852 12000
rect 19916 11936 19924 12000
rect 19604 11935 19924 11936
rect 17493 11658 17559 11661
rect 19425 11658 19491 11661
rect 17493 11656 19491 11658
rect 17493 11600 17498 11656
rect 17554 11600 19430 11656
rect 19486 11600 19491 11656
rect 17493 11598 19491 11600
rect 17493 11595 17559 11598
rect 19425 11595 19491 11598
rect 20529 11658 20595 11661
rect 23800 11658 24600 11688
rect 20529 11656 24600 11658
rect 20529 11600 20534 11656
rect 20590 11600 24600 11656
rect 20529 11598 24600 11600
rect 20529 11595 20595 11598
rect 23800 11568 24600 11598
rect 8408 11456 8728 11457
rect 8408 11392 8416 11456
rect 8480 11392 8496 11456
rect 8560 11392 8576 11456
rect 8640 11392 8656 11456
rect 8720 11392 8728 11456
rect 8408 11391 8728 11392
rect 15872 11456 16192 11457
rect 15872 11392 15880 11456
rect 15944 11392 15960 11456
rect 16024 11392 16040 11456
rect 16104 11392 16120 11456
rect 16184 11392 16192 11456
rect 15872 11391 16192 11392
rect 19425 11250 19491 11253
rect 21173 11250 21239 11253
rect 19425 11248 21239 11250
rect 19425 11192 19430 11248
rect 19486 11192 21178 11248
rect 21234 11192 21239 11248
rect 19425 11190 21239 11192
rect 19425 11187 19491 11190
rect 21173 11187 21239 11190
rect 20161 11116 20227 11117
rect 20110 11114 20116 11116
rect 20070 11054 20116 11114
rect 20180 11112 20227 11116
rect 20437 11116 20503 11117
rect 20437 11114 20484 11116
rect 20222 11056 20227 11112
rect 20110 11052 20116 11054
rect 20180 11052 20227 11056
rect 20392 11112 20484 11114
rect 20392 11056 20442 11112
rect 20392 11054 20484 11056
rect 20161 11051 20227 11052
rect 20437 11052 20484 11054
rect 20548 11052 20554 11116
rect 20437 11051 20503 11052
rect 20253 10978 20319 10981
rect 23800 10978 24600 11008
rect 20253 10976 24600 10978
rect 20253 10920 20258 10976
rect 20314 10920 24600 10976
rect 20253 10918 24600 10920
rect 20253 10915 20319 10918
rect 4676 10912 4996 10913
rect 4676 10848 4684 10912
rect 4748 10848 4764 10912
rect 4828 10848 4844 10912
rect 4908 10848 4924 10912
rect 4988 10848 4996 10912
rect 4676 10847 4996 10848
rect 12140 10912 12460 10913
rect 12140 10848 12148 10912
rect 12212 10848 12228 10912
rect 12292 10848 12308 10912
rect 12372 10848 12388 10912
rect 12452 10848 12460 10912
rect 12140 10847 12460 10848
rect 19604 10912 19924 10913
rect 19604 10848 19612 10912
rect 19676 10848 19692 10912
rect 19756 10848 19772 10912
rect 19836 10848 19852 10912
rect 19916 10848 19924 10912
rect 23800 10888 24600 10918
rect 19604 10847 19924 10848
rect 19333 10706 19399 10709
rect 19198 10704 19399 10706
rect 19198 10648 19338 10704
rect 19394 10648 19399 10704
rect 19198 10646 19399 10648
rect 16481 10434 16547 10437
rect 18045 10434 18111 10437
rect 16481 10432 18111 10434
rect 16481 10376 16486 10432
rect 16542 10376 18050 10432
rect 18106 10376 18111 10432
rect 16481 10374 18111 10376
rect 16481 10371 16547 10374
rect 18045 10371 18111 10374
rect 18689 10434 18755 10437
rect 19198 10434 19258 10646
rect 19333 10643 19399 10646
rect 19609 10706 19675 10709
rect 19793 10706 19859 10709
rect 19609 10704 19859 10706
rect 19609 10648 19614 10704
rect 19670 10648 19798 10704
rect 19854 10648 19859 10704
rect 19609 10646 19859 10648
rect 19609 10643 19675 10646
rect 19793 10643 19859 10646
rect 19425 10570 19491 10573
rect 21909 10570 21975 10573
rect 19425 10568 21975 10570
rect 19425 10512 19430 10568
rect 19486 10512 21914 10568
rect 21970 10512 21975 10568
rect 19425 10510 21975 10512
rect 19425 10507 19491 10510
rect 21909 10507 21975 10510
rect 19701 10434 19767 10437
rect 18689 10432 19767 10434
rect 18689 10376 18694 10432
rect 18750 10376 19706 10432
rect 19762 10376 19767 10432
rect 18689 10374 19767 10376
rect 18689 10371 18755 10374
rect 19701 10371 19767 10374
rect 8408 10368 8728 10369
rect 8408 10304 8416 10368
rect 8480 10304 8496 10368
rect 8560 10304 8576 10368
rect 8640 10304 8656 10368
rect 8720 10304 8728 10368
rect 8408 10303 8728 10304
rect 15872 10368 16192 10369
rect 15872 10304 15880 10368
rect 15944 10304 15960 10368
rect 16024 10304 16040 10368
rect 16104 10304 16120 10368
rect 16184 10304 16192 10368
rect 15872 10303 16192 10304
rect 19333 10298 19399 10301
rect 23800 10298 24600 10328
rect 19333 10296 24600 10298
rect 19333 10240 19338 10296
rect 19394 10240 24600 10296
rect 19333 10238 24600 10240
rect 19333 10235 19399 10238
rect 23800 10208 24600 10238
rect 17401 10162 17467 10165
rect 19149 10162 19215 10165
rect 17401 10160 19215 10162
rect 17401 10104 17406 10160
rect 17462 10104 19154 10160
rect 19210 10104 19215 10160
rect 17401 10102 19215 10104
rect 17401 10099 17467 10102
rect 19149 10099 19215 10102
rect 4676 9824 4996 9825
rect 4676 9760 4684 9824
rect 4748 9760 4764 9824
rect 4828 9760 4844 9824
rect 4908 9760 4924 9824
rect 4988 9760 4996 9824
rect 4676 9759 4996 9760
rect 12140 9824 12460 9825
rect 12140 9760 12148 9824
rect 12212 9760 12228 9824
rect 12292 9760 12308 9824
rect 12372 9760 12388 9824
rect 12452 9760 12460 9824
rect 12140 9759 12460 9760
rect 19604 9824 19924 9825
rect 19604 9760 19612 9824
rect 19676 9760 19692 9824
rect 19756 9760 19772 9824
rect 19836 9760 19852 9824
rect 19916 9760 19924 9824
rect 19604 9759 19924 9760
rect 16849 9618 16915 9621
rect 18965 9618 19031 9621
rect 16849 9616 19031 9618
rect 16849 9560 16854 9616
rect 16910 9560 18970 9616
rect 19026 9560 19031 9616
rect 16849 9558 19031 9560
rect 16849 9555 16915 9558
rect 18965 9555 19031 9558
rect 19241 9618 19307 9621
rect 23800 9618 24600 9648
rect 19241 9616 24600 9618
rect 19241 9560 19246 9616
rect 19302 9560 24600 9616
rect 19241 9558 24600 9560
rect 19241 9555 19307 9558
rect 23800 9528 24600 9558
rect 8408 9280 8728 9281
rect 0 9210 800 9240
rect 8408 9216 8416 9280
rect 8480 9216 8496 9280
rect 8560 9216 8576 9280
rect 8640 9216 8656 9280
rect 8720 9216 8728 9280
rect 8408 9215 8728 9216
rect 15872 9280 16192 9281
rect 15872 9216 15880 9280
rect 15944 9216 15960 9280
rect 16024 9216 16040 9280
rect 16104 9216 16120 9280
rect 16184 9216 16192 9280
rect 15872 9215 16192 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 20345 8938 20411 8941
rect 23800 8938 24600 8968
rect 20345 8936 24600 8938
rect 20345 8880 20350 8936
rect 20406 8880 24600 8936
rect 20345 8878 24600 8880
rect 20345 8875 20411 8878
rect 23800 8848 24600 8878
rect 4676 8736 4996 8737
rect 4676 8672 4684 8736
rect 4748 8672 4764 8736
rect 4828 8672 4844 8736
rect 4908 8672 4924 8736
rect 4988 8672 4996 8736
rect 4676 8671 4996 8672
rect 12140 8736 12460 8737
rect 12140 8672 12148 8736
rect 12212 8672 12228 8736
rect 12292 8672 12308 8736
rect 12372 8672 12388 8736
rect 12452 8672 12460 8736
rect 12140 8671 12460 8672
rect 19604 8736 19924 8737
rect 19604 8672 19612 8736
rect 19676 8672 19692 8736
rect 19756 8672 19772 8736
rect 19836 8672 19852 8736
rect 19916 8672 19924 8736
rect 19604 8671 19924 8672
rect 21173 8258 21239 8261
rect 23800 8258 24600 8288
rect 21173 8256 24600 8258
rect 21173 8200 21178 8256
rect 21234 8200 24600 8256
rect 21173 8198 24600 8200
rect 21173 8195 21239 8198
rect 8408 8192 8728 8193
rect 8408 8128 8416 8192
rect 8480 8128 8496 8192
rect 8560 8128 8576 8192
rect 8640 8128 8656 8192
rect 8720 8128 8728 8192
rect 8408 8127 8728 8128
rect 15872 8192 16192 8193
rect 15872 8128 15880 8192
rect 15944 8128 15960 8192
rect 16024 8128 16040 8192
rect 16104 8128 16120 8192
rect 16184 8128 16192 8192
rect 23800 8168 24600 8198
rect 15872 8127 16192 8128
rect 15285 7986 15351 7989
rect 17309 7986 17375 7989
rect 15285 7984 17375 7986
rect 15285 7928 15290 7984
rect 15346 7928 17314 7984
rect 17370 7928 17375 7984
rect 15285 7926 17375 7928
rect 15285 7923 15351 7926
rect 17309 7923 17375 7926
rect 14549 7850 14615 7853
rect 16481 7850 16547 7853
rect 18137 7850 18203 7853
rect 14549 7848 18203 7850
rect 14549 7792 14554 7848
rect 14610 7792 16486 7848
rect 16542 7792 18142 7848
rect 18198 7792 18203 7848
rect 14549 7790 18203 7792
rect 14549 7787 14615 7790
rect 16481 7787 16547 7790
rect 18137 7787 18203 7790
rect 19701 7850 19767 7853
rect 20805 7850 20871 7853
rect 19701 7848 20871 7850
rect 19701 7792 19706 7848
rect 19762 7792 20810 7848
rect 20866 7792 20871 7848
rect 19701 7790 20871 7792
rect 19701 7787 19767 7790
rect 20805 7787 20871 7790
rect 4676 7648 4996 7649
rect 4676 7584 4684 7648
rect 4748 7584 4764 7648
rect 4828 7584 4844 7648
rect 4908 7584 4924 7648
rect 4988 7584 4996 7648
rect 4676 7583 4996 7584
rect 12140 7648 12460 7649
rect 12140 7584 12148 7648
rect 12212 7584 12228 7648
rect 12292 7584 12308 7648
rect 12372 7584 12388 7648
rect 12452 7584 12460 7648
rect 12140 7583 12460 7584
rect 19604 7648 19924 7649
rect 19604 7584 19612 7648
rect 19676 7584 19692 7648
rect 19756 7584 19772 7648
rect 19836 7584 19852 7648
rect 19916 7584 19924 7648
rect 19604 7583 19924 7584
rect 23289 7578 23355 7581
rect 23800 7578 24600 7608
rect 23289 7576 24600 7578
rect 23289 7520 23294 7576
rect 23350 7520 24600 7576
rect 23289 7518 24600 7520
rect 23289 7515 23355 7518
rect 23800 7488 24600 7518
rect 15837 7442 15903 7445
rect 19241 7442 19307 7445
rect 20161 7442 20227 7445
rect 15837 7440 20227 7442
rect 15837 7384 15842 7440
rect 15898 7384 19246 7440
rect 19302 7384 20166 7440
rect 20222 7384 20227 7440
rect 15837 7382 20227 7384
rect 15837 7379 15903 7382
rect 19241 7379 19307 7382
rect 20161 7379 20227 7382
rect 11881 7306 11947 7309
rect 17401 7306 17467 7309
rect 11881 7304 17467 7306
rect 11881 7248 11886 7304
rect 11942 7248 17406 7304
rect 17462 7248 17467 7304
rect 11881 7246 17467 7248
rect 11881 7243 11947 7246
rect 17401 7243 17467 7246
rect 20437 7306 20503 7309
rect 22093 7306 22159 7309
rect 20437 7304 22159 7306
rect 20437 7248 20442 7304
rect 20498 7248 22098 7304
rect 22154 7248 22159 7304
rect 20437 7246 22159 7248
rect 20437 7243 20503 7246
rect 22093 7243 22159 7246
rect 8408 7104 8728 7105
rect 8408 7040 8416 7104
rect 8480 7040 8496 7104
rect 8560 7040 8576 7104
rect 8640 7040 8656 7104
rect 8720 7040 8728 7104
rect 8408 7039 8728 7040
rect 15872 7104 16192 7105
rect 15872 7040 15880 7104
rect 15944 7040 15960 7104
rect 16024 7040 16040 7104
rect 16104 7040 16120 7104
rect 16184 7040 16192 7104
rect 15872 7039 16192 7040
rect 19333 7034 19399 7037
rect 23289 7034 23355 7037
rect 19333 7032 23355 7034
rect 19333 6976 19338 7032
rect 19394 6976 23294 7032
rect 23350 6976 23355 7032
rect 19333 6974 23355 6976
rect 19333 6971 19399 6974
rect 23289 6971 23355 6974
rect 20069 6898 20135 6901
rect 23800 6898 24600 6928
rect 20069 6896 24600 6898
rect 20069 6840 20074 6896
rect 20130 6840 24600 6896
rect 20069 6838 24600 6840
rect 20069 6835 20135 6838
rect 23800 6808 24600 6838
rect 4676 6560 4996 6561
rect 4676 6496 4684 6560
rect 4748 6496 4764 6560
rect 4828 6496 4844 6560
rect 4908 6496 4924 6560
rect 4988 6496 4996 6560
rect 4676 6495 4996 6496
rect 12140 6560 12460 6561
rect 12140 6496 12148 6560
rect 12212 6496 12228 6560
rect 12292 6496 12308 6560
rect 12372 6496 12388 6560
rect 12452 6496 12460 6560
rect 12140 6495 12460 6496
rect 19604 6560 19924 6561
rect 19604 6496 19612 6560
rect 19676 6496 19692 6560
rect 19756 6496 19772 6560
rect 19836 6496 19852 6560
rect 19916 6496 19924 6560
rect 19604 6495 19924 6496
rect 19977 6354 20043 6357
rect 23800 6354 24600 6384
rect 19977 6352 24600 6354
rect 19977 6296 19982 6352
rect 20038 6296 24600 6352
rect 19977 6294 24600 6296
rect 19977 6291 20043 6294
rect 23800 6264 24600 6294
rect 8408 6016 8728 6017
rect 8408 5952 8416 6016
rect 8480 5952 8496 6016
rect 8560 5952 8576 6016
rect 8640 5952 8656 6016
rect 8720 5952 8728 6016
rect 8408 5951 8728 5952
rect 15872 6016 16192 6017
rect 15872 5952 15880 6016
rect 15944 5952 15960 6016
rect 16024 5952 16040 6016
rect 16104 5952 16120 6016
rect 16184 5952 16192 6016
rect 15872 5951 16192 5952
rect 21357 5674 21423 5677
rect 23800 5674 24600 5704
rect 21357 5672 24600 5674
rect 21357 5616 21362 5672
rect 21418 5616 24600 5672
rect 21357 5614 24600 5616
rect 21357 5611 21423 5614
rect 23800 5584 24600 5614
rect 4676 5472 4996 5473
rect 4676 5408 4684 5472
rect 4748 5408 4764 5472
rect 4828 5408 4844 5472
rect 4908 5408 4924 5472
rect 4988 5408 4996 5472
rect 4676 5407 4996 5408
rect 12140 5472 12460 5473
rect 12140 5408 12148 5472
rect 12212 5408 12228 5472
rect 12292 5408 12308 5472
rect 12372 5408 12388 5472
rect 12452 5408 12460 5472
rect 12140 5407 12460 5408
rect 19604 5472 19924 5473
rect 19604 5408 19612 5472
rect 19676 5408 19692 5472
rect 19756 5408 19772 5472
rect 19836 5408 19852 5472
rect 19916 5408 19924 5472
rect 19604 5407 19924 5408
rect 20161 4994 20227 4997
rect 23800 4994 24600 5024
rect 20161 4992 24600 4994
rect 20161 4936 20166 4992
rect 20222 4936 24600 4992
rect 20161 4934 24600 4936
rect 20161 4931 20227 4934
rect 8408 4928 8728 4929
rect 8408 4864 8416 4928
rect 8480 4864 8496 4928
rect 8560 4864 8576 4928
rect 8640 4864 8656 4928
rect 8720 4864 8728 4928
rect 8408 4863 8728 4864
rect 15872 4928 16192 4929
rect 15872 4864 15880 4928
rect 15944 4864 15960 4928
rect 16024 4864 16040 4928
rect 16104 4864 16120 4928
rect 16184 4864 16192 4928
rect 23800 4904 24600 4934
rect 15872 4863 16192 4864
rect 4676 4384 4996 4385
rect 4676 4320 4684 4384
rect 4748 4320 4764 4384
rect 4828 4320 4844 4384
rect 4908 4320 4924 4384
rect 4988 4320 4996 4384
rect 4676 4319 4996 4320
rect 12140 4384 12460 4385
rect 12140 4320 12148 4384
rect 12212 4320 12228 4384
rect 12292 4320 12308 4384
rect 12372 4320 12388 4384
rect 12452 4320 12460 4384
rect 12140 4319 12460 4320
rect 19604 4384 19924 4385
rect 19604 4320 19612 4384
rect 19676 4320 19692 4384
rect 19756 4320 19772 4384
rect 19836 4320 19852 4384
rect 19916 4320 19924 4384
rect 19604 4319 19924 4320
rect 20529 4314 20595 4317
rect 23800 4314 24600 4344
rect 20529 4312 24600 4314
rect 20529 4256 20534 4312
rect 20590 4256 24600 4312
rect 20529 4254 24600 4256
rect 20529 4251 20595 4254
rect 23800 4224 24600 4254
rect 8408 3840 8728 3841
rect 8408 3776 8416 3840
rect 8480 3776 8496 3840
rect 8560 3776 8576 3840
rect 8640 3776 8656 3840
rect 8720 3776 8728 3840
rect 8408 3775 8728 3776
rect 15872 3840 16192 3841
rect 15872 3776 15880 3840
rect 15944 3776 15960 3840
rect 16024 3776 16040 3840
rect 16104 3776 16120 3840
rect 16184 3776 16192 3840
rect 15872 3775 16192 3776
rect 19885 3634 19951 3637
rect 23800 3634 24600 3664
rect 19885 3632 24600 3634
rect 19885 3576 19890 3632
rect 19946 3576 24600 3632
rect 19885 3574 24600 3576
rect 19885 3571 19951 3574
rect 23800 3544 24600 3574
rect 4676 3296 4996 3297
rect 4676 3232 4684 3296
rect 4748 3232 4764 3296
rect 4828 3232 4844 3296
rect 4908 3232 4924 3296
rect 4988 3232 4996 3296
rect 4676 3231 4996 3232
rect 12140 3296 12460 3297
rect 12140 3232 12148 3296
rect 12212 3232 12228 3296
rect 12292 3232 12308 3296
rect 12372 3232 12388 3296
rect 12452 3232 12460 3296
rect 12140 3231 12460 3232
rect 19604 3296 19924 3297
rect 19604 3232 19612 3296
rect 19676 3232 19692 3296
rect 19756 3232 19772 3296
rect 19836 3232 19852 3296
rect 19916 3232 19924 3296
rect 19604 3231 19924 3232
rect 0 3090 800 3120
rect 1393 3090 1459 3093
rect 0 3088 1459 3090
rect 0 3032 1398 3088
rect 1454 3032 1459 3088
rect 0 3030 1459 3032
rect 0 3000 800 3030
rect 1393 3027 1459 3030
rect 20253 3090 20319 3093
rect 21357 3090 21423 3093
rect 20253 3088 21423 3090
rect 20253 3032 20258 3088
rect 20314 3032 21362 3088
rect 21418 3032 21423 3088
rect 20253 3030 21423 3032
rect 20253 3027 20319 3030
rect 21357 3027 21423 3030
rect 20529 2954 20595 2957
rect 23800 2954 24600 2984
rect 20529 2952 24600 2954
rect 20529 2896 20534 2952
rect 20590 2896 24600 2952
rect 20529 2894 24600 2896
rect 20529 2891 20595 2894
rect 23800 2864 24600 2894
rect 8408 2752 8728 2753
rect 8408 2688 8416 2752
rect 8480 2688 8496 2752
rect 8560 2688 8576 2752
rect 8640 2688 8656 2752
rect 8720 2688 8728 2752
rect 8408 2687 8728 2688
rect 15872 2752 16192 2753
rect 15872 2688 15880 2752
rect 15944 2688 15960 2752
rect 16024 2688 16040 2752
rect 16104 2688 16120 2752
rect 16184 2688 16192 2752
rect 15872 2687 16192 2688
rect 21909 2274 21975 2277
rect 23800 2274 24600 2304
rect 21909 2272 24600 2274
rect 21909 2216 21914 2272
rect 21970 2216 24600 2272
rect 21909 2214 24600 2216
rect 21909 2211 21975 2214
rect 4676 2208 4996 2209
rect 4676 2144 4684 2208
rect 4748 2144 4764 2208
rect 4828 2144 4844 2208
rect 4908 2144 4924 2208
rect 4988 2144 4996 2208
rect 4676 2143 4996 2144
rect 12140 2208 12460 2209
rect 12140 2144 12148 2208
rect 12212 2144 12228 2208
rect 12292 2144 12308 2208
rect 12372 2144 12388 2208
rect 12452 2144 12460 2208
rect 12140 2143 12460 2144
rect 19604 2208 19924 2209
rect 19604 2144 19612 2208
rect 19676 2144 19692 2208
rect 19756 2144 19772 2208
rect 19836 2144 19852 2208
rect 19916 2144 19924 2208
rect 23800 2184 24600 2214
rect 19604 2143 19924 2144
rect 23013 1594 23079 1597
rect 23800 1594 24600 1624
rect 23013 1592 24600 1594
rect 23013 1536 23018 1592
rect 23074 1536 24600 1592
rect 23013 1534 24600 1536
rect 23013 1531 23079 1534
rect 23800 1504 24600 1534
rect 22001 914 22067 917
rect 23800 914 24600 944
rect 22001 912 24600 914
rect 22001 856 22006 912
rect 22062 856 24600 912
rect 22001 854 24600 856
rect 22001 851 22067 854
rect 23800 824 24600 854
rect 23565 370 23631 373
rect 23800 370 24600 400
rect 23565 368 24600 370
rect 23565 312 23570 368
rect 23626 312 24600 368
rect 23565 310 24600 312
rect 23565 307 23631 310
rect 23800 280 24600 310
<< via3 >>
rect 8416 22332 8480 22336
rect 8416 22276 8420 22332
rect 8420 22276 8476 22332
rect 8476 22276 8480 22332
rect 8416 22272 8480 22276
rect 8496 22332 8560 22336
rect 8496 22276 8500 22332
rect 8500 22276 8556 22332
rect 8556 22276 8560 22332
rect 8496 22272 8560 22276
rect 8576 22332 8640 22336
rect 8576 22276 8580 22332
rect 8580 22276 8636 22332
rect 8636 22276 8640 22332
rect 8576 22272 8640 22276
rect 8656 22332 8720 22336
rect 8656 22276 8660 22332
rect 8660 22276 8716 22332
rect 8716 22276 8720 22332
rect 8656 22272 8720 22276
rect 15880 22332 15944 22336
rect 15880 22276 15884 22332
rect 15884 22276 15940 22332
rect 15940 22276 15944 22332
rect 15880 22272 15944 22276
rect 15960 22332 16024 22336
rect 15960 22276 15964 22332
rect 15964 22276 16020 22332
rect 16020 22276 16024 22332
rect 15960 22272 16024 22276
rect 16040 22332 16104 22336
rect 16040 22276 16044 22332
rect 16044 22276 16100 22332
rect 16100 22276 16104 22332
rect 16040 22272 16104 22276
rect 16120 22332 16184 22336
rect 16120 22276 16124 22332
rect 16124 22276 16180 22332
rect 16180 22276 16184 22332
rect 16120 22272 16184 22276
rect 4684 21788 4748 21792
rect 4684 21732 4688 21788
rect 4688 21732 4744 21788
rect 4744 21732 4748 21788
rect 4684 21728 4748 21732
rect 4764 21788 4828 21792
rect 4764 21732 4768 21788
rect 4768 21732 4824 21788
rect 4824 21732 4828 21788
rect 4764 21728 4828 21732
rect 4844 21788 4908 21792
rect 4844 21732 4848 21788
rect 4848 21732 4904 21788
rect 4904 21732 4908 21788
rect 4844 21728 4908 21732
rect 4924 21788 4988 21792
rect 4924 21732 4928 21788
rect 4928 21732 4984 21788
rect 4984 21732 4988 21788
rect 4924 21728 4988 21732
rect 12148 21788 12212 21792
rect 12148 21732 12152 21788
rect 12152 21732 12208 21788
rect 12208 21732 12212 21788
rect 12148 21728 12212 21732
rect 12228 21788 12292 21792
rect 12228 21732 12232 21788
rect 12232 21732 12288 21788
rect 12288 21732 12292 21788
rect 12228 21728 12292 21732
rect 12308 21788 12372 21792
rect 12308 21732 12312 21788
rect 12312 21732 12368 21788
rect 12368 21732 12372 21788
rect 12308 21728 12372 21732
rect 12388 21788 12452 21792
rect 12388 21732 12392 21788
rect 12392 21732 12448 21788
rect 12448 21732 12452 21788
rect 12388 21728 12452 21732
rect 19612 21788 19676 21792
rect 19612 21732 19616 21788
rect 19616 21732 19672 21788
rect 19672 21732 19676 21788
rect 19612 21728 19676 21732
rect 19692 21788 19756 21792
rect 19692 21732 19696 21788
rect 19696 21732 19752 21788
rect 19752 21732 19756 21788
rect 19692 21728 19756 21732
rect 19772 21788 19836 21792
rect 19772 21732 19776 21788
rect 19776 21732 19832 21788
rect 19832 21732 19836 21788
rect 19772 21728 19836 21732
rect 19852 21788 19916 21792
rect 19852 21732 19856 21788
rect 19856 21732 19912 21788
rect 19912 21732 19916 21788
rect 19852 21728 19916 21732
rect 8416 21244 8480 21248
rect 8416 21188 8420 21244
rect 8420 21188 8476 21244
rect 8476 21188 8480 21244
rect 8416 21184 8480 21188
rect 8496 21244 8560 21248
rect 8496 21188 8500 21244
rect 8500 21188 8556 21244
rect 8556 21188 8560 21244
rect 8496 21184 8560 21188
rect 8576 21244 8640 21248
rect 8576 21188 8580 21244
rect 8580 21188 8636 21244
rect 8636 21188 8640 21244
rect 8576 21184 8640 21188
rect 8656 21244 8720 21248
rect 8656 21188 8660 21244
rect 8660 21188 8716 21244
rect 8716 21188 8720 21244
rect 8656 21184 8720 21188
rect 15880 21244 15944 21248
rect 15880 21188 15884 21244
rect 15884 21188 15940 21244
rect 15940 21188 15944 21244
rect 15880 21184 15944 21188
rect 15960 21244 16024 21248
rect 15960 21188 15964 21244
rect 15964 21188 16020 21244
rect 16020 21188 16024 21244
rect 15960 21184 16024 21188
rect 16040 21244 16104 21248
rect 16040 21188 16044 21244
rect 16044 21188 16100 21244
rect 16100 21188 16104 21244
rect 16040 21184 16104 21188
rect 16120 21244 16184 21248
rect 16120 21188 16124 21244
rect 16124 21188 16180 21244
rect 16180 21188 16184 21244
rect 16120 21184 16184 21188
rect 4684 20700 4748 20704
rect 4684 20644 4688 20700
rect 4688 20644 4744 20700
rect 4744 20644 4748 20700
rect 4684 20640 4748 20644
rect 4764 20700 4828 20704
rect 4764 20644 4768 20700
rect 4768 20644 4824 20700
rect 4824 20644 4828 20700
rect 4764 20640 4828 20644
rect 4844 20700 4908 20704
rect 4844 20644 4848 20700
rect 4848 20644 4904 20700
rect 4904 20644 4908 20700
rect 4844 20640 4908 20644
rect 4924 20700 4988 20704
rect 4924 20644 4928 20700
rect 4928 20644 4984 20700
rect 4984 20644 4988 20700
rect 4924 20640 4988 20644
rect 12148 20700 12212 20704
rect 12148 20644 12152 20700
rect 12152 20644 12208 20700
rect 12208 20644 12212 20700
rect 12148 20640 12212 20644
rect 12228 20700 12292 20704
rect 12228 20644 12232 20700
rect 12232 20644 12288 20700
rect 12288 20644 12292 20700
rect 12228 20640 12292 20644
rect 12308 20700 12372 20704
rect 12308 20644 12312 20700
rect 12312 20644 12368 20700
rect 12368 20644 12372 20700
rect 12308 20640 12372 20644
rect 12388 20700 12452 20704
rect 12388 20644 12392 20700
rect 12392 20644 12448 20700
rect 12448 20644 12452 20700
rect 12388 20640 12452 20644
rect 19612 20700 19676 20704
rect 19612 20644 19616 20700
rect 19616 20644 19672 20700
rect 19672 20644 19676 20700
rect 19612 20640 19676 20644
rect 19692 20700 19756 20704
rect 19692 20644 19696 20700
rect 19696 20644 19752 20700
rect 19752 20644 19756 20700
rect 19692 20640 19756 20644
rect 19772 20700 19836 20704
rect 19772 20644 19776 20700
rect 19776 20644 19832 20700
rect 19832 20644 19836 20700
rect 19772 20640 19836 20644
rect 19852 20700 19916 20704
rect 19852 20644 19856 20700
rect 19856 20644 19912 20700
rect 19912 20644 19916 20700
rect 19852 20640 19916 20644
rect 8416 20156 8480 20160
rect 8416 20100 8420 20156
rect 8420 20100 8476 20156
rect 8476 20100 8480 20156
rect 8416 20096 8480 20100
rect 8496 20156 8560 20160
rect 8496 20100 8500 20156
rect 8500 20100 8556 20156
rect 8556 20100 8560 20156
rect 8496 20096 8560 20100
rect 8576 20156 8640 20160
rect 8576 20100 8580 20156
rect 8580 20100 8636 20156
rect 8636 20100 8640 20156
rect 8576 20096 8640 20100
rect 8656 20156 8720 20160
rect 8656 20100 8660 20156
rect 8660 20100 8716 20156
rect 8716 20100 8720 20156
rect 8656 20096 8720 20100
rect 15880 20156 15944 20160
rect 15880 20100 15884 20156
rect 15884 20100 15940 20156
rect 15940 20100 15944 20156
rect 15880 20096 15944 20100
rect 15960 20156 16024 20160
rect 15960 20100 15964 20156
rect 15964 20100 16020 20156
rect 16020 20100 16024 20156
rect 15960 20096 16024 20100
rect 16040 20156 16104 20160
rect 16040 20100 16044 20156
rect 16044 20100 16100 20156
rect 16100 20100 16104 20156
rect 16040 20096 16104 20100
rect 16120 20156 16184 20160
rect 16120 20100 16124 20156
rect 16124 20100 16180 20156
rect 16180 20100 16184 20156
rect 16120 20096 16184 20100
rect 4684 19612 4748 19616
rect 4684 19556 4688 19612
rect 4688 19556 4744 19612
rect 4744 19556 4748 19612
rect 4684 19552 4748 19556
rect 4764 19612 4828 19616
rect 4764 19556 4768 19612
rect 4768 19556 4824 19612
rect 4824 19556 4828 19612
rect 4764 19552 4828 19556
rect 4844 19612 4908 19616
rect 4844 19556 4848 19612
rect 4848 19556 4904 19612
rect 4904 19556 4908 19612
rect 4844 19552 4908 19556
rect 4924 19612 4988 19616
rect 4924 19556 4928 19612
rect 4928 19556 4984 19612
rect 4984 19556 4988 19612
rect 4924 19552 4988 19556
rect 12148 19612 12212 19616
rect 12148 19556 12152 19612
rect 12152 19556 12208 19612
rect 12208 19556 12212 19612
rect 12148 19552 12212 19556
rect 12228 19612 12292 19616
rect 12228 19556 12232 19612
rect 12232 19556 12288 19612
rect 12288 19556 12292 19612
rect 12228 19552 12292 19556
rect 12308 19612 12372 19616
rect 12308 19556 12312 19612
rect 12312 19556 12368 19612
rect 12368 19556 12372 19612
rect 12308 19552 12372 19556
rect 12388 19612 12452 19616
rect 12388 19556 12392 19612
rect 12392 19556 12448 19612
rect 12448 19556 12452 19612
rect 12388 19552 12452 19556
rect 19612 19612 19676 19616
rect 19612 19556 19616 19612
rect 19616 19556 19672 19612
rect 19672 19556 19676 19612
rect 19612 19552 19676 19556
rect 19692 19612 19756 19616
rect 19692 19556 19696 19612
rect 19696 19556 19752 19612
rect 19752 19556 19756 19612
rect 19692 19552 19756 19556
rect 19772 19612 19836 19616
rect 19772 19556 19776 19612
rect 19776 19556 19832 19612
rect 19832 19556 19836 19612
rect 19772 19552 19836 19556
rect 19852 19612 19916 19616
rect 19852 19556 19856 19612
rect 19856 19556 19912 19612
rect 19912 19556 19916 19612
rect 19852 19552 19916 19556
rect 8416 19068 8480 19072
rect 8416 19012 8420 19068
rect 8420 19012 8476 19068
rect 8476 19012 8480 19068
rect 8416 19008 8480 19012
rect 8496 19068 8560 19072
rect 8496 19012 8500 19068
rect 8500 19012 8556 19068
rect 8556 19012 8560 19068
rect 8496 19008 8560 19012
rect 8576 19068 8640 19072
rect 8576 19012 8580 19068
rect 8580 19012 8636 19068
rect 8636 19012 8640 19068
rect 8576 19008 8640 19012
rect 8656 19068 8720 19072
rect 8656 19012 8660 19068
rect 8660 19012 8716 19068
rect 8716 19012 8720 19068
rect 8656 19008 8720 19012
rect 15880 19068 15944 19072
rect 15880 19012 15884 19068
rect 15884 19012 15940 19068
rect 15940 19012 15944 19068
rect 15880 19008 15944 19012
rect 15960 19068 16024 19072
rect 15960 19012 15964 19068
rect 15964 19012 16020 19068
rect 16020 19012 16024 19068
rect 15960 19008 16024 19012
rect 16040 19068 16104 19072
rect 16040 19012 16044 19068
rect 16044 19012 16100 19068
rect 16100 19012 16104 19068
rect 16040 19008 16104 19012
rect 16120 19068 16184 19072
rect 16120 19012 16124 19068
rect 16124 19012 16180 19068
rect 16180 19012 16184 19068
rect 16120 19008 16184 19012
rect 4684 18524 4748 18528
rect 4684 18468 4688 18524
rect 4688 18468 4744 18524
rect 4744 18468 4748 18524
rect 4684 18464 4748 18468
rect 4764 18524 4828 18528
rect 4764 18468 4768 18524
rect 4768 18468 4824 18524
rect 4824 18468 4828 18524
rect 4764 18464 4828 18468
rect 4844 18524 4908 18528
rect 4844 18468 4848 18524
rect 4848 18468 4904 18524
rect 4904 18468 4908 18524
rect 4844 18464 4908 18468
rect 4924 18524 4988 18528
rect 4924 18468 4928 18524
rect 4928 18468 4984 18524
rect 4984 18468 4988 18524
rect 4924 18464 4988 18468
rect 12148 18524 12212 18528
rect 12148 18468 12152 18524
rect 12152 18468 12208 18524
rect 12208 18468 12212 18524
rect 12148 18464 12212 18468
rect 12228 18524 12292 18528
rect 12228 18468 12232 18524
rect 12232 18468 12288 18524
rect 12288 18468 12292 18524
rect 12228 18464 12292 18468
rect 12308 18524 12372 18528
rect 12308 18468 12312 18524
rect 12312 18468 12368 18524
rect 12368 18468 12372 18524
rect 12308 18464 12372 18468
rect 12388 18524 12452 18528
rect 12388 18468 12392 18524
rect 12392 18468 12448 18524
rect 12448 18468 12452 18524
rect 12388 18464 12452 18468
rect 19612 18524 19676 18528
rect 19612 18468 19616 18524
rect 19616 18468 19672 18524
rect 19672 18468 19676 18524
rect 19612 18464 19676 18468
rect 19692 18524 19756 18528
rect 19692 18468 19696 18524
rect 19696 18468 19752 18524
rect 19752 18468 19756 18524
rect 19692 18464 19756 18468
rect 19772 18524 19836 18528
rect 19772 18468 19776 18524
rect 19776 18468 19832 18524
rect 19832 18468 19836 18524
rect 19772 18464 19836 18468
rect 19852 18524 19916 18528
rect 19852 18468 19856 18524
rect 19856 18468 19912 18524
rect 19912 18468 19916 18524
rect 19852 18464 19916 18468
rect 8416 17980 8480 17984
rect 8416 17924 8420 17980
rect 8420 17924 8476 17980
rect 8476 17924 8480 17980
rect 8416 17920 8480 17924
rect 8496 17980 8560 17984
rect 8496 17924 8500 17980
rect 8500 17924 8556 17980
rect 8556 17924 8560 17980
rect 8496 17920 8560 17924
rect 8576 17980 8640 17984
rect 8576 17924 8580 17980
rect 8580 17924 8636 17980
rect 8636 17924 8640 17980
rect 8576 17920 8640 17924
rect 8656 17980 8720 17984
rect 8656 17924 8660 17980
rect 8660 17924 8716 17980
rect 8716 17924 8720 17980
rect 8656 17920 8720 17924
rect 15880 17980 15944 17984
rect 15880 17924 15884 17980
rect 15884 17924 15940 17980
rect 15940 17924 15944 17980
rect 15880 17920 15944 17924
rect 15960 17980 16024 17984
rect 15960 17924 15964 17980
rect 15964 17924 16020 17980
rect 16020 17924 16024 17980
rect 15960 17920 16024 17924
rect 16040 17980 16104 17984
rect 16040 17924 16044 17980
rect 16044 17924 16100 17980
rect 16100 17924 16104 17980
rect 16040 17920 16104 17924
rect 16120 17980 16184 17984
rect 16120 17924 16124 17980
rect 16124 17924 16180 17980
rect 16180 17924 16184 17980
rect 16120 17920 16184 17924
rect 4684 17436 4748 17440
rect 4684 17380 4688 17436
rect 4688 17380 4744 17436
rect 4744 17380 4748 17436
rect 4684 17376 4748 17380
rect 4764 17436 4828 17440
rect 4764 17380 4768 17436
rect 4768 17380 4824 17436
rect 4824 17380 4828 17436
rect 4764 17376 4828 17380
rect 4844 17436 4908 17440
rect 4844 17380 4848 17436
rect 4848 17380 4904 17436
rect 4904 17380 4908 17436
rect 4844 17376 4908 17380
rect 4924 17436 4988 17440
rect 4924 17380 4928 17436
rect 4928 17380 4984 17436
rect 4984 17380 4988 17436
rect 4924 17376 4988 17380
rect 12148 17436 12212 17440
rect 12148 17380 12152 17436
rect 12152 17380 12208 17436
rect 12208 17380 12212 17436
rect 12148 17376 12212 17380
rect 12228 17436 12292 17440
rect 12228 17380 12232 17436
rect 12232 17380 12288 17436
rect 12288 17380 12292 17436
rect 12228 17376 12292 17380
rect 12308 17436 12372 17440
rect 12308 17380 12312 17436
rect 12312 17380 12368 17436
rect 12368 17380 12372 17436
rect 12308 17376 12372 17380
rect 12388 17436 12452 17440
rect 12388 17380 12392 17436
rect 12392 17380 12448 17436
rect 12448 17380 12452 17436
rect 12388 17376 12452 17380
rect 19612 17436 19676 17440
rect 19612 17380 19616 17436
rect 19616 17380 19672 17436
rect 19672 17380 19676 17436
rect 19612 17376 19676 17380
rect 19692 17436 19756 17440
rect 19692 17380 19696 17436
rect 19696 17380 19752 17436
rect 19752 17380 19756 17436
rect 19692 17376 19756 17380
rect 19772 17436 19836 17440
rect 19772 17380 19776 17436
rect 19776 17380 19832 17436
rect 19832 17380 19836 17436
rect 19772 17376 19836 17380
rect 19852 17436 19916 17440
rect 19852 17380 19856 17436
rect 19856 17380 19912 17436
rect 19912 17380 19916 17436
rect 19852 17376 19916 17380
rect 8416 16892 8480 16896
rect 8416 16836 8420 16892
rect 8420 16836 8476 16892
rect 8476 16836 8480 16892
rect 8416 16832 8480 16836
rect 8496 16892 8560 16896
rect 8496 16836 8500 16892
rect 8500 16836 8556 16892
rect 8556 16836 8560 16892
rect 8496 16832 8560 16836
rect 8576 16892 8640 16896
rect 8576 16836 8580 16892
rect 8580 16836 8636 16892
rect 8636 16836 8640 16892
rect 8576 16832 8640 16836
rect 8656 16892 8720 16896
rect 8656 16836 8660 16892
rect 8660 16836 8716 16892
rect 8716 16836 8720 16892
rect 8656 16832 8720 16836
rect 15880 16892 15944 16896
rect 15880 16836 15884 16892
rect 15884 16836 15940 16892
rect 15940 16836 15944 16892
rect 15880 16832 15944 16836
rect 15960 16892 16024 16896
rect 15960 16836 15964 16892
rect 15964 16836 16020 16892
rect 16020 16836 16024 16892
rect 15960 16832 16024 16836
rect 16040 16892 16104 16896
rect 16040 16836 16044 16892
rect 16044 16836 16100 16892
rect 16100 16836 16104 16892
rect 16040 16832 16104 16836
rect 16120 16892 16184 16896
rect 16120 16836 16124 16892
rect 16124 16836 16180 16892
rect 16180 16836 16184 16892
rect 16120 16832 16184 16836
rect 4684 16348 4748 16352
rect 4684 16292 4688 16348
rect 4688 16292 4744 16348
rect 4744 16292 4748 16348
rect 4684 16288 4748 16292
rect 4764 16348 4828 16352
rect 4764 16292 4768 16348
rect 4768 16292 4824 16348
rect 4824 16292 4828 16348
rect 4764 16288 4828 16292
rect 4844 16348 4908 16352
rect 4844 16292 4848 16348
rect 4848 16292 4904 16348
rect 4904 16292 4908 16348
rect 4844 16288 4908 16292
rect 4924 16348 4988 16352
rect 4924 16292 4928 16348
rect 4928 16292 4984 16348
rect 4984 16292 4988 16348
rect 4924 16288 4988 16292
rect 12148 16348 12212 16352
rect 12148 16292 12152 16348
rect 12152 16292 12208 16348
rect 12208 16292 12212 16348
rect 12148 16288 12212 16292
rect 12228 16348 12292 16352
rect 12228 16292 12232 16348
rect 12232 16292 12288 16348
rect 12288 16292 12292 16348
rect 12228 16288 12292 16292
rect 12308 16348 12372 16352
rect 12308 16292 12312 16348
rect 12312 16292 12368 16348
rect 12368 16292 12372 16348
rect 12308 16288 12372 16292
rect 12388 16348 12452 16352
rect 12388 16292 12392 16348
rect 12392 16292 12448 16348
rect 12448 16292 12452 16348
rect 12388 16288 12452 16292
rect 19612 16348 19676 16352
rect 19612 16292 19616 16348
rect 19616 16292 19672 16348
rect 19672 16292 19676 16348
rect 19612 16288 19676 16292
rect 19692 16348 19756 16352
rect 19692 16292 19696 16348
rect 19696 16292 19752 16348
rect 19752 16292 19756 16348
rect 19692 16288 19756 16292
rect 19772 16348 19836 16352
rect 19772 16292 19776 16348
rect 19776 16292 19832 16348
rect 19832 16292 19836 16348
rect 19772 16288 19836 16292
rect 19852 16348 19916 16352
rect 19852 16292 19856 16348
rect 19856 16292 19912 16348
rect 19912 16292 19916 16348
rect 19852 16288 19916 16292
rect 8416 15804 8480 15808
rect 8416 15748 8420 15804
rect 8420 15748 8476 15804
rect 8476 15748 8480 15804
rect 8416 15744 8480 15748
rect 8496 15804 8560 15808
rect 8496 15748 8500 15804
rect 8500 15748 8556 15804
rect 8556 15748 8560 15804
rect 8496 15744 8560 15748
rect 8576 15804 8640 15808
rect 8576 15748 8580 15804
rect 8580 15748 8636 15804
rect 8636 15748 8640 15804
rect 8576 15744 8640 15748
rect 8656 15804 8720 15808
rect 8656 15748 8660 15804
rect 8660 15748 8716 15804
rect 8716 15748 8720 15804
rect 8656 15744 8720 15748
rect 15880 15804 15944 15808
rect 15880 15748 15884 15804
rect 15884 15748 15940 15804
rect 15940 15748 15944 15804
rect 15880 15744 15944 15748
rect 15960 15804 16024 15808
rect 15960 15748 15964 15804
rect 15964 15748 16020 15804
rect 16020 15748 16024 15804
rect 15960 15744 16024 15748
rect 16040 15804 16104 15808
rect 16040 15748 16044 15804
rect 16044 15748 16100 15804
rect 16100 15748 16104 15804
rect 16040 15744 16104 15748
rect 16120 15804 16184 15808
rect 16120 15748 16124 15804
rect 16124 15748 16180 15804
rect 16180 15748 16184 15804
rect 16120 15744 16184 15748
rect 20116 15676 20180 15740
rect 4684 15260 4748 15264
rect 4684 15204 4688 15260
rect 4688 15204 4744 15260
rect 4744 15204 4748 15260
rect 4684 15200 4748 15204
rect 4764 15260 4828 15264
rect 4764 15204 4768 15260
rect 4768 15204 4824 15260
rect 4824 15204 4828 15260
rect 4764 15200 4828 15204
rect 4844 15260 4908 15264
rect 4844 15204 4848 15260
rect 4848 15204 4904 15260
rect 4904 15204 4908 15260
rect 4844 15200 4908 15204
rect 4924 15260 4988 15264
rect 4924 15204 4928 15260
rect 4928 15204 4984 15260
rect 4984 15204 4988 15260
rect 4924 15200 4988 15204
rect 12148 15260 12212 15264
rect 12148 15204 12152 15260
rect 12152 15204 12208 15260
rect 12208 15204 12212 15260
rect 12148 15200 12212 15204
rect 12228 15260 12292 15264
rect 12228 15204 12232 15260
rect 12232 15204 12288 15260
rect 12288 15204 12292 15260
rect 12228 15200 12292 15204
rect 12308 15260 12372 15264
rect 12308 15204 12312 15260
rect 12312 15204 12368 15260
rect 12368 15204 12372 15260
rect 12308 15200 12372 15204
rect 12388 15260 12452 15264
rect 12388 15204 12392 15260
rect 12392 15204 12448 15260
rect 12448 15204 12452 15260
rect 12388 15200 12452 15204
rect 19612 15260 19676 15264
rect 19612 15204 19616 15260
rect 19616 15204 19672 15260
rect 19672 15204 19676 15260
rect 19612 15200 19676 15204
rect 19692 15260 19756 15264
rect 19692 15204 19696 15260
rect 19696 15204 19752 15260
rect 19752 15204 19756 15260
rect 19692 15200 19756 15204
rect 19772 15260 19836 15264
rect 19772 15204 19776 15260
rect 19776 15204 19832 15260
rect 19832 15204 19836 15260
rect 19772 15200 19836 15204
rect 19852 15260 19916 15264
rect 19852 15204 19856 15260
rect 19856 15204 19912 15260
rect 19912 15204 19916 15260
rect 19852 15200 19916 15204
rect 8416 14716 8480 14720
rect 8416 14660 8420 14716
rect 8420 14660 8476 14716
rect 8476 14660 8480 14716
rect 8416 14656 8480 14660
rect 8496 14716 8560 14720
rect 8496 14660 8500 14716
rect 8500 14660 8556 14716
rect 8556 14660 8560 14716
rect 8496 14656 8560 14660
rect 8576 14716 8640 14720
rect 8576 14660 8580 14716
rect 8580 14660 8636 14716
rect 8636 14660 8640 14716
rect 8576 14656 8640 14660
rect 8656 14716 8720 14720
rect 8656 14660 8660 14716
rect 8660 14660 8716 14716
rect 8716 14660 8720 14716
rect 8656 14656 8720 14660
rect 15880 14716 15944 14720
rect 15880 14660 15884 14716
rect 15884 14660 15940 14716
rect 15940 14660 15944 14716
rect 15880 14656 15944 14660
rect 15960 14716 16024 14720
rect 15960 14660 15964 14716
rect 15964 14660 16020 14716
rect 16020 14660 16024 14716
rect 15960 14656 16024 14660
rect 16040 14716 16104 14720
rect 16040 14660 16044 14716
rect 16044 14660 16100 14716
rect 16100 14660 16104 14716
rect 16040 14656 16104 14660
rect 16120 14716 16184 14720
rect 16120 14660 16124 14716
rect 16124 14660 16180 14716
rect 16180 14660 16184 14716
rect 16120 14656 16184 14660
rect 4684 14172 4748 14176
rect 4684 14116 4688 14172
rect 4688 14116 4744 14172
rect 4744 14116 4748 14172
rect 4684 14112 4748 14116
rect 4764 14172 4828 14176
rect 4764 14116 4768 14172
rect 4768 14116 4824 14172
rect 4824 14116 4828 14172
rect 4764 14112 4828 14116
rect 4844 14172 4908 14176
rect 4844 14116 4848 14172
rect 4848 14116 4904 14172
rect 4904 14116 4908 14172
rect 4844 14112 4908 14116
rect 4924 14172 4988 14176
rect 4924 14116 4928 14172
rect 4928 14116 4984 14172
rect 4984 14116 4988 14172
rect 4924 14112 4988 14116
rect 12148 14172 12212 14176
rect 12148 14116 12152 14172
rect 12152 14116 12208 14172
rect 12208 14116 12212 14172
rect 12148 14112 12212 14116
rect 12228 14172 12292 14176
rect 12228 14116 12232 14172
rect 12232 14116 12288 14172
rect 12288 14116 12292 14172
rect 12228 14112 12292 14116
rect 12308 14172 12372 14176
rect 12308 14116 12312 14172
rect 12312 14116 12368 14172
rect 12368 14116 12372 14172
rect 12308 14112 12372 14116
rect 12388 14172 12452 14176
rect 12388 14116 12392 14172
rect 12392 14116 12448 14172
rect 12448 14116 12452 14172
rect 12388 14112 12452 14116
rect 19612 14172 19676 14176
rect 19612 14116 19616 14172
rect 19616 14116 19672 14172
rect 19672 14116 19676 14172
rect 19612 14112 19676 14116
rect 19692 14172 19756 14176
rect 19692 14116 19696 14172
rect 19696 14116 19752 14172
rect 19752 14116 19756 14172
rect 19692 14112 19756 14116
rect 19772 14172 19836 14176
rect 19772 14116 19776 14172
rect 19776 14116 19832 14172
rect 19832 14116 19836 14172
rect 19772 14112 19836 14116
rect 19852 14172 19916 14176
rect 19852 14116 19856 14172
rect 19856 14116 19912 14172
rect 19912 14116 19916 14172
rect 19852 14112 19916 14116
rect 8416 13628 8480 13632
rect 8416 13572 8420 13628
rect 8420 13572 8476 13628
rect 8476 13572 8480 13628
rect 8416 13568 8480 13572
rect 8496 13628 8560 13632
rect 8496 13572 8500 13628
rect 8500 13572 8556 13628
rect 8556 13572 8560 13628
rect 8496 13568 8560 13572
rect 8576 13628 8640 13632
rect 8576 13572 8580 13628
rect 8580 13572 8636 13628
rect 8636 13572 8640 13628
rect 8576 13568 8640 13572
rect 8656 13628 8720 13632
rect 8656 13572 8660 13628
rect 8660 13572 8716 13628
rect 8716 13572 8720 13628
rect 8656 13568 8720 13572
rect 15880 13628 15944 13632
rect 15880 13572 15884 13628
rect 15884 13572 15940 13628
rect 15940 13572 15944 13628
rect 15880 13568 15944 13572
rect 15960 13628 16024 13632
rect 15960 13572 15964 13628
rect 15964 13572 16020 13628
rect 16020 13572 16024 13628
rect 15960 13568 16024 13572
rect 16040 13628 16104 13632
rect 16040 13572 16044 13628
rect 16044 13572 16100 13628
rect 16100 13572 16104 13628
rect 16040 13568 16104 13572
rect 16120 13628 16184 13632
rect 16120 13572 16124 13628
rect 16124 13572 16180 13628
rect 16180 13572 16184 13628
rect 16120 13568 16184 13572
rect 20484 13288 20548 13292
rect 20484 13232 20498 13288
rect 20498 13232 20548 13288
rect 20484 13228 20548 13232
rect 4684 13084 4748 13088
rect 4684 13028 4688 13084
rect 4688 13028 4744 13084
rect 4744 13028 4748 13084
rect 4684 13024 4748 13028
rect 4764 13084 4828 13088
rect 4764 13028 4768 13084
rect 4768 13028 4824 13084
rect 4824 13028 4828 13084
rect 4764 13024 4828 13028
rect 4844 13084 4908 13088
rect 4844 13028 4848 13084
rect 4848 13028 4904 13084
rect 4904 13028 4908 13084
rect 4844 13024 4908 13028
rect 4924 13084 4988 13088
rect 4924 13028 4928 13084
rect 4928 13028 4984 13084
rect 4984 13028 4988 13084
rect 4924 13024 4988 13028
rect 12148 13084 12212 13088
rect 12148 13028 12152 13084
rect 12152 13028 12208 13084
rect 12208 13028 12212 13084
rect 12148 13024 12212 13028
rect 12228 13084 12292 13088
rect 12228 13028 12232 13084
rect 12232 13028 12288 13084
rect 12288 13028 12292 13084
rect 12228 13024 12292 13028
rect 12308 13084 12372 13088
rect 12308 13028 12312 13084
rect 12312 13028 12368 13084
rect 12368 13028 12372 13084
rect 12308 13024 12372 13028
rect 12388 13084 12452 13088
rect 12388 13028 12392 13084
rect 12392 13028 12448 13084
rect 12448 13028 12452 13084
rect 12388 13024 12452 13028
rect 19612 13084 19676 13088
rect 19612 13028 19616 13084
rect 19616 13028 19672 13084
rect 19672 13028 19676 13084
rect 19612 13024 19676 13028
rect 19692 13084 19756 13088
rect 19692 13028 19696 13084
rect 19696 13028 19752 13084
rect 19752 13028 19756 13084
rect 19692 13024 19756 13028
rect 19772 13084 19836 13088
rect 19772 13028 19776 13084
rect 19776 13028 19832 13084
rect 19832 13028 19836 13084
rect 19772 13024 19836 13028
rect 19852 13084 19916 13088
rect 19852 13028 19856 13084
rect 19856 13028 19912 13084
rect 19912 13028 19916 13084
rect 19852 13024 19916 13028
rect 8416 12540 8480 12544
rect 8416 12484 8420 12540
rect 8420 12484 8476 12540
rect 8476 12484 8480 12540
rect 8416 12480 8480 12484
rect 8496 12540 8560 12544
rect 8496 12484 8500 12540
rect 8500 12484 8556 12540
rect 8556 12484 8560 12540
rect 8496 12480 8560 12484
rect 8576 12540 8640 12544
rect 8576 12484 8580 12540
rect 8580 12484 8636 12540
rect 8636 12484 8640 12540
rect 8576 12480 8640 12484
rect 8656 12540 8720 12544
rect 8656 12484 8660 12540
rect 8660 12484 8716 12540
rect 8716 12484 8720 12540
rect 8656 12480 8720 12484
rect 15880 12540 15944 12544
rect 15880 12484 15884 12540
rect 15884 12484 15940 12540
rect 15940 12484 15944 12540
rect 15880 12480 15944 12484
rect 15960 12540 16024 12544
rect 15960 12484 15964 12540
rect 15964 12484 16020 12540
rect 16020 12484 16024 12540
rect 15960 12480 16024 12484
rect 16040 12540 16104 12544
rect 16040 12484 16044 12540
rect 16044 12484 16100 12540
rect 16100 12484 16104 12540
rect 16040 12480 16104 12484
rect 16120 12540 16184 12544
rect 16120 12484 16124 12540
rect 16124 12484 16180 12540
rect 16180 12484 16184 12540
rect 16120 12480 16184 12484
rect 4684 11996 4748 12000
rect 4684 11940 4688 11996
rect 4688 11940 4744 11996
rect 4744 11940 4748 11996
rect 4684 11936 4748 11940
rect 4764 11996 4828 12000
rect 4764 11940 4768 11996
rect 4768 11940 4824 11996
rect 4824 11940 4828 11996
rect 4764 11936 4828 11940
rect 4844 11996 4908 12000
rect 4844 11940 4848 11996
rect 4848 11940 4904 11996
rect 4904 11940 4908 11996
rect 4844 11936 4908 11940
rect 4924 11996 4988 12000
rect 4924 11940 4928 11996
rect 4928 11940 4984 11996
rect 4984 11940 4988 11996
rect 4924 11936 4988 11940
rect 12148 11996 12212 12000
rect 12148 11940 12152 11996
rect 12152 11940 12208 11996
rect 12208 11940 12212 11996
rect 12148 11936 12212 11940
rect 12228 11996 12292 12000
rect 12228 11940 12232 11996
rect 12232 11940 12288 11996
rect 12288 11940 12292 11996
rect 12228 11936 12292 11940
rect 12308 11996 12372 12000
rect 12308 11940 12312 11996
rect 12312 11940 12368 11996
rect 12368 11940 12372 11996
rect 12308 11936 12372 11940
rect 12388 11996 12452 12000
rect 12388 11940 12392 11996
rect 12392 11940 12448 11996
rect 12448 11940 12452 11996
rect 12388 11936 12452 11940
rect 19612 11996 19676 12000
rect 19612 11940 19616 11996
rect 19616 11940 19672 11996
rect 19672 11940 19676 11996
rect 19612 11936 19676 11940
rect 19692 11996 19756 12000
rect 19692 11940 19696 11996
rect 19696 11940 19752 11996
rect 19752 11940 19756 11996
rect 19692 11936 19756 11940
rect 19772 11996 19836 12000
rect 19772 11940 19776 11996
rect 19776 11940 19832 11996
rect 19832 11940 19836 11996
rect 19772 11936 19836 11940
rect 19852 11996 19916 12000
rect 19852 11940 19856 11996
rect 19856 11940 19912 11996
rect 19912 11940 19916 11996
rect 19852 11936 19916 11940
rect 8416 11452 8480 11456
rect 8416 11396 8420 11452
rect 8420 11396 8476 11452
rect 8476 11396 8480 11452
rect 8416 11392 8480 11396
rect 8496 11452 8560 11456
rect 8496 11396 8500 11452
rect 8500 11396 8556 11452
rect 8556 11396 8560 11452
rect 8496 11392 8560 11396
rect 8576 11452 8640 11456
rect 8576 11396 8580 11452
rect 8580 11396 8636 11452
rect 8636 11396 8640 11452
rect 8576 11392 8640 11396
rect 8656 11452 8720 11456
rect 8656 11396 8660 11452
rect 8660 11396 8716 11452
rect 8716 11396 8720 11452
rect 8656 11392 8720 11396
rect 15880 11452 15944 11456
rect 15880 11396 15884 11452
rect 15884 11396 15940 11452
rect 15940 11396 15944 11452
rect 15880 11392 15944 11396
rect 15960 11452 16024 11456
rect 15960 11396 15964 11452
rect 15964 11396 16020 11452
rect 16020 11396 16024 11452
rect 15960 11392 16024 11396
rect 16040 11452 16104 11456
rect 16040 11396 16044 11452
rect 16044 11396 16100 11452
rect 16100 11396 16104 11452
rect 16040 11392 16104 11396
rect 16120 11452 16184 11456
rect 16120 11396 16124 11452
rect 16124 11396 16180 11452
rect 16180 11396 16184 11452
rect 16120 11392 16184 11396
rect 20116 11112 20180 11116
rect 20116 11056 20166 11112
rect 20166 11056 20180 11112
rect 20116 11052 20180 11056
rect 20484 11112 20548 11116
rect 20484 11056 20498 11112
rect 20498 11056 20548 11112
rect 20484 11052 20548 11056
rect 4684 10908 4748 10912
rect 4684 10852 4688 10908
rect 4688 10852 4744 10908
rect 4744 10852 4748 10908
rect 4684 10848 4748 10852
rect 4764 10908 4828 10912
rect 4764 10852 4768 10908
rect 4768 10852 4824 10908
rect 4824 10852 4828 10908
rect 4764 10848 4828 10852
rect 4844 10908 4908 10912
rect 4844 10852 4848 10908
rect 4848 10852 4904 10908
rect 4904 10852 4908 10908
rect 4844 10848 4908 10852
rect 4924 10908 4988 10912
rect 4924 10852 4928 10908
rect 4928 10852 4984 10908
rect 4984 10852 4988 10908
rect 4924 10848 4988 10852
rect 12148 10908 12212 10912
rect 12148 10852 12152 10908
rect 12152 10852 12208 10908
rect 12208 10852 12212 10908
rect 12148 10848 12212 10852
rect 12228 10908 12292 10912
rect 12228 10852 12232 10908
rect 12232 10852 12288 10908
rect 12288 10852 12292 10908
rect 12228 10848 12292 10852
rect 12308 10908 12372 10912
rect 12308 10852 12312 10908
rect 12312 10852 12368 10908
rect 12368 10852 12372 10908
rect 12308 10848 12372 10852
rect 12388 10908 12452 10912
rect 12388 10852 12392 10908
rect 12392 10852 12448 10908
rect 12448 10852 12452 10908
rect 12388 10848 12452 10852
rect 19612 10908 19676 10912
rect 19612 10852 19616 10908
rect 19616 10852 19672 10908
rect 19672 10852 19676 10908
rect 19612 10848 19676 10852
rect 19692 10908 19756 10912
rect 19692 10852 19696 10908
rect 19696 10852 19752 10908
rect 19752 10852 19756 10908
rect 19692 10848 19756 10852
rect 19772 10908 19836 10912
rect 19772 10852 19776 10908
rect 19776 10852 19832 10908
rect 19832 10852 19836 10908
rect 19772 10848 19836 10852
rect 19852 10908 19916 10912
rect 19852 10852 19856 10908
rect 19856 10852 19912 10908
rect 19912 10852 19916 10908
rect 19852 10848 19916 10852
rect 8416 10364 8480 10368
rect 8416 10308 8420 10364
rect 8420 10308 8476 10364
rect 8476 10308 8480 10364
rect 8416 10304 8480 10308
rect 8496 10364 8560 10368
rect 8496 10308 8500 10364
rect 8500 10308 8556 10364
rect 8556 10308 8560 10364
rect 8496 10304 8560 10308
rect 8576 10364 8640 10368
rect 8576 10308 8580 10364
rect 8580 10308 8636 10364
rect 8636 10308 8640 10364
rect 8576 10304 8640 10308
rect 8656 10364 8720 10368
rect 8656 10308 8660 10364
rect 8660 10308 8716 10364
rect 8716 10308 8720 10364
rect 8656 10304 8720 10308
rect 15880 10364 15944 10368
rect 15880 10308 15884 10364
rect 15884 10308 15940 10364
rect 15940 10308 15944 10364
rect 15880 10304 15944 10308
rect 15960 10364 16024 10368
rect 15960 10308 15964 10364
rect 15964 10308 16020 10364
rect 16020 10308 16024 10364
rect 15960 10304 16024 10308
rect 16040 10364 16104 10368
rect 16040 10308 16044 10364
rect 16044 10308 16100 10364
rect 16100 10308 16104 10364
rect 16040 10304 16104 10308
rect 16120 10364 16184 10368
rect 16120 10308 16124 10364
rect 16124 10308 16180 10364
rect 16180 10308 16184 10364
rect 16120 10304 16184 10308
rect 4684 9820 4748 9824
rect 4684 9764 4688 9820
rect 4688 9764 4744 9820
rect 4744 9764 4748 9820
rect 4684 9760 4748 9764
rect 4764 9820 4828 9824
rect 4764 9764 4768 9820
rect 4768 9764 4824 9820
rect 4824 9764 4828 9820
rect 4764 9760 4828 9764
rect 4844 9820 4908 9824
rect 4844 9764 4848 9820
rect 4848 9764 4904 9820
rect 4904 9764 4908 9820
rect 4844 9760 4908 9764
rect 4924 9820 4988 9824
rect 4924 9764 4928 9820
rect 4928 9764 4984 9820
rect 4984 9764 4988 9820
rect 4924 9760 4988 9764
rect 12148 9820 12212 9824
rect 12148 9764 12152 9820
rect 12152 9764 12208 9820
rect 12208 9764 12212 9820
rect 12148 9760 12212 9764
rect 12228 9820 12292 9824
rect 12228 9764 12232 9820
rect 12232 9764 12288 9820
rect 12288 9764 12292 9820
rect 12228 9760 12292 9764
rect 12308 9820 12372 9824
rect 12308 9764 12312 9820
rect 12312 9764 12368 9820
rect 12368 9764 12372 9820
rect 12308 9760 12372 9764
rect 12388 9820 12452 9824
rect 12388 9764 12392 9820
rect 12392 9764 12448 9820
rect 12448 9764 12452 9820
rect 12388 9760 12452 9764
rect 19612 9820 19676 9824
rect 19612 9764 19616 9820
rect 19616 9764 19672 9820
rect 19672 9764 19676 9820
rect 19612 9760 19676 9764
rect 19692 9820 19756 9824
rect 19692 9764 19696 9820
rect 19696 9764 19752 9820
rect 19752 9764 19756 9820
rect 19692 9760 19756 9764
rect 19772 9820 19836 9824
rect 19772 9764 19776 9820
rect 19776 9764 19832 9820
rect 19832 9764 19836 9820
rect 19772 9760 19836 9764
rect 19852 9820 19916 9824
rect 19852 9764 19856 9820
rect 19856 9764 19912 9820
rect 19912 9764 19916 9820
rect 19852 9760 19916 9764
rect 8416 9276 8480 9280
rect 8416 9220 8420 9276
rect 8420 9220 8476 9276
rect 8476 9220 8480 9276
rect 8416 9216 8480 9220
rect 8496 9276 8560 9280
rect 8496 9220 8500 9276
rect 8500 9220 8556 9276
rect 8556 9220 8560 9276
rect 8496 9216 8560 9220
rect 8576 9276 8640 9280
rect 8576 9220 8580 9276
rect 8580 9220 8636 9276
rect 8636 9220 8640 9276
rect 8576 9216 8640 9220
rect 8656 9276 8720 9280
rect 8656 9220 8660 9276
rect 8660 9220 8716 9276
rect 8716 9220 8720 9276
rect 8656 9216 8720 9220
rect 15880 9276 15944 9280
rect 15880 9220 15884 9276
rect 15884 9220 15940 9276
rect 15940 9220 15944 9276
rect 15880 9216 15944 9220
rect 15960 9276 16024 9280
rect 15960 9220 15964 9276
rect 15964 9220 16020 9276
rect 16020 9220 16024 9276
rect 15960 9216 16024 9220
rect 16040 9276 16104 9280
rect 16040 9220 16044 9276
rect 16044 9220 16100 9276
rect 16100 9220 16104 9276
rect 16040 9216 16104 9220
rect 16120 9276 16184 9280
rect 16120 9220 16124 9276
rect 16124 9220 16180 9276
rect 16180 9220 16184 9276
rect 16120 9216 16184 9220
rect 4684 8732 4748 8736
rect 4684 8676 4688 8732
rect 4688 8676 4744 8732
rect 4744 8676 4748 8732
rect 4684 8672 4748 8676
rect 4764 8732 4828 8736
rect 4764 8676 4768 8732
rect 4768 8676 4824 8732
rect 4824 8676 4828 8732
rect 4764 8672 4828 8676
rect 4844 8732 4908 8736
rect 4844 8676 4848 8732
rect 4848 8676 4904 8732
rect 4904 8676 4908 8732
rect 4844 8672 4908 8676
rect 4924 8732 4988 8736
rect 4924 8676 4928 8732
rect 4928 8676 4984 8732
rect 4984 8676 4988 8732
rect 4924 8672 4988 8676
rect 12148 8732 12212 8736
rect 12148 8676 12152 8732
rect 12152 8676 12208 8732
rect 12208 8676 12212 8732
rect 12148 8672 12212 8676
rect 12228 8732 12292 8736
rect 12228 8676 12232 8732
rect 12232 8676 12288 8732
rect 12288 8676 12292 8732
rect 12228 8672 12292 8676
rect 12308 8732 12372 8736
rect 12308 8676 12312 8732
rect 12312 8676 12368 8732
rect 12368 8676 12372 8732
rect 12308 8672 12372 8676
rect 12388 8732 12452 8736
rect 12388 8676 12392 8732
rect 12392 8676 12448 8732
rect 12448 8676 12452 8732
rect 12388 8672 12452 8676
rect 19612 8732 19676 8736
rect 19612 8676 19616 8732
rect 19616 8676 19672 8732
rect 19672 8676 19676 8732
rect 19612 8672 19676 8676
rect 19692 8732 19756 8736
rect 19692 8676 19696 8732
rect 19696 8676 19752 8732
rect 19752 8676 19756 8732
rect 19692 8672 19756 8676
rect 19772 8732 19836 8736
rect 19772 8676 19776 8732
rect 19776 8676 19832 8732
rect 19832 8676 19836 8732
rect 19772 8672 19836 8676
rect 19852 8732 19916 8736
rect 19852 8676 19856 8732
rect 19856 8676 19912 8732
rect 19912 8676 19916 8732
rect 19852 8672 19916 8676
rect 8416 8188 8480 8192
rect 8416 8132 8420 8188
rect 8420 8132 8476 8188
rect 8476 8132 8480 8188
rect 8416 8128 8480 8132
rect 8496 8188 8560 8192
rect 8496 8132 8500 8188
rect 8500 8132 8556 8188
rect 8556 8132 8560 8188
rect 8496 8128 8560 8132
rect 8576 8188 8640 8192
rect 8576 8132 8580 8188
rect 8580 8132 8636 8188
rect 8636 8132 8640 8188
rect 8576 8128 8640 8132
rect 8656 8188 8720 8192
rect 8656 8132 8660 8188
rect 8660 8132 8716 8188
rect 8716 8132 8720 8188
rect 8656 8128 8720 8132
rect 15880 8188 15944 8192
rect 15880 8132 15884 8188
rect 15884 8132 15940 8188
rect 15940 8132 15944 8188
rect 15880 8128 15944 8132
rect 15960 8188 16024 8192
rect 15960 8132 15964 8188
rect 15964 8132 16020 8188
rect 16020 8132 16024 8188
rect 15960 8128 16024 8132
rect 16040 8188 16104 8192
rect 16040 8132 16044 8188
rect 16044 8132 16100 8188
rect 16100 8132 16104 8188
rect 16040 8128 16104 8132
rect 16120 8188 16184 8192
rect 16120 8132 16124 8188
rect 16124 8132 16180 8188
rect 16180 8132 16184 8188
rect 16120 8128 16184 8132
rect 4684 7644 4748 7648
rect 4684 7588 4688 7644
rect 4688 7588 4744 7644
rect 4744 7588 4748 7644
rect 4684 7584 4748 7588
rect 4764 7644 4828 7648
rect 4764 7588 4768 7644
rect 4768 7588 4824 7644
rect 4824 7588 4828 7644
rect 4764 7584 4828 7588
rect 4844 7644 4908 7648
rect 4844 7588 4848 7644
rect 4848 7588 4904 7644
rect 4904 7588 4908 7644
rect 4844 7584 4908 7588
rect 4924 7644 4988 7648
rect 4924 7588 4928 7644
rect 4928 7588 4984 7644
rect 4984 7588 4988 7644
rect 4924 7584 4988 7588
rect 12148 7644 12212 7648
rect 12148 7588 12152 7644
rect 12152 7588 12208 7644
rect 12208 7588 12212 7644
rect 12148 7584 12212 7588
rect 12228 7644 12292 7648
rect 12228 7588 12232 7644
rect 12232 7588 12288 7644
rect 12288 7588 12292 7644
rect 12228 7584 12292 7588
rect 12308 7644 12372 7648
rect 12308 7588 12312 7644
rect 12312 7588 12368 7644
rect 12368 7588 12372 7644
rect 12308 7584 12372 7588
rect 12388 7644 12452 7648
rect 12388 7588 12392 7644
rect 12392 7588 12448 7644
rect 12448 7588 12452 7644
rect 12388 7584 12452 7588
rect 19612 7644 19676 7648
rect 19612 7588 19616 7644
rect 19616 7588 19672 7644
rect 19672 7588 19676 7644
rect 19612 7584 19676 7588
rect 19692 7644 19756 7648
rect 19692 7588 19696 7644
rect 19696 7588 19752 7644
rect 19752 7588 19756 7644
rect 19692 7584 19756 7588
rect 19772 7644 19836 7648
rect 19772 7588 19776 7644
rect 19776 7588 19832 7644
rect 19832 7588 19836 7644
rect 19772 7584 19836 7588
rect 19852 7644 19916 7648
rect 19852 7588 19856 7644
rect 19856 7588 19912 7644
rect 19912 7588 19916 7644
rect 19852 7584 19916 7588
rect 8416 7100 8480 7104
rect 8416 7044 8420 7100
rect 8420 7044 8476 7100
rect 8476 7044 8480 7100
rect 8416 7040 8480 7044
rect 8496 7100 8560 7104
rect 8496 7044 8500 7100
rect 8500 7044 8556 7100
rect 8556 7044 8560 7100
rect 8496 7040 8560 7044
rect 8576 7100 8640 7104
rect 8576 7044 8580 7100
rect 8580 7044 8636 7100
rect 8636 7044 8640 7100
rect 8576 7040 8640 7044
rect 8656 7100 8720 7104
rect 8656 7044 8660 7100
rect 8660 7044 8716 7100
rect 8716 7044 8720 7100
rect 8656 7040 8720 7044
rect 15880 7100 15944 7104
rect 15880 7044 15884 7100
rect 15884 7044 15940 7100
rect 15940 7044 15944 7100
rect 15880 7040 15944 7044
rect 15960 7100 16024 7104
rect 15960 7044 15964 7100
rect 15964 7044 16020 7100
rect 16020 7044 16024 7100
rect 15960 7040 16024 7044
rect 16040 7100 16104 7104
rect 16040 7044 16044 7100
rect 16044 7044 16100 7100
rect 16100 7044 16104 7100
rect 16040 7040 16104 7044
rect 16120 7100 16184 7104
rect 16120 7044 16124 7100
rect 16124 7044 16180 7100
rect 16180 7044 16184 7100
rect 16120 7040 16184 7044
rect 4684 6556 4748 6560
rect 4684 6500 4688 6556
rect 4688 6500 4744 6556
rect 4744 6500 4748 6556
rect 4684 6496 4748 6500
rect 4764 6556 4828 6560
rect 4764 6500 4768 6556
rect 4768 6500 4824 6556
rect 4824 6500 4828 6556
rect 4764 6496 4828 6500
rect 4844 6556 4908 6560
rect 4844 6500 4848 6556
rect 4848 6500 4904 6556
rect 4904 6500 4908 6556
rect 4844 6496 4908 6500
rect 4924 6556 4988 6560
rect 4924 6500 4928 6556
rect 4928 6500 4984 6556
rect 4984 6500 4988 6556
rect 4924 6496 4988 6500
rect 12148 6556 12212 6560
rect 12148 6500 12152 6556
rect 12152 6500 12208 6556
rect 12208 6500 12212 6556
rect 12148 6496 12212 6500
rect 12228 6556 12292 6560
rect 12228 6500 12232 6556
rect 12232 6500 12288 6556
rect 12288 6500 12292 6556
rect 12228 6496 12292 6500
rect 12308 6556 12372 6560
rect 12308 6500 12312 6556
rect 12312 6500 12368 6556
rect 12368 6500 12372 6556
rect 12308 6496 12372 6500
rect 12388 6556 12452 6560
rect 12388 6500 12392 6556
rect 12392 6500 12448 6556
rect 12448 6500 12452 6556
rect 12388 6496 12452 6500
rect 19612 6556 19676 6560
rect 19612 6500 19616 6556
rect 19616 6500 19672 6556
rect 19672 6500 19676 6556
rect 19612 6496 19676 6500
rect 19692 6556 19756 6560
rect 19692 6500 19696 6556
rect 19696 6500 19752 6556
rect 19752 6500 19756 6556
rect 19692 6496 19756 6500
rect 19772 6556 19836 6560
rect 19772 6500 19776 6556
rect 19776 6500 19832 6556
rect 19832 6500 19836 6556
rect 19772 6496 19836 6500
rect 19852 6556 19916 6560
rect 19852 6500 19856 6556
rect 19856 6500 19912 6556
rect 19912 6500 19916 6556
rect 19852 6496 19916 6500
rect 8416 6012 8480 6016
rect 8416 5956 8420 6012
rect 8420 5956 8476 6012
rect 8476 5956 8480 6012
rect 8416 5952 8480 5956
rect 8496 6012 8560 6016
rect 8496 5956 8500 6012
rect 8500 5956 8556 6012
rect 8556 5956 8560 6012
rect 8496 5952 8560 5956
rect 8576 6012 8640 6016
rect 8576 5956 8580 6012
rect 8580 5956 8636 6012
rect 8636 5956 8640 6012
rect 8576 5952 8640 5956
rect 8656 6012 8720 6016
rect 8656 5956 8660 6012
rect 8660 5956 8716 6012
rect 8716 5956 8720 6012
rect 8656 5952 8720 5956
rect 15880 6012 15944 6016
rect 15880 5956 15884 6012
rect 15884 5956 15940 6012
rect 15940 5956 15944 6012
rect 15880 5952 15944 5956
rect 15960 6012 16024 6016
rect 15960 5956 15964 6012
rect 15964 5956 16020 6012
rect 16020 5956 16024 6012
rect 15960 5952 16024 5956
rect 16040 6012 16104 6016
rect 16040 5956 16044 6012
rect 16044 5956 16100 6012
rect 16100 5956 16104 6012
rect 16040 5952 16104 5956
rect 16120 6012 16184 6016
rect 16120 5956 16124 6012
rect 16124 5956 16180 6012
rect 16180 5956 16184 6012
rect 16120 5952 16184 5956
rect 4684 5468 4748 5472
rect 4684 5412 4688 5468
rect 4688 5412 4744 5468
rect 4744 5412 4748 5468
rect 4684 5408 4748 5412
rect 4764 5468 4828 5472
rect 4764 5412 4768 5468
rect 4768 5412 4824 5468
rect 4824 5412 4828 5468
rect 4764 5408 4828 5412
rect 4844 5468 4908 5472
rect 4844 5412 4848 5468
rect 4848 5412 4904 5468
rect 4904 5412 4908 5468
rect 4844 5408 4908 5412
rect 4924 5468 4988 5472
rect 4924 5412 4928 5468
rect 4928 5412 4984 5468
rect 4984 5412 4988 5468
rect 4924 5408 4988 5412
rect 12148 5468 12212 5472
rect 12148 5412 12152 5468
rect 12152 5412 12208 5468
rect 12208 5412 12212 5468
rect 12148 5408 12212 5412
rect 12228 5468 12292 5472
rect 12228 5412 12232 5468
rect 12232 5412 12288 5468
rect 12288 5412 12292 5468
rect 12228 5408 12292 5412
rect 12308 5468 12372 5472
rect 12308 5412 12312 5468
rect 12312 5412 12368 5468
rect 12368 5412 12372 5468
rect 12308 5408 12372 5412
rect 12388 5468 12452 5472
rect 12388 5412 12392 5468
rect 12392 5412 12448 5468
rect 12448 5412 12452 5468
rect 12388 5408 12452 5412
rect 19612 5468 19676 5472
rect 19612 5412 19616 5468
rect 19616 5412 19672 5468
rect 19672 5412 19676 5468
rect 19612 5408 19676 5412
rect 19692 5468 19756 5472
rect 19692 5412 19696 5468
rect 19696 5412 19752 5468
rect 19752 5412 19756 5468
rect 19692 5408 19756 5412
rect 19772 5468 19836 5472
rect 19772 5412 19776 5468
rect 19776 5412 19832 5468
rect 19832 5412 19836 5468
rect 19772 5408 19836 5412
rect 19852 5468 19916 5472
rect 19852 5412 19856 5468
rect 19856 5412 19912 5468
rect 19912 5412 19916 5468
rect 19852 5408 19916 5412
rect 8416 4924 8480 4928
rect 8416 4868 8420 4924
rect 8420 4868 8476 4924
rect 8476 4868 8480 4924
rect 8416 4864 8480 4868
rect 8496 4924 8560 4928
rect 8496 4868 8500 4924
rect 8500 4868 8556 4924
rect 8556 4868 8560 4924
rect 8496 4864 8560 4868
rect 8576 4924 8640 4928
rect 8576 4868 8580 4924
rect 8580 4868 8636 4924
rect 8636 4868 8640 4924
rect 8576 4864 8640 4868
rect 8656 4924 8720 4928
rect 8656 4868 8660 4924
rect 8660 4868 8716 4924
rect 8716 4868 8720 4924
rect 8656 4864 8720 4868
rect 15880 4924 15944 4928
rect 15880 4868 15884 4924
rect 15884 4868 15940 4924
rect 15940 4868 15944 4924
rect 15880 4864 15944 4868
rect 15960 4924 16024 4928
rect 15960 4868 15964 4924
rect 15964 4868 16020 4924
rect 16020 4868 16024 4924
rect 15960 4864 16024 4868
rect 16040 4924 16104 4928
rect 16040 4868 16044 4924
rect 16044 4868 16100 4924
rect 16100 4868 16104 4924
rect 16040 4864 16104 4868
rect 16120 4924 16184 4928
rect 16120 4868 16124 4924
rect 16124 4868 16180 4924
rect 16180 4868 16184 4924
rect 16120 4864 16184 4868
rect 4684 4380 4748 4384
rect 4684 4324 4688 4380
rect 4688 4324 4744 4380
rect 4744 4324 4748 4380
rect 4684 4320 4748 4324
rect 4764 4380 4828 4384
rect 4764 4324 4768 4380
rect 4768 4324 4824 4380
rect 4824 4324 4828 4380
rect 4764 4320 4828 4324
rect 4844 4380 4908 4384
rect 4844 4324 4848 4380
rect 4848 4324 4904 4380
rect 4904 4324 4908 4380
rect 4844 4320 4908 4324
rect 4924 4380 4988 4384
rect 4924 4324 4928 4380
rect 4928 4324 4984 4380
rect 4984 4324 4988 4380
rect 4924 4320 4988 4324
rect 12148 4380 12212 4384
rect 12148 4324 12152 4380
rect 12152 4324 12208 4380
rect 12208 4324 12212 4380
rect 12148 4320 12212 4324
rect 12228 4380 12292 4384
rect 12228 4324 12232 4380
rect 12232 4324 12288 4380
rect 12288 4324 12292 4380
rect 12228 4320 12292 4324
rect 12308 4380 12372 4384
rect 12308 4324 12312 4380
rect 12312 4324 12368 4380
rect 12368 4324 12372 4380
rect 12308 4320 12372 4324
rect 12388 4380 12452 4384
rect 12388 4324 12392 4380
rect 12392 4324 12448 4380
rect 12448 4324 12452 4380
rect 12388 4320 12452 4324
rect 19612 4380 19676 4384
rect 19612 4324 19616 4380
rect 19616 4324 19672 4380
rect 19672 4324 19676 4380
rect 19612 4320 19676 4324
rect 19692 4380 19756 4384
rect 19692 4324 19696 4380
rect 19696 4324 19752 4380
rect 19752 4324 19756 4380
rect 19692 4320 19756 4324
rect 19772 4380 19836 4384
rect 19772 4324 19776 4380
rect 19776 4324 19832 4380
rect 19832 4324 19836 4380
rect 19772 4320 19836 4324
rect 19852 4380 19916 4384
rect 19852 4324 19856 4380
rect 19856 4324 19912 4380
rect 19912 4324 19916 4380
rect 19852 4320 19916 4324
rect 8416 3836 8480 3840
rect 8416 3780 8420 3836
rect 8420 3780 8476 3836
rect 8476 3780 8480 3836
rect 8416 3776 8480 3780
rect 8496 3836 8560 3840
rect 8496 3780 8500 3836
rect 8500 3780 8556 3836
rect 8556 3780 8560 3836
rect 8496 3776 8560 3780
rect 8576 3836 8640 3840
rect 8576 3780 8580 3836
rect 8580 3780 8636 3836
rect 8636 3780 8640 3836
rect 8576 3776 8640 3780
rect 8656 3836 8720 3840
rect 8656 3780 8660 3836
rect 8660 3780 8716 3836
rect 8716 3780 8720 3836
rect 8656 3776 8720 3780
rect 15880 3836 15944 3840
rect 15880 3780 15884 3836
rect 15884 3780 15940 3836
rect 15940 3780 15944 3836
rect 15880 3776 15944 3780
rect 15960 3836 16024 3840
rect 15960 3780 15964 3836
rect 15964 3780 16020 3836
rect 16020 3780 16024 3836
rect 15960 3776 16024 3780
rect 16040 3836 16104 3840
rect 16040 3780 16044 3836
rect 16044 3780 16100 3836
rect 16100 3780 16104 3836
rect 16040 3776 16104 3780
rect 16120 3836 16184 3840
rect 16120 3780 16124 3836
rect 16124 3780 16180 3836
rect 16180 3780 16184 3836
rect 16120 3776 16184 3780
rect 4684 3292 4748 3296
rect 4684 3236 4688 3292
rect 4688 3236 4744 3292
rect 4744 3236 4748 3292
rect 4684 3232 4748 3236
rect 4764 3292 4828 3296
rect 4764 3236 4768 3292
rect 4768 3236 4824 3292
rect 4824 3236 4828 3292
rect 4764 3232 4828 3236
rect 4844 3292 4908 3296
rect 4844 3236 4848 3292
rect 4848 3236 4904 3292
rect 4904 3236 4908 3292
rect 4844 3232 4908 3236
rect 4924 3292 4988 3296
rect 4924 3236 4928 3292
rect 4928 3236 4984 3292
rect 4984 3236 4988 3292
rect 4924 3232 4988 3236
rect 12148 3292 12212 3296
rect 12148 3236 12152 3292
rect 12152 3236 12208 3292
rect 12208 3236 12212 3292
rect 12148 3232 12212 3236
rect 12228 3292 12292 3296
rect 12228 3236 12232 3292
rect 12232 3236 12288 3292
rect 12288 3236 12292 3292
rect 12228 3232 12292 3236
rect 12308 3292 12372 3296
rect 12308 3236 12312 3292
rect 12312 3236 12368 3292
rect 12368 3236 12372 3292
rect 12308 3232 12372 3236
rect 12388 3292 12452 3296
rect 12388 3236 12392 3292
rect 12392 3236 12448 3292
rect 12448 3236 12452 3292
rect 12388 3232 12452 3236
rect 19612 3292 19676 3296
rect 19612 3236 19616 3292
rect 19616 3236 19672 3292
rect 19672 3236 19676 3292
rect 19612 3232 19676 3236
rect 19692 3292 19756 3296
rect 19692 3236 19696 3292
rect 19696 3236 19752 3292
rect 19752 3236 19756 3292
rect 19692 3232 19756 3236
rect 19772 3292 19836 3296
rect 19772 3236 19776 3292
rect 19776 3236 19832 3292
rect 19832 3236 19836 3292
rect 19772 3232 19836 3236
rect 19852 3292 19916 3296
rect 19852 3236 19856 3292
rect 19856 3236 19912 3292
rect 19912 3236 19916 3292
rect 19852 3232 19916 3236
rect 8416 2748 8480 2752
rect 8416 2692 8420 2748
rect 8420 2692 8476 2748
rect 8476 2692 8480 2748
rect 8416 2688 8480 2692
rect 8496 2748 8560 2752
rect 8496 2692 8500 2748
rect 8500 2692 8556 2748
rect 8556 2692 8560 2748
rect 8496 2688 8560 2692
rect 8576 2748 8640 2752
rect 8576 2692 8580 2748
rect 8580 2692 8636 2748
rect 8636 2692 8640 2748
rect 8576 2688 8640 2692
rect 8656 2748 8720 2752
rect 8656 2692 8660 2748
rect 8660 2692 8716 2748
rect 8716 2692 8720 2748
rect 8656 2688 8720 2692
rect 15880 2748 15944 2752
rect 15880 2692 15884 2748
rect 15884 2692 15940 2748
rect 15940 2692 15944 2748
rect 15880 2688 15944 2692
rect 15960 2748 16024 2752
rect 15960 2692 15964 2748
rect 15964 2692 16020 2748
rect 16020 2692 16024 2748
rect 15960 2688 16024 2692
rect 16040 2748 16104 2752
rect 16040 2692 16044 2748
rect 16044 2692 16100 2748
rect 16100 2692 16104 2748
rect 16040 2688 16104 2692
rect 16120 2748 16184 2752
rect 16120 2692 16124 2748
rect 16124 2692 16180 2748
rect 16180 2692 16184 2748
rect 16120 2688 16184 2692
rect 4684 2204 4748 2208
rect 4684 2148 4688 2204
rect 4688 2148 4744 2204
rect 4744 2148 4748 2204
rect 4684 2144 4748 2148
rect 4764 2204 4828 2208
rect 4764 2148 4768 2204
rect 4768 2148 4824 2204
rect 4824 2148 4828 2204
rect 4764 2144 4828 2148
rect 4844 2204 4908 2208
rect 4844 2148 4848 2204
rect 4848 2148 4904 2204
rect 4904 2148 4908 2204
rect 4844 2144 4908 2148
rect 4924 2204 4988 2208
rect 4924 2148 4928 2204
rect 4928 2148 4984 2204
rect 4984 2148 4988 2204
rect 4924 2144 4988 2148
rect 12148 2204 12212 2208
rect 12148 2148 12152 2204
rect 12152 2148 12208 2204
rect 12208 2148 12212 2204
rect 12148 2144 12212 2148
rect 12228 2204 12292 2208
rect 12228 2148 12232 2204
rect 12232 2148 12288 2204
rect 12288 2148 12292 2204
rect 12228 2144 12292 2148
rect 12308 2204 12372 2208
rect 12308 2148 12312 2204
rect 12312 2148 12368 2204
rect 12368 2148 12372 2204
rect 12308 2144 12372 2148
rect 12388 2204 12452 2208
rect 12388 2148 12392 2204
rect 12392 2148 12448 2204
rect 12448 2148 12452 2204
rect 12388 2144 12452 2148
rect 19612 2204 19676 2208
rect 19612 2148 19616 2204
rect 19616 2148 19672 2204
rect 19672 2148 19676 2204
rect 19612 2144 19676 2148
rect 19692 2204 19756 2208
rect 19692 2148 19696 2204
rect 19696 2148 19752 2204
rect 19752 2148 19756 2204
rect 19692 2144 19756 2148
rect 19772 2204 19836 2208
rect 19772 2148 19776 2204
rect 19776 2148 19832 2204
rect 19832 2148 19836 2204
rect 19772 2144 19836 2148
rect 19852 2204 19916 2208
rect 19852 2148 19856 2204
rect 19856 2148 19912 2204
rect 19912 2148 19916 2204
rect 19852 2144 19916 2148
<< metal4 >>
rect 4676 21792 4996 22352
rect 4676 21728 4684 21792
rect 4748 21728 4764 21792
rect 4828 21728 4844 21792
rect 4908 21728 4924 21792
rect 4988 21728 4996 21792
rect 4676 20704 4996 21728
rect 4676 20640 4684 20704
rect 4748 20640 4764 20704
rect 4828 20640 4844 20704
rect 4908 20640 4924 20704
rect 4988 20640 4996 20704
rect 4676 19616 4996 20640
rect 4676 19552 4684 19616
rect 4748 19552 4764 19616
rect 4828 19552 4844 19616
rect 4908 19552 4924 19616
rect 4988 19552 4996 19616
rect 4676 18528 4996 19552
rect 4676 18464 4684 18528
rect 4748 18464 4764 18528
rect 4828 18464 4844 18528
rect 4908 18464 4924 18528
rect 4988 18464 4996 18528
rect 4676 17440 4996 18464
rect 4676 17376 4684 17440
rect 4748 17376 4764 17440
rect 4828 17376 4844 17440
rect 4908 17376 4924 17440
rect 4988 17376 4996 17440
rect 4676 16352 4996 17376
rect 4676 16288 4684 16352
rect 4748 16288 4764 16352
rect 4828 16288 4844 16352
rect 4908 16288 4924 16352
rect 4988 16288 4996 16352
rect 4676 15264 4996 16288
rect 4676 15200 4684 15264
rect 4748 15200 4764 15264
rect 4828 15200 4844 15264
rect 4908 15200 4924 15264
rect 4988 15200 4996 15264
rect 4676 14176 4996 15200
rect 4676 14112 4684 14176
rect 4748 14112 4764 14176
rect 4828 14112 4844 14176
rect 4908 14112 4924 14176
rect 4988 14112 4996 14176
rect 4676 13088 4996 14112
rect 4676 13024 4684 13088
rect 4748 13024 4764 13088
rect 4828 13024 4844 13088
rect 4908 13024 4924 13088
rect 4988 13024 4996 13088
rect 4676 12000 4996 13024
rect 4676 11936 4684 12000
rect 4748 11936 4764 12000
rect 4828 11936 4844 12000
rect 4908 11936 4924 12000
rect 4988 11936 4996 12000
rect 4676 10912 4996 11936
rect 4676 10848 4684 10912
rect 4748 10848 4764 10912
rect 4828 10848 4844 10912
rect 4908 10848 4924 10912
rect 4988 10848 4996 10912
rect 4676 9824 4996 10848
rect 4676 9760 4684 9824
rect 4748 9760 4764 9824
rect 4828 9760 4844 9824
rect 4908 9760 4924 9824
rect 4988 9760 4996 9824
rect 4676 8736 4996 9760
rect 4676 8672 4684 8736
rect 4748 8672 4764 8736
rect 4828 8672 4844 8736
rect 4908 8672 4924 8736
rect 4988 8672 4996 8736
rect 4676 7648 4996 8672
rect 4676 7584 4684 7648
rect 4748 7584 4764 7648
rect 4828 7584 4844 7648
rect 4908 7584 4924 7648
rect 4988 7584 4996 7648
rect 4676 6560 4996 7584
rect 4676 6496 4684 6560
rect 4748 6496 4764 6560
rect 4828 6496 4844 6560
rect 4908 6496 4924 6560
rect 4988 6496 4996 6560
rect 4676 5472 4996 6496
rect 4676 5408 4684 5472
rect 4748 5408 4764 5472
rect 4828 5408 4844 5472
rect 4908 5408 4924 5472
rect 4988 5408 4996 5472
rect 4676 4384 4996 5408
rect 4676 4320 4684 4384
rect 4748 4320 4764 4384
rect 4828 4320 4844 4384
rect 4908 4320 4924 4384
rect 4988 4320 4996 4384
rect 4676 3296 4996 4320
rect 4676 3232 4684 3296
rect 4748 3232 4764 3296
rect 4828 3232 4844 3296
rect 4908 3232 4924 3296
rect 4988 3232 4996 3296
rect 4676 2208 4996 3232
rect 4676 2144 4684 2208
rect 4748 2144 4764 2208
rect 4828 2144 4844 2208
rect 4908 2144 4924 2208
rect 4988 2144 4996 2208
rect 4676 2128 4996 2144
rect 8408 22336 8728 22352
rect 8408 22272 8416 22336
rect 8480 22272 8496 22336
rect 8560 22272 8576 22336
rect 8640 22272 8656 22336
rect 8720 22272 8728 22336
rect 8408 21248 8728 22272
rect 8408 21184 8416 21248
rect 8480 21184 8496 21248
rect 8560 21184 8576 21248
rect 8640 21184 8656 21248
rect 8720 21184 8728 21248
rect 8408 20160 8728 21184
rect 8408 20096 8416 20160
rect 8480 20096 8496 20160
rect 8560 20096 8576 20160
rect 8640 20096 8656 20160
rect 8720 20096 8728 20160
rect 8408 19072 8728 20096
rect 8408 19008 8416 19072
rect 8480 19008 8496 19072
rect 8560 19008 8576 19072
rect 8640 19008 8656 19072
rect 8720 19008 8728 19072
rect 8408 17984 8728 19008
rect 8408 17920 8416 17984
rect 8480 17920 8496 17984
rect 8560 17920 8576 17984
rect 8640 17920 8656 17984
rect 8720 17920 8728 17984
rect 8408 16896 8728 17920
rect 8408 16832 8416 16896
rect 8480 16832 8496 16896
rect 8560 16832 8576 16896
rect 8640 16832 8656 16896
rect 8720 16832 8728 16896
rect 8408 15808 8728 16832
rect 8408 15744 8416 15808
rect 8480 15744 8496 15808
rect 8560 15744 8576 15808
rect 8640 15744 8656 15808
rect 8720 15744 8728 15808
rect 8408 14720 8728 15744
rect 8408 14656 8416 14720
rect 8480 14656 8496 14720
rect 8560 14656 8576 14720
rect 8640 14656 8656 14720
rect 8720 14656 8728 14720
rect 8408 13632 8728 14656
rect 8408 13568 8416 13632
rect 8480 13568 8496 13632
rect 8560 13568 8576 13632
rect 8640 13568 8656 13632
rect 8720 13568 8728 13632
rect 8408 12544 8728 13568
rect 8408 12480 8416 12544
rect 8480 12480 8496 12544
rect 8560 12480 8576 12544
rect 8640 12480 8656 12544
rect 8720 12480 8728 12544
rect 8408 11456 8728 12480
rect 8408 11392 8416 11456
rect 8480 11392 8496 11456
rect 8560 11392 8576 11456
rect 8640 11392 8656 11456
rect 8720 11392 8728 11456
rect 8408 10368 8728 11392
rect 8408 10304 8416 10368
rect 8480 10304 8496 10368
rect 8560 10304 8576 10368
rect 8640 10304 8656 10368
rect 8720 10304 8728 10368
rect 8408 9280 8728 10304
rect 8408 9216 8416 9280
rect 8480 9216 8496 9280
rect 8560 9216 8576 9280
rect 8640 9216 8656 9280
rect 8720 9216 8728 9280
rect 8408 8192 8728 9216
rect 8408 8128 8416 8192
rect 8480 8128 8496 8192
rect 8560 8128 8576 8192
rect 8640 8128 8656 8192
rect 8720 8128 8728 8192
rect 8408 7104 8728 8128
rect 8408 7040 8416 7104
rect 8480 7040 8496 7104
rect 8560 7040 8576 7104
rect 8640 7040 8656 7104
rect 8720 7040 8728 7104
rect 8408 6016 8728 7040
rect 8408 5952 8416 6016
rect 8480 5952 8496 6016
rect 8560 5952 8576 6016
rect 8640 5952 8656 6016
rect 8720 5952 8728 6016
rect 8408 4928 8728 5952
rect 8408 4864 8416 4928
rect 8480 4864 8496 4928
rect 8560 4864 8576 4928
rect 8640 4864 8656 4928
rect 8720 4864 8728 4928
rect 8408 3840 8728 4864
rect 8408 3776 8416 3840
rect 8480 3776 8496 3840
rect 8560 3776 8576 3840
rect 8640 3776 8656 3840
rect 8720 3776 8728 3840
rect 8408 2752 8728 3776
rect 8408 2688 8416 2752
rect 8480 2688 8496 2752
rect 8560 2688 8576 2752
rect 8640 2688 8656 2752
rect 8720 2688 8728 2752
rect 8408 2128 8728 2688
rect 12140 21792 12460 22352
rect 12140 21728 12148 21792
rect 12212 21728 12228 21792
rect 12292 21728 12308 21792
rect 12372 21728 12388 21792
rect 12452 21728 12460 21792
rect 12140 20704 12460 21728
rect 12140 20640 12148 20704
rect 12212 20640 12228 20704
rect 12292 20640 12308 20704
rect 12372 20640 12388 20704
rect 12452 20640 12460 20704
rect 12140 19616 12460 20640
rect 12140 19552 12148 19616
rect 12212 19552 12228 19616
rect 12292 19552 12308 19616
rect 12372 19552 12388 19616
rect 12452 19552 12460 19616
rect 12140 18528 12460 19552
rect 12140 18464 12148 18528
rect 12212 18464 12228 18528
rect 12292 18464 12308 18528
rect 12372 18464 12388 18528
rect 12452 18464 12460 18528
rect 12140 17440 12460 18464
rect 12140 17376 12148 17440
rect 12212 17376 12228 17440
rect 12292 17376 12308 17440
rect 12372 17376 12388 17440
rect 12452 17376 12460 17440
rect 12140 16352 12460 17376
rect 12140 16288 12148 16352
rect 12212 16288 12228 16352
rect 12292 16288 12308 16352
rect 12372 16288 12388 16352
rect 12452 16288 12460 16352
rect 12140 15264 12460 16288
rect 12140 15200 12148 15264
rect 12212 15200 12228 15264
rect 12292 15200 12308 15264
rect 12372 15200 12388 15264
rect 12452 15200 12460 15264
rect 12140 14176 12460 15200
rect 12140 14112 12148 14176
rect 12212 14112 12228 14176
rect 12292 14112 12308 14176
rect 12372 14112 12388 14176
rect 12452 14112 12460 14176
rect 12140 13088 12460 14112
rect 12140 13024 12148 13088
rect 12212 13024 12228 13088
rect 12292 13024 12308 13088
rect 12372 13024 12388 13088
rect 12452 13024 12460 13088
rect 12140 12000 12460 13024
rect 12140 11936 12148 12000
rect 12212 11936 12228 12000
rect 12292 11936 12308 12000
rect 12372 11936 12388 12000
rect 12452 11936 12460 12000
rect 12140 10912 12460 11936
rect 12140 10848 12148 10912
rect 12212 10848 12228 10912
rect 12292 10848 12308 10912
rect 12372 10848 12388 10912
rect 12452 10848 12460 10912
rect 12140 9824 12460 10848
rect 12140 9760 12148 9824
rect 12212 9760 12228 9824
rect 12292 9760 12308 9824
rect 12372 9760 12388 9824
rect 12452 9760 12460 9824
rect 12140 8736 12460 9760
rect 12140 8672 12148 8736
rect 12212 8672 12228 8736
rect 12292 8672 12308 8736
rect 12372 8672 12388 8736
rect 12452 8672 12460 8736
rect 12140 7648 12460 8672
rect 12140 7584 12148 7648
rect 12212 7584 12228 7648
rect 12292 7584 12308 7648
rect 12372 7584 12388 7648
rect 12452 7584 12460 7648
rect 12140 6560 12460 7584
rect 12140 6496 12148 6560
rect 12212 6496 12228 6560
rect 12292 6496 12308 6560
rect 12372 6496 12388 6560
rect 12452 6496 12460 6560
rect 12140 5472 12460 6496
rect 12140 5408 12148 5472
rect 12212 5408 12228 5472
rect 12292 5408 12308 5472
rect 12372 5408 12388 5472
rect 12452 5408 12460 5472
rect 12140 4384 12460 5408
rect 12140 4320 12148 4384
rect 12212 4320 12228 4384
rect 12292 4320 12308 4384
rect 12372 4320 12388 4384
rect 12452 4320 12460 4384
rect 12140 3296 12460 4320
rect 12140 3232 12148 3296
rect 12212 3232 12228 3296
rect 12292 3232 12308 3296
rect 12372 3232 12388 3296
rect 12452 3232 12460 3296
rect 12140 2208 12460 3232
rect 12140 2144 12148 2208
rect 12212 2144 12228 2208
rect 12292 2144 12308 2208
rect 12372 2144 12388 2208
rect 12452 2144 12460 2208
rect 12140 2128 12460 2144
rect 15872 22336 16192 22352
rect 15872 22272 15880 22336
rect 15944 22272 15960 22336
rect 16024 22272 16040 22336
rect 16104 22272 16120 22336
rect 16184 22272 16192 22336
rect 15872 21248 16192 22272
rect 15872 21184 15880 21248
rect 15944 21184 15960 21248
rect 16024 21184 16040 21248
rect 16104 21184 16120 21248
rect 16184 21184 16192 21248
rect 15872 20160 16192 21184
rect 15872 20096 15880 20160
rect 15944 20096 15960 20160
rect 16024 20096 16040 20160
rect 16104 20096 16120 20160
rect 16184 20096 16192 20160
rect 15872 19072 16192 20096
rect 15872 19008 15880 19072
rect 15944 19008 15960 19072
rect 16024 19008 16040 19072
rect 16104 19008 16120 19072
rect 16184 19008 16192 19072
rect 15872 17984 16192 19008
rect 15872 17920 15880 17984
rect 15944 17920 15960 17984
rect 16024 17920 16040 17984
rect 16104 17920 16120 17984
rect 16184 17920 16192 17984
rect 15872 16896 16192 17920
rect 15872 16832 15880 16896
rect 15944 16832 15960 16896
rect 16024 16832 16040 16896
rect 16104 16832 16120 16896
rect 16184 16832 16192 16896
rect 15872 15808 16192 16832
rect 15872 15744 15880 15808
rect 15944 15744 15960 15808
rect 16024 15744 16040 15808
rect 16104 15744 16120 15808
rect 16184 15744 16192 15808
rect 15872 14720 16192 15744
rect 15872 14656 15880 14720
rect 15944 14656 15960 14720
rect 16024 14656 16040 14720
rect 16104 14656 16120 14720
rect 16184 14656 16192 14720
rect 15872 13632 16192 14656
rect 15872 13568 15880 13632
rect 15944 13568 15960 13632
rect 16024 13568 16040 13632
rect 16104 13568 16120 13632
rect 16184 13568 16192 13632
rect 15872 12544 16192 13568
rect 15872 12480 15880 12544
rect 15944 12480 15960 12544
rect 16024 12480 16040 12544
rect 16104 12480 16120 12544
rect 16184 12480 16192 12544
rect 15872 11456 16192 12480
rect 15872 11392 15880 11456
rect 15944 11392 15960 11456
rect 16024 11392 16040 11456
rect 16104 11392 16120 11456
rect 16184 11392 16192 11456
rect 15872 10368 16192 11392
rect 15872 10304 15880 10368
rect 15944 10304 15960 10368
rect 16024 10304 16040 10368
rect 16104 10304 16120 10368
rect 16184 10304 16192 10368
rect 15872 9280 16192 10304
rect 15872 9216 15880 9280
rect 15944 9216 15960 9280
rect 16024 9216 16040 9280
rect 16104 9216 16120 9280
rect 16184 9216 16192 9280
rect 15872 8192 16192 9216
rect 15872 8128 15880 8192
rect 15944 8128 15960 8192
rect 16024 8128 16040 8192
rect 16104 8128 16120 8192
rect 16184 8128 16192 8192
rect 15872 7104 16192 8128
rect 15872 7040 15880 7104
rect 15944 7040 15960 7104
rect 16024 7040 16040 7104
rect 16104 7040 16120 7104
rect 16184 7040 16192 7104
rect 15872 6016 16192 7040
rect 15872 5952 15880 6016
rect 15944 5952 15960 6016
rect 16024 5952 16040 6016
rect 16104 5952 16120 6016
rect 16184 5952 16192 6016
rect 15872 4928 16192 5952
rect 15872 4864 15880 4928
rect 15944 4864 15960 4928
rect 16024 4864 16040 4928
rect 16104 4864 16120 4928
rect 16184 4864 16192 4928
rect 15872 3840 16192 4864
rect 15872 3776 15880 3840
rect 15944 3776 15960 3840
rect 16024 3776 16040 3840
rect 16104 3776 16120 3840
rect 16184 3776 16192 3840
rect 15872 2752 16192 3776
rect 15872 2688 15880 2752
rect 15944 2688 15960 2752
rect 16024 2688 16040 2752
rect 16104 2688 16120 2752
rect 16184 2688 16192 2752
rect 15872 2128 16192 2688
rect 19604 21792 19924 22352
rect 19604 21728 19612 21792
rect 19676 21728 19692 21792
rect 19756 21728 19772 21792
rect 19836 21728 19852 21792
rect 19916 21728 19924 21792
rect 19604 20704 19924 21728
rect 19604 20640 19612 20704
rect 19676 20640 19692 20704
rect 19756 20640 19772 20704
rect 19836 20640 19852 20704
rect 19916 20640 19924 20704
rect 19604 19616 19924 20640
rect 19604 19552 19612 19616
rect 19676 19552 19692 19616
rect 19756 19552 19772 19616
rect 19836 19552 19852 19616
rect 19916 19552 19924 19616
rect 19604 18528 19924 19552
rect 19604 18464 19612 18528
rect 19676 18464 19692 18528
rect 19756 18464 19772 18528
rect 19836 18464 19852 18528
rect 19916 18464 19924 18528
rect 19604 17440 19924 18464
rect 19604 17376 19612 17440
rect 19676 17376 19692 17440
rect 19756 17376 19772 17440
rect 19836 17376 19852 17440
rect 19916 17376 19924 17440
rect 19604 16352 19924 17376
rect 19604 16288 19612 16352
rect 19676 16288 19692 16352
rect 19756 16288 19772 16352
rect 19836 16288 19852 16352
rect 19916 16288 19924 16352
rect 19604 15264 19924 16288
rect 20115 15740 20181 15741
rect 20115 15676 20116 15740
rect 20180 15676 20181 15740
rect 20115 15675 20181 15676
rect 19604 15200 19612 15264
rect 19676 15200 19692 15264
rect 19756 15200 19772 15264
rect 19836 15200 19852 15264
rect 19916 15200 19924 15264
rect 19604 14176 19924 15200
rect 19604 14112 19612 14176
rect 19676 14112 19692 14176
rect 19756 14112 19772 14176
rect 19836 14112 19852 14176
rect 19916 14112 19924 14176
rect 19604 13088 19924 14112
rect 19604 13024 19612 13088
rect 19676 13024 19692 13088
rect 19756 13024 19772 13088
rect 19836 13024 19852 13088
rect 19916 13024 19924 13088
rect 19604 12000 19924 13024
rect 19604 11936 19612 12000
rect 19676 11936 19692 12000
rect 19756 11936 19772 12000
rect 19836 11936 19852 12000
rect 19916 11936 19924 12000
rect 19604 10912 19924 11936
rect 20118 11117 20178 15675
rect 20483 13292 20549 13293
rect 20483 13228 20484 13292
rect 20548 13228 20549 13292
rect 20483 13227 20549 13228
rect 20486 11117 20546 13227
rect 20115 11116 20181 11117
rect 20115 11052 20116 11116
rect 20180 11052 20181 11116
rect 20115 11051 20181 11052
rect 20483 11116 20549 11117
rect 20483 11052 20484 11116
rect 20548 11052 20549 11116
rect 20483 11051 20549 11052
rect 19604 10848 19612 10912
rect 19676 10848 19692 10912
rect 19756 10848 19772 10912
rect 19836 10848 19852 10912
rect 19916 10848 19924 10912
rect 19604 9824 19924 10848
rect 19604 9760 19612 9824
rect 19676 9760 19692 9824
rect 19756 9760 19772 9824
rect 19836 9760 19852 9824
rect 19916 9760 19924 9824
rect 19604 8736 19924 9760
rect 19604 8672 19612 8736
rect 19676 8672 19692 8736
rect 19756 8672 19772 8736
rect 19836 8672 19852 8736
rect 19916 8672 19924 8736
rect 19604 7648 19924 8672
rect 19604 7584 19612 7648
rect 19676 7584 19692 7648
rect 19756 7584 19772 7648
rect 19836 7584 19852 7648
rect 19916 7584 19924 7648
rect 19604 6560 19924 7584
rect 19604 6496 19612 6560
rect 19676 6496 19692 6560
rect 19756 6496 19772 6560
rect 19836 6496 19852 6560
rect 19916 6496 19924 6560
rect 19604 5472 19924 6496
rect 19604 5408 19612 5472
rect 19676 5408 19692 5472
rect 19756 5408 19772 5472
rect 19836 5408 19852 5472
rect 19916 5408 19924 5472
rect 19604 4384 19924 5408
rect 19604 4320 19612 4384
rect 19676 4320 19692 4384
rect 19756 4320 19772 4384
rect 19836 4320 19852 4384
rect 19916 4320 19924 4384
rect 19604 3296 19924 4320
rect 19604 3232 19612 3296
rect 19676 3232 19692 3296
rect 19756 3232 19772 3296
rect 19836 3232 19852 3296
rect 19916 3232 19924 3296
rect 19604 2208 19924 3232
rect 19604 2144 19612 2208
rect 19676 2144 19692 2208
rect 19756 2144 19772 2208
rect 19836 2144 19852 2208
rect 19916 2144 19924 2208
rect 19604 2128 19924 2144
use sky130_fd_sc_hd__fill_1  FILLER_1_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1656 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9
timestamp 1624635492
transform 1 0 1932 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output52 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 1656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2392 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2300 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1624635492
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _66_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2484 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2944 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_14
timestamp 1624635492
transform 1 0 2392 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26
timestamp 1624635492
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_30
timestamp 1624635492
transform 1 0 3864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42
timestamp 1624635492
transform 1 0 4968 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1624635492
transform 1 0 4048 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5152 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _64_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output47
timestamp 1624635492
transform -1 0 6440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_59
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_58
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_71
timestamp 1624635492
transform 1 0 7636 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_88
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_70
timestamp 1624635492
transform 1 0 7544 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_82
timestamp 1624635492
transform 1 0 8648 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output42
timestamp 1624635492
transform -1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output42_A
timestamp 1624635492
transform -1 0 10764 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_96
timestamp 1624635492
transform 1 0 9936 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_105
timestamp 1624635492
transform 1 0 10764 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1624635492
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_94
timestamp 1624635492
transform 1 0 9752 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_106
timestamp 1624635492
transform 1 0 10856 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_117
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_129
timestamp 1624635492
transform 1 0 12972 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_115
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_127
timestamp 1624635492
transform 1 0 12788 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1624635492
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1624635492
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_151
timestamp 1624635492
transform 1 0 14996 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_139
timestamp 1624635492
transform 1 0 13892 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_151
timestamp 1624635492
transform 1 0 14996 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1624635492
transform 1 0 17204 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output61_A
timestamp 1624635492
transform -1 0 17112 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_163
timestamp 1624635492
transform 1 0 16100 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_171
timestamp 1624635492
transform 1 0 16836 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_163
timestamp 1624635492
transform 1 0 16100 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 19136 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1624635492
transform -1 0 18952 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 18400 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_204
timestamp 1624635492
transform 1 0 19872 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output59_A
timestamp 1624635492
transform -1 0 19320 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output57_A
timestamp 1624635492
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output55_A
timestamp 1624635492
transform -1 0 19504 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  output51
timestamp 1624635492
transform 1 0 19504 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1624635492
transform -1 0 20240 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1624635492
transform -1 0 20884 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1624635492
transform 1 0 20884 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1624635492
transform 1 0 20608 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output55
timestamp 1624635492
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output59
timestamp 1624635492
transform 1 0 21712 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output61
timestamp 1624635492
transform 1 0 20240 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform 1 0 22540 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1624635492
transform -1 0 22724 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 23460 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 23460 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output53
timestamp 1624635492
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output57
timestamp 1624635492
transform 1 0 22816 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_235
timestamp 1624635492
transform 1 0 22724 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1624635492
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_30
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_42
timestamp 1624635492
transform 1 0 4968 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_54
timestamp 1624635492
transform 1 0 6072 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_66
timestamp 1624635492
transform 1 0 7176 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_78
timestamp 1624635492
transform 1 0 8280 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_87
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_99
timestamp 1624635492
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_111
timestamp 1624635492
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1624635492
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_135
timestamp 1624635492
transform 1 0 13524 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_144
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_156
timestamp 1624635492
transform 1 0 15456 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform -1 0 17940 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output63_A
timestamp 1624635492
transform -1 0 16468 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_164
timestamp 1624635492
transform 1 0 16192 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1624635492
transform 1 0 19964 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1624635492
transform 1 0 17940 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output63
timestamp 1624635492
transform 1 0 19596 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_199
timestamp 1624635492
transform 1 0 19412 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1624635492
transform 1 0 21436 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1624635492
transform 1 0 22908 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 23460 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1624635492
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1624635492
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1624635492
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_51
timestamp 1624635492
transform 1 0 5796 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1624635492
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1624635492
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1624635492
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1624635492
transform 1 0 9752 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_106
timestamp 1624635492
transform 1 0 10856 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1624635492
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1624635492
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_151
timestamp 1624635492
transform 1 0 14996 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_159
timestamp 1624635492
transform 1 0 15732 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1624635492
transform 1 0 16008 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output67_A
timestamp 1624635492
transform -1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1624635492
transform 1 0 18400 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output67
timestamp 1624635492
transform 1 0 19872 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1624635492
transform 1 0 20608 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output65
timestamp 1624635492
transform 1 0 20240 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1624635492
transform 1 0 22172 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 23460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1624635492
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1624635492
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1624635492
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1624635492
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1624635492
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1624635492
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1624635492
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_99
timestamp 1624635492
transform 1 0 10212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1624635492
transform 1 0 11316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1624635492
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1624635492
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_156
timestamp 1624635492
transform 1 0 15456 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1624635492
transform -1 0 18676 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1624635492
transform -1 0 16376 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 17848 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_4_162
timestamp 1624635492
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1624635492
transform 1 0 18676 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1624635492
transform 1 0 19596 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1624635492
transform -1 0 22908 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output48
timestamp 1624635492
transform 1 0 21068 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform 1 0 22908 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 23460 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1624635492
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1624635492
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1624635492
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_51
timestamp 1624635492
transform 1 0 5796 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1624635492
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1624635492
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1624635492
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1624635492
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1624635492
transform -1 0 13708 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_5_115
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1624635492
transform 1 0 13708 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1624635492
transform 1 0 14812 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_157
timestamp 1624635492
transform 1 0 15548 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1624635492
transform 1 0 16100 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform -1 0 16836 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16928 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 16100 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1624635492
transform 1 0 16376 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1624635492
transform -1 0 19504 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18400 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1624635492
transform -1 0 20332 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1624635492
transform 1 0 20332 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1624635492
transform -1 0 21988 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_227
timestamp 1624635492
transform 1 0 21988 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1624635492
transform 1 0 22172 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 23460 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output48_A
timestamp 1624635492
transform -1 0 23184 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1624635492
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1624635492
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1624635492
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1624635492
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1624635492
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1624635492
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1624635492
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1624635492
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1624635492
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1624635492
transform 1 0 8648 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1624635492
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_87
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1624635492
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1624635492
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1624635492
transform 1 0 10120 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1624635492
transform 1 0 11132 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1624635492
transform 1 0 12604 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1624635492
transform 1 0 13156 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform -1 0 14628 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14628 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 15824 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 14904 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1624635492
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_150
timestamp 1624635492
transform 1 0 14904 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18216 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15916 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 16928 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 16100 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_6_160
timestamp 1624635492
transform 1 0 15824 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_170
timestamp 1624635492
transform 1 0 16744 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1624635492
transform -1 0 19504 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform -1 0 18676 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 19596 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 19412 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 19412 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform -1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output65_A
timestamp 1624635492
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1624635492
transform 1 0 20884 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 22080 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 21068 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1624635492
transform -1 0 23000 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 22080 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 22172 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 23460 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 23460 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_238
timestamp 1624635492
transform 1 0 23000 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_238
timestamp 1624635492
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1624635492
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1624635492
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1624635492
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1624635492
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1624635492
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1624635492
transform -1 0 10580 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1624635492
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1624635492
transform -1 0 11408 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1624635492
transform 1 0 11408 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1624635492
transform 1 0 12236 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1624635492
transform 1 0 13064 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform -1 0 14260 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1624635492
transform 1 0 13892 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15824 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 18768 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1624635492
transform 1 0 18768 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output44
timestamp 1624635492
transform 1 0 19688 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1624635492
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_201
timestamp 1624635492
transform 1 0 19596 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1624635492
transform -1 0 20884 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 23092 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  output49
timestamp 1624635492
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform -1 0 21344 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_220
timestamp 1624635492
transform 1 0 21344 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 23460 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_239
timestamp 1624635492
transform 1 0 23092 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1624635492
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1624635492
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1624635492
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51
timestamp 1624635492
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1624635492
transform 1 0 9108 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1624635492
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1624635492
transform 1 0 8648 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_86
timestamp 1624635492
transform 1 0 9016 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1624635492
transform -1 0 11408 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_112
timestamp 1624635492
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1624635492
transform 1 0 11960 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1624635492
transform -1 0 13616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1624635492
transform -1 0 11960 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1624635492
transform -1 0 14076 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1624635492
transform -1 0 14904 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 15732 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_4  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1624635492
transform 1 0 17756 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 16928 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 19780 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1624635492
transform 1 0 19964 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 19964 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_E_FTB01
timestamp 1624635492
transform 1 0 21804 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 20332 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 23000 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 23460 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_E_FTB01_A
timestamp 1624635492
transform -1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1624635492
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624635492
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1624635492
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  Test_en_FTB00
timestamp 1624635492
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1624635492
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1624635492
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1624635492
transform -1 0 10580 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_FTB00_A
timestamp 1624635492
transform 1 0 8464 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_82
timestamp 1624635492
transform 1 0 8648 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1624635492
transform -1 0 11408 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1624635492
transform -1 0 11684 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12972 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1624635492
transform -1 0 13800 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1624635492
transform -1 0 12144 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_115
timestamp 1624635492
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14536 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform -1 0 14260 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 14352 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1624635492
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 16468 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1624635492
transform -1 0 19872 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1624635492
transform -1 0 18676 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 19872 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 19504 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 22080 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 22080 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 23460 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_W_FTB01
timestamp 1624635492
transform 1 0 1748 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_W_FTB01_A
timestamp 1624635492
transform -1 0 2208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_12
timestamp 1624635492
transform 1 0 2208 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_24
timestamp 1624635492
transform 1 0 3312 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_36
timestamp 1624635492
transform 1 0 4416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1624635492
transform 1 0 5520 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_56
timestamp 1624635492
transform 1 0 6256 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform -1 0 10304 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1624635492
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp 1624635492
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1624635492
transform -1 0 11132 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform -1 0 11592 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1624635492
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1624635492
transform 1 0 13156 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 13156 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1624635492
transform 1 0 15548 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 15548 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_140
timestamp 1624635492
transform 1 0 13984 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform -1 0 17204 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 17204 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1624635492
transform -1 0 16836 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1624635492
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 18308 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1624635492
transform -1 0 20608 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 20608 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_208
timestamp 1624635492
transform 1 0 20240 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 22172 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 23460 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_238
timestamp 1624635492
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1624635492
transform -1 0 1656 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 1840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_8
timestamp 1624635492
transform 1 0 1840 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1624635492
transform 1 0 2944 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_28
timestamp 1624635492
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1624635492
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1624635492
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_66
timestamp 1624635492
transform 1 0 7176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1624635492
transform 1 0 9108 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1624635492
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11408 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_12_112
timestamp 1624635492
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1624635492
transform -1 0 13984 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11684 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 15824 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_140
timestamp 1624635492
transform 1 0 13984 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 18032 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 15824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 16284 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1624635492
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 19504 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 20424 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 21528 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_4  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 21528 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 23460 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_238
timestamp 1624635492
transform 1 0 23000 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1624635492
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1624635492
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1624635492
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1624635492
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1624635492
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1624635492
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1624635492
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1624635492
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_66
timestamp 1624635492
transform 1 0 7176 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1624635492
transform -1 0 8740 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1624635492
transform -1 0 10120 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1624635492
transform -1 0 9016 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_70
timestamp 1624635492
transform 1 0 7544 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_83
timestamp 1624635492
transform 1 0 8740 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_87
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1624635492
transform 1 0 10120 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11592 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 10120 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_98
timestamp 1624635492
transform 1 0 10120 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_104
timestamp 1624635492
transform 1 0 10672 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_114
timestamp 1624635492
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 13616 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 13248 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 13248 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14260 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1624635492
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_132
timestamp 1624635492
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_6  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform -1 0 15180 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 14628 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14628 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 17204 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_153
timestamp 1624635492
transform 1 0 15180 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 17388 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17204 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1624635492
transform -1 0 16836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 16560 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform 1 0 17204 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18676 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 19596 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 20332 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624635492
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_198
timestamp 1624635492
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1624635492
transform -1 0 20608 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 21068 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 20608 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624635492
transform 1 0 22080 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 22172 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_E_FTB01
timestamp 1624635492
transform -1 0 23184 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 23460 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 23460 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_E_FTB01_A
timestamp 1624635492
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_233
timestamp 1624635492
transform 1 0 22540 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1624635492
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1624635492
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1624635492
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1624635492
transform -1 0 8648 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1624635492
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_58
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1624635492
transform 1 0 9200 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 9200 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_82
timestamp 1624635492
transform 1 0 8648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform -1 0 11500 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1624635492
transform 1 0 11500 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform -1 0 14260 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_124
timestamp 1624635492
transform 1 0 12512 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 16468 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 14352 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 14996 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_143
timestamp 1624635492
transform 1 0 14260 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_147
timestamp 1624635492
transform 1 0 14628 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 18492 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1624635492
transform -1 0 16836 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1624635492
transform 1 0 16468 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_172
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1624635492
transform -1 0 18768 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform 1 0 18952 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 19228 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1624635492
transform -1 0 22080 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624635492
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_218
timestamp 1624635492
transform 1 0 21160 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1624635492
transform -1 0 23000 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 23460 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_238
timestamp 1624635492
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1624635492
transform 1 0 2852 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1624635492
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1624635492
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1624635492
transform -1 0 8280 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_54
timestamp 1624635492
transform 1 0 6072 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_78
timestamp 1624635492
transform 1 0 8280 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1624635492
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_87
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1624635492
transform -1 0 11224 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1624635492
transform -1 0 12696 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1624635492
transform 1 0 9660 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1624635492
transform 1 0 12788 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_126
timestamp 1624635492
transform 1 0 12696 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 15364 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_153
timestamp 1624635492
transform 1 0 15180 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1624635492
transform -1 0 17664 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform -1 0 18032 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_180
timestamp 1624635492
transform 1 0 17664 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 18032 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 21252 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624635492
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 21252 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1624635492
transform 1 0 22724 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 23460 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_238
timestamp 1624635492
transform 1 0 23000 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 2024 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_9
timestamp 1624635492
transform 1 0 1932 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 3772 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_26
timestamp 1624635492
transform 1 0 3496 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1624635492
transform 1 0 4048 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1624635492
transform 1 0 5152 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1624635492
transform 1 0 6992 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_56
timestamp 1624635492
transform 1 0 6256 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_58
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1624635492
transform 1 0 8556 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_80
timestamp 1624635492
transform 1 0 8464 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1624635492
transform -1 0 10948 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 11224 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_97
timestamp 1624635492
transform 1 0 10028 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_110
timestamp 1624635492
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1624635492
transform -1 0 13524 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1624635492
transform 1 0 13524 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_17_115
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1624635492
transform -1 0 16468 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1624635492
transform -1 0 17756 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform -1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624635492
transform -1 0 16836 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1624635492
transform 1 0 16468 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1624635492
transform 1 0 19504 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1624635492
transform 1 0 19872 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 19504 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_203
timestamp 1624635492
transform 1 0 19780 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 20148 0 1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624635492
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 22172 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 23460 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_238
timestamp 1624635492
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1624635492
transform -1 0 3680 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_15
timestamp 1624635492
transform 1 0 2484 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_28
timestamp 1624635492
transform 1 0 3680 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1624635492
transform 1 0 5336 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform 1 0 6900 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_62
timestamp 1624635492
transform 1 0 6808 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1624635492
transform -1 0 9936 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1624635492
transform -1 0 8924 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 8372 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1624635492
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1624635492
transform -1 0 10304 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1624635492
transform -1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1624635492
transform 1 0 10580 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_96
timestamp 1624635492
transform 1 0 9936 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 12236 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_18_119
timestamp 1624635492
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1624635492
transform -1 0 15456 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_ltile_clb_mode__0.clb_clk
timestamp 1624635492
transform -1 0 15732 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 15916 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1624635492
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16744 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1624635492
transform 1 0 16744 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1624635492
transform -1 0 18400 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1624635492
transform -1 0 19228 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1624635492
transform 1 0 19596 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 19504 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624635492
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 22080 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_4  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 23184 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 23460 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1624635492
transform -1 0 3772 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 2576 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_15
timestamp 1624635492
transform 1 0 2484 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_15
timestamp 1624635492
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_19
timestamp 1624635492
transform 1 0 2852 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform 1 0 4048 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1624635492
transform 1 0 4692 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1624635492
transform 1 0 5520 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1624635492
transform 1 0 6164 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1624635492
transform -1 0 7912 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 7360 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 6992 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_67
timestamp 1624635492
transform 1 0 7268 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1624635492
transform -1 0 9936 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1624635492
transform 1 0 9384 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 9384 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1624635492
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1624635492
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1624635492
transform 1 0 10212 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform -1 0 10212 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1624635492
transform 1 0 11040 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_99
timestamp 1624635492
transform 1 0 10212 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 12788 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1624635492
transform -1 0 14260 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1624635492
transform 1 0 13340 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1624635492
transform -1 0 13340 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1624635492
transform -1 0 16284 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1624635492
transform -1 0 17756 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1624635492
transform 1 0 16008 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1624635492
transform 1 0 17480 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17756 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 16560 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_160
timestamp 1624635492
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1624635492
transform 1 0 19228 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform 1 0 19596 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1624635492
transform 1 0 18952 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__sdfxtp_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 19964 0 -1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624635492
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_199
timestamp 1624635492
transform 1 0 19412 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_204
timestamp 1624635492
transform 1 0 19872 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1624635492
transform 1 0 21804 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform -1 0 20332 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 21988 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 21804 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624635492
transform 1 0 22080 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1624635492
transform 1 0 22816 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1624635492
transform -1 0 23000 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 23460 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 23460 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_238
timestamp 1624635492
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_239
timestamp 1624635492
transform 1 0 23092 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1624635492
transform -1 0 3680 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1624635492
transform -1 0 2852 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1624635492
transform 1 0 3680 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1624635492
transform -1 0 5796 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform -1 0 4784 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1624635492
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1624635492
transform -1 0 6072 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8832 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_54
timestamp 1624635492
transform 1 0 6072 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_58
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_66
timestamp 1624635492
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9660 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _60_
timestamp 1624635492
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9660 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1624635492
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 13524 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 13156 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 16008 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.clb_clk
timestamp 1624635492
transform -1 0 15640 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1624635492
transform 1 0 16928 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17848 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 16008 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_181
timestamp 1624635492
transform 1 0 17756 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 19780 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1624635492
transform -1 0 19780 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 20608 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624635492
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 22172 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 23460 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1624635492
transform -1 0 3220 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1624635492
transform -1 0 4140 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1624635492
transform 1 0 4600 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_23
timestamp 1624635492
transform 1 0 3220 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_33
timestamp 1624635492
transform 1 0 4140 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_37
timestamp 1624635492
transform 1 0 4508 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_6  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform 1 0 6072 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7176 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 6900 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform -1 0 9384 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform -1 0 9016 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10856 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_82
timestamp 1624635492
transform 1 0 8648 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1624635492
transform -1 0 11684 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1624635492
transform -1 0 12512 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1624635492
transform 1 0 12512 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1624635492
transform -1 0 14260 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_22_133
timestamp 1624635492
transform 1 0 13340 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1624635492
transform -1 0 14996 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1624635492
transform 1 0 14996 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_ltile_clb_mode__0.clb_clk
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_147
timestamp 1624635492
transform 1 0 14628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1624635492
transform 1 0 16468 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1624635492
transform -1 0 19044 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 17940 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1624635492
transform -1 0 20424 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624635492
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1624635492
transform -1 0 19504 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 19228 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 22724 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 21252 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform 1 0 22724 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 23460 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_238
timestamp 1624635492
transform 1 0 23000 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1624635492
transform 1 0 2024 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1624635492
transform 1 0 1380 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1624635492
transform 1 0 1932 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1624635492
transform 1 0 4968 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1624635492
transform 1 0 3496 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1624635492
transform -1 0 8096 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1624635492
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform -1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 10120 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9292 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_79
timestamp 1624635492
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10120 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1624635492
transform 1 0 12512 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 11684 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 13064 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_23_129
timestamp 1624635492
transform 1 0 12972 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 15732 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1624635492
transform 1 0 14536 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 15732 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_155
timestamp 1624635492
transform 1 0 15364 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1624635492
transform 1 0 16560 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform 1 0 17112 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624635492
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_172
timestamp 1624635492
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 18400 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 19872 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1624635492
transform 1 0 18124 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 18124 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1624635492
transform -1 0 22080 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform 1 0 21344 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624635492
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_223
timestamp 1624635492
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 23000 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 23460 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_238
timestamp 1624635492
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1624635492
transform -1 0 3772 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1624635492
transform 1 0 1472 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1624635492
transform 1 0 1380 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1624635492
transform 1 0 5336 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1624635492
transform 1 0 6808 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform -1 0 8556 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 8832 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 9936 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1624635492
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 10764 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10764 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 12236 0 -1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 15824 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_142
timestamp 1624635492
transform 1 0 14168 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 17296 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform -1 0 18952 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 17480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 21068 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624635492
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1624635492
transform -1 0 19504 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1624635492
transform -1 0 19228 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 21252 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform -1 0 23000 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 23460 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_238
timestamp 1624635492
transform 1 0 23000 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1624635492
transform 1 0 2024 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output45
timestamp 1624635492
transform -1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_7
timestamp 1624635492
transform 1 0 1748 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1624635492
transform 1 0 4692 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1624635492
transform -1 0 4692 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_26
timestamp 1624635492
transform 1 0 3496 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1624635492
transform -1 0 6348 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1624635492
transform -1 0 6900 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6900 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8372 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 9384 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _63_
timestamp 1624635492
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _61_
timestamp 1624635492
transform -1 0 11960 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12144 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14444 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _62_
timestamp 1624635492
transform -1 0 14720 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 14904 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform 1 0 16928 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1624635492
transform 1 0 17572 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624635492
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1624635492
transform 1 0 17296 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_175
timestamp 1624635492
transform 1 0 17204 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1624635492
transform -1 0 20240 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform -1 0 19412 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_195
timestamp 1624635492
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1624635492
transform -1 0 21068 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1624635492
transform -1 0 21896 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624635492
transform 1 0 22080 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_226
timestamp 1624635492
transform 1 0 21896 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1624635492
transform -1 0 23000 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 23460 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_238
timestamp 1624635492
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform 1 0 1564 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1624635492
transform -1 0 3220 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1624635492
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_21
timestamp 1624635492
transform 1 0 3036 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1624635492
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1624635492
transform 1 0 4508 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 4784 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 6256 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1624635492
transform -1 0 4692 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 4232 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_30
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_39
timestamp 1624635492
transform 1 0 4692 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 6624 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 7452 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_56
timestamp 1624635492
transform 1 0 6256 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_67
timestamp 1624635492
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform 1 0 9384 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8924 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 8280 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 8280 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1624635492
transform 1 0 8924 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11132 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10028 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11132 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624635492
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 10028 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 11500 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_106
timestamp 1624635492
transform 1 0 10856 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1624635492
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 12604 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 11960 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 13432 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_26_137
timestamp 1624635492
transform 1 0 13708 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_115
timestamp 1624635492
transform 1 0 11684 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1624635492
transform -1 0 15180 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1624635492
transform -1 0 16376 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16008 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1624635492
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 16560 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624635492
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_178
timestamp 1624635492
transform 1 0 17480 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 17112 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1624635492
transform 1 0 17112 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1624635492
transform 1 0 17388 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1624635492
transform 1 0 17664 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1624635492
transform -1 0 19044 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 17480 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1624635492
transform -1 0 19964 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1624635492
transform 1 0 19964 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1624635492
transform 1 0 19596 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1624635492
transform -1 0 19504 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624635492
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform -1 0 19228 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1624635492
transform 1 0 20424 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1624635492
transform 1 0 20976 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform -1 0 22080 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 21436 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624635492
transform 1 0 22080 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_219
timestamp 1624635492
transform 1 0 21252 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_214
timestamp 1624635492
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1624635492
transform 1 0 22172 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform 1 0 22908 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 23460 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 23460 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_238
timestamp 1624635492
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1624635492
transform 1 0 2116 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1624635492
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1624635492
transform 1 0 3864 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 6256 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624635492
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1624635492
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_39
timestamp 1624635492
transform 1 0 4692 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8372 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 6440 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_56
timestamp 1624635492
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_61
timestamp 1624635492
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624635492
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_79
timestamp 1624635492
transform 1 0 8372 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1624635492
transform 1 0 8740 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11500 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_96
timestamp 1624635492
transform 1 0 9936 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_113
timestamp 1624635492
transform 1 0 11500 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12788 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__S
timestamp 1624635492
transform -1 0 13800 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_117
timestamp 1624635492
transform 1 0 11868 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1624635492
transform 1 0 14352 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624635492
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_138
timestamp 1624635492
transform 1 0 13800 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_142
timestamp 1624635492
transform 1 0 14168 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1624635492
transform -1 0 17296 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1624635492
transform -1 0 17572 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1624635492
transform -1 0 17848 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 18032 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1624635492
transform 1 0 18032 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1624635492
transform -1 0 21068 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624635492
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1624635492
transform -1 0 21344 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1624635492
transform 1 0 21344 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 23184 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 23460 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1624635492
transform -1 0 2208 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1624635492
transform -1 0 3680 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1624635492
transform 1 0 3680 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1624635492
transform -1 0 4784 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 4784 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1624635492
transform 1 0 6900 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform -1 0 9108 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1624635492
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_56
timestamp 1624635492
transform 1 0 6256 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_58
timestamp 1624635492
transform 1 0 6440 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_62
timestamp 1624635492
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1624635492
transform -1 0 9660 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_89
timestamp 1624635492
transform 1 0 9292 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform -1 0 11592 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1624635492
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1624635492
transform -1 0 13156 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 13340 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_133
timestamp 1624635492
transform 1 0 13340 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13892 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1624635492
transform -1 0 16192 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18308 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1624635492
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 16468 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 17480 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 17296 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_167
timestamp 1624635492
transform 1 0 16468 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_172
timestamp 1624635492
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1624635492
transform 1 0 18676 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform 1 0 18400 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_187
timestamp 1624635492
transform 1 0 18308 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1624635492
transform -1 0 20424 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1624635492
transform 1 0 20608 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1624635492
transform 1 0 22080 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1624635492
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1624635492
transform 1 0 22172 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 23460 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_238
timestamp 1624635492
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1624635492
transform -1 0 3220 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1624635492
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1624635492
transform 1 0 5244 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1624635492
transform -1 0 4692 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform -1 0 5060 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_23
timestamp 1624635492
transform 1 0 3220 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_39
timestamp 1624635492
transform 1 0 4692 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_43
timestamp 1624635492
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 8188 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 6348 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_57
timestamp 1624635492
transform 1 0 6348 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 9108 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1624635492
transform -1 0 9016 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 11040 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1624635492
transform -1 0 14260 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1624635492
transform 1 0 11868 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_133
timestamp 1624635492
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform -1 0 14628 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1624635492
transform -1 0 14904 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1624635492
transform 1 0 14904 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1624635492
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 16652 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_166
timestamp 1624635492
transform 1 0 16376 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1624635492
transform -1 0 19412 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1624635492
transform 1 0 19596 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1624635492
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_199
timestamp 1624635492
transform 1 0 19412 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1624635492
transform 1 0 21068 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 23460 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_233
timestamp 1624635492
transform 1 0 22540 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_239
timestamp 1624635492
transform 1 0 23092 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1624635492
transform -1 0 3956 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1624635492
transform 1 0 1656 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1624635492
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1624635492
transform 1 0 4784 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1624635492
transform 1 0 3956 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform -1 0 5888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 6164 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 7268 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1624635492
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_55
timestamp 1624635492
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_67
timestamp 1624635492
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1624635492
transform 1 0 7452 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 9660 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11316 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1624635492
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1624635492
transform -1 0 11592 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_92
timestamp 1624635492
transform 1 0 9568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1624635492
transform -1 0 13984 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1624635492
transform 1 0 11684 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1624635492
transform 1 0 14812 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1624635492
transform 1 0 15640 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1624635492
transform -1 0 14812 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1624635492
transform -1 0 16836 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 18400 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1624635492
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1624635492
transform 1 0 16468 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1624635492
transform -1 0 19872 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1624635492
transform 1 0 19872 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_188
timestamp 1624635492
transform 1 0 18400 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_194
timestamp 1624635492
transform 1 0 18952 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1624635492
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1624635492
transform 1 0 21620 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1624635492
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1624635492
transform 1 0 22172 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 23460 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1624635492
transform -1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1624635492
transform -1 0 3036 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1624635492
transform -1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1624635492
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1624635492
transform 1 0 3864 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1624635492
transform -1 0 5520 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1624635492
transform -1 0 3772 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1624635492
transform -1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1624635492
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1624635492
transform -1 0 6348 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform 1 0 6348 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8556 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1624635492
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_62
timestamp 1624635492
transform 1 0 6808 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1624635492
transform -1 0 8832 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1624635492
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0__SCE
timestamp 1624635492
transform -1 0 9292 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1624635492
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_89
timestamp 1624635492
transform 1 0 9292 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9660 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1624635492
transform 1 0 11132 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1624635492
transform -1 0 13340 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1624635492
transform -1 0 14168 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1624635492
transform -1 0 12512 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 12144 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_120
timestamp 1624635492
transform 1 0 12144 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1624635492
transform -1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform -1 0 16008 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1624635492
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1624635492
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 15732 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_142
timestamp 1624635492
transform 1 0 14168 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_144
timestamp 1624635492
transform 1 0 14352 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 17112 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16836 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 19044 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 17296 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624635492
transform -1 0 17480 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_178
timestamp 1624635492
transform 1 0 17480 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1624635492
transform -1 0 20424 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1624635492
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_195
timestamp 1624635492
transform 1 0 19044 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1624635492
transform 1 0 19412 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1624635492
transform 1 0 20976 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1624635492
transform -1 0 20976 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 20700 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_210
timestamp 1624635492
transform 1 0 20424 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1624635492
transform -1 0 22724 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 23460 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output54
timestamp 1624635492
transform 1 0 22816 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_235
timestamp 1624635492
transform 1 0 22724 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1624635492
transform -1 0 2024 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1624635492
transform -1 0 3864 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1624635492
transform 1 0 1564 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1624635492
transform 1 0 2024 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1624635492
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1624635492
transform -1 0 1748 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1624635492
transform -1 0 1564 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1624635492
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1624635492
transform 1 0 3496 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1624635492
transform -1 0 4692 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1624635492
transform -1 0 5520 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1624635492
transform 1 0 3864 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1624635492
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1624635492
transform -1 0 6716 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform 1 0 6716 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 5336 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 6348 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6808 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 7176 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1624635492
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 7176 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1624635492
transform 1 0 8280 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_85
timestamp 1624635492
transform 1 0 8924 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 9200 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 9292 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 9016 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1624635492
transform 1 0 8556 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1624635492
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform -1 0 8924 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9292 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10672 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1624635492
transform 1 0 10764 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1624635492
transform 1 0 11040 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11500 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1624635492
transform -1 0 12972 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1624635492
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 11500 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_113
timestamp 1624635492
transform 1 0 11500 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1624635492
transform -1 0 13800 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform 1 0 13340 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1624635492
transform -1 0 13156 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 13340 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1624635492
transform 1 0 13892 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1624635492
transform -1 0 15548 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1624635492
transform -1 0 16376 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 14168 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1624635492
transform 1 0 14352 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1624635492
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_142
timestamp 1624635492
transform 1 0 14168 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1624635492
transform -1 0 17204 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform 1 0 16376 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15824 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17296 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 18768 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1624635492
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 16836 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_175
timestamp 1624635492
transform 1 0 17204 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1624635492
transform 1 0 18768 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1624635492
transform 1 0 19044 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 19596 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 19596 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1624635492
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1624635492
transform 1 0 19320 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1624635492
transform -1 0 19780 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_203
timestamp 1624635492
transform 1 0 19780 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1624635492
transform -1 0 20608 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_211
timestamp 1624635492
transform 1 0 20516 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1624635492
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1624635492
transform 1 0 20792 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1624635492
transform -1 0 20792 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 20976 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1624635492
transform -1 0 21252 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1624635492
transform -1 0 21528 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1624635492
transform -1 0 21252 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1624635492
transform -1 0 21528 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1624635492
transform -1 0 21804 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1624635492
transform -1 0 21804 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform 1 0 22080 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1624635492
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1624635492
transform -1 0 22080 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1624635492
transform -1 0 22080 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform 1 0 22356 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 23460 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1624635492
transform -1 0 23460 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output56
timestamp 1624635492
transform 1 0 22816 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output58
timestamp 1624635492
transform 1 0 22448 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 22356 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1624635492
transform 1 0 1840 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1624635492
transform 1 0 2116 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1624635492
transform 1 0 2576 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1624635492
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform -1 0 1656 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 1840 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1624635492
transform 1 0 2392 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1624635492
transform 1 0 4048 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 4416 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_35
timestamp 1624635492
transform 1 0 4324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform -1 0 6716 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1624635492
transform -1 0 6348 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8372 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1624635492
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 6900 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 10856 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_6  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1624635492
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 9384 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform 1 0 11040 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1624635492
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1624635492
transform 1 0 11316 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 11040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1624635492
transform 1 0 11776 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1624635492
transform 1 0 13248 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_115
timestamp 1624635492
transform 1 0 11684 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1624635492
transform 1 0 14720 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1624635492
transform 1 0 16192 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16928 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1624635492
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 16836 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 16652 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_6  clk_0_FTB00
timestamp 1624635492
transform 1 0 18400 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform 1 0 19228 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output69_A
timestamp 1624635492
transform 1 0 19688 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1624635492
transform -1 0 20056 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_201
timestamp 1624635492
transform 1 0 19596 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_208
timestamp 1624635492
transform 1 0 20240 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output71_A
timestamp 1624635492
transform 1 0 20056 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_215
timestamp 1624635492
transform 1 0 20884 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_212
timestamp 1624635492
transform 1 0 20608 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output73_A
timestamp 1624635492
transform 1 0 20700 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_219
timestamp 1624635492
transform 1 0 21252 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1624635492
transform -1 0 21528 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_222
timestamp 1624635492
transform 1 0 21528 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output81_A
timestamp 1624635492
transform 1 0 21896 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1624635492
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1624635492
transform -1 0 23460 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output60
timestamp 1624635492
transform 1 0 22816 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform 1 0 22448 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1624635492
transform -1 0 22356 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_231
timestamp 1624635492
transform 1 0 22356 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1624635492
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output70
timestamp 1624635492
transform -1 0 1748 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform -1 0 2116 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform -1 0 2484 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform -1 0 2852 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform -1 0 3220 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1624635492
transform -1 0 3772 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1624635492
transform 1 0 5152 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1624635492
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform -1 0 4232 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform -1 0 4600 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform -1 0 5152 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 4784 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1624635492
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_25
timestamp 1624635492
transform 1 0 3404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1624635492
transform 1 0 5796 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1624635492
transform -1 0 5796 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1624635492
transform 1 0 6440 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1624635492
transform -1 0 6348 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1624635492
transform 1 0 6532 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1624635492
transform 1 0 6808 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1624635492
transform 1 0 7176 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_57
timestamp 1624635492
transform 1 0 6348 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_65
timestamp 1624635492
transform 1 0 7084 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1624635492
transform 1 0 9200 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9476 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 8280 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 9108 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1624635492
transform 1 0 9108 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11408 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1624635492
transform -1 0 11776 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1624635492
transform 1 0 13340 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1624635492
transform 1 0 11776 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1624635492
transform 1 0 11868 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1624635492
transform 1 0 12512 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1624635492
transform -1 0 13340 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1624635492
transform 1 0 12144 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1624635492
transform -1 0 13064 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_123
timestamp 1624635492
transform 1 0 12420 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1624635492
transform 1 0 14536 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1624635492
transform -1 0 15640 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1624635492
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1624635492
transform 1 0 14168 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1624635492
transform 1 0 14812 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1624635492
transform 1 0 15640 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_152
timestamp 1624635492
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_4  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1624635492
transform -1 0 18492 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1624635492
transform 1 0 17112 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1624635492
transform 1 0 16836 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1624635492
transform -1 0 16836 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1624635492
transform 1 0 15916 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1624635492
transform -1 0 16560 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 17388 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_164
timestamp 1624635492
transform 1 0 16192 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1624635492
transform 1 0 19780 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output43
timestamp 1624635492
transform -1 0 18860 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output69
timestamp 1624635492
transform -1 0 20240 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform 1 0 19412 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform 1 0 19044 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 19044 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  output50
timestamp 1624635492
transform -1 0 20884 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output64
timestamp 1624635492
transform 1 0 22080 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output66
timestamp 1624635492
transform 1 0 21712 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output68
timestamp 1624635492
transform 1 0 21344 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output71
timestamp 1624635492
transform -1 0 20608 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform -1 0 21252 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_219
timestamp 1624635492
transform 1 0 21252 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1624635492
transform -1 0 23460 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1624635492
transform 1 0 22448 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output62
timestamp 1624635492
transform 1 0 22816 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_233
timestamp 1624635492
transform 1 0 22540 0 -1 22304
box -38 -48 314 592
<< labels >>
rlabel metal2 s 17038 23800 17094 24600 6 SC_IN_TOP
port 0 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal2 s 17682 23800 17738 24600 6 SC_OUT_TOP
port 2 nsew signal tristate
rlabel metal3 s 23800 6808 24600 6928 6 Test_en_E_in
port 3 nsew signal input
rlabel metal3 s 23800 6264 24600 6384 6 Test_en_E_out
port 4 nsew signal tristate
rlabel metal3 s 0 21360 800 21480 6 Test_en_W_in
port 5 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 Test_en_W_out
port 6 nsew signal tristate
rlabel metal2 s 2042 0 2098 800 6 bottom_width_0_height_0__pin_50_
port 7 nsew signal tristate
rlabel metal2 s 6090 0 6146 800 6 bottom_width_0_height_0__pin_51_
port 8 nsew signal tristate
rlabel metal3 s 0 9120 800 9240 6 ccff_head
port 9 nsew signal input
rlabel metal3 s 23800 5584 24600 5704 6 ccff_tail
port 10 nsew signal tristate
rlabel metal2 s 18326 23800 18382 24600 6 clk_0_N_in
port 11 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 clk_0_S_in
port 12 nsew signal input
rlabel metal3 s 23800 8168 24600 8288 6 prog_clk_0_E_out
port 13 nsew signal tristate
rlabel metal3 s 23800 7488 24600 7608 6 prog_clk_0_N_in
port 14 nsew signal input
rlabel metal2 s 18970 23800 19026 24600 6 prog_clk_0_N_out
port 15 nsew signal tristate
rlabel metal2 s 18418 0 18474 800 6 prog_clk_0_S_in
port 16 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 prog_clk_0_S_out
port 17 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 prog_clk_0_W_out
port 18 nsew signal tristate
rlabel metal3 s 23800 8848 24600 8968 6 right_width_0_height_0__pin_16_
port 19 nsew signal input
rlabel metal3 s 23800 9528 24600 9648 6 right_width_0_height_0__pin_17_
port 20 nsew signal input
rlabel metal3 s 23800 10208 24600 10328 6 right_width_0_height_0__pin_18_
port 21 nsew signal input
rlabel metal3 s 23800 10888 24600 11008 6 right_width_0_height_0__pin_19_
port 22 nsew signal input
rlabel metal3 s 23800 11568 24600 11688 6 right_width_0_height_0__pin_20_
port 23 nsew signal input
rlabel metal3 s 23800 12248 24600 12368 6 right_width_0_height_0__pin_21_
port 24 nsew signal input
rlabel metal3 s 23800 12792 24600 12912 6 right_width_0_height_0__pin_22_
port 25 nsew signal input
rlabel metal3 s 23800 13472 24600 13592 6 right_width_0_height_0__pin_23_
port 26 nsew signal input
rlabel metal3 s 23800 14152 24600 14272 6 right_width_0_height_0__pin_24_
port 27 nsew signal input
rlabel metal3 s 23800 14832 24600 14952 6 right_width_0_height_0__pin_25_
port 28 nsew signal input
rlabel metal3 s 23800 15512 24600 15632 6 right_width_0_height_0__pin_26_
port 29 nsew signal input
rlabel metal3 s 23800 16192 24600 16312 6 right_width_0_height_0__pin_27_
port 30 nsew signal input
rlabel metal3 s 23800 16872 24600 16992 6 right_width_0_height_0__pin_28_
port 31 nsew signal input
rlabel metal3 s 23800 17552 24600 17672 6 right_width_0_height_0__pin_29_
port 32 nsew signal input
rlabel metal3 s 23800 18232 24600 18352 6 right_width_0_height_0__pin_30_
port 33 nsew signal input
rlabel metal3 s 23800 18776 24600 18896 6 right_width_0_height_0__pin_31_
port 34 nsew signal input
rlabel metal3 s 23800 280 24600 400 6 right_width_0_height_0__pin_42_lower
port 35 nsew signal tristate
rlabel metal3 s 23800 19456 24600 19576 6 right_width_0_height_0__pin_42_upper
port 36 nsew signal tristate
rlabel metal3 s 23800 824 24600 944 6 right_width_0_height_0__pin_43_lower
port 37 nsew signal tristate
rlabel metal3 s 23800 20136 24600 20256 6 right_width_0_height_0__pin_43_upper
port 38 nsew signal tristate
rlabel metal3 s 23800 1504 24600 1624 6 right_width_0_height_0__pin_44_lower
port 39 nsew signal tristate
rlabel metal3 s 23800 20816 24600 20936 6 right_width_0_height_0__pin_44_upper
port 40 nsew signal tristate
rlabel metal3 s 23800 2184 24600 2304 6 right_width_0_height_0__pin_45_lower
port 41 nsew signal tristate
rlabel metal3 s 23800 21496 24600 21616 6 right_width_0_height_0__pin_45_upper
port 42 nsew signal tristate
rlabel metal3 s 23800 2864 24600 2984 6 right_width_0_height_0__pin_46_lower
port 43 nsew signal tristate
rlabel metal3 s 23800 22176 24600 22296 6 right_width_0_height_0__pin_46_upper
port 44 nsew signal tristate
rlabel metal3 s 23800 3544 24600 3664 6 right_width_0_height_0__pin_47_lower
port 45 nsew signal tristate
rlabel metal3 s 23800 22856 24600 22976 6 right_width_0_height_0__pin_47_upper
port 46 nsew signal tristate
rlabel metal3 s 23800 4224 24600 4344 6 right_width_0_height_0__pin_48_lower
port 47 nsew signal tristate
rlabel metal3 s 23800 23536 24600 23656 6 right_width_0_height_0__pin_48_upper
port 48 nsew signal tristate
rlabel metal3 s 23800 4904 24600 5024 6 right_width_0_height_0__pin_49_lower
port 49 nsew signal tristate
rlabel metal3 s 23800 24216 24600 24336 6 right_width_0_height_0__pin_49_upper
port 50 nsew signal tristate
rlabel metal2 s 5446 23800 5502 24600 6 top_width_0_height_0__pin_0_
port 51 nsew signal input
rlabel metal2 s 11886 23800 11942 24600 6 top_width_0_height_0__pin_10_
port 52 nsew signal input
rlabel metal2 s 12530 23800 12586 24600 6 top_width_0_height_0__pin_11_
port 53 nsew signal input
rlabel metal2 s 13174 23800 13230 24600 6 top_width_0_height_0__pin_12_
port 54 nsew signal input
rlabel metal2 s 13818 23800 13874 24600 6 top_width_0_height_0__pin_13_
port 55 nsew signal input
rlabel metal2 s 14462 23800 14518 24600 6 top_width_0_height_0__pin_14_
port 56 nsew signal input
rlabel metal2 s 15106 23800 15162 24600 6 top_width_0_height_0__pin_15_
port 57 nsew signal input
rlabel metal2 s 6090 23800 6146 24600 6 top_width_0_height_0__pin_1_
port 58 nsew signal input
rlabel metal2 s 6734 23800 6790 24600 6 top_width_0_height_0__pin_2_
port 59 nsew signal input
rlabel metal2 s 15750 23800 15806 24600 6 top_width_0_height_0__pin_32_
port 60 nsew signal input
rlabel metal2 s 16394 23800 16450 24600 6 top_width_0_height_0__pin_33_
port 61 nsew signal input
rlabel metal2 s 19614 23800 19670 24600 6 top_width_0_height_0__pin_34_lower
port 62 nsew signal tristate
rlabel metal2 s 294 23800 350 24600 6 top_width_0_height_0__pin_34_upper
port 63 nsew signal tristate
rlabel metal2 s 20258 23800 20314 24600 6 top_width_0_height_0__pin_35_lower
port 64 nsew signal tristate
rlabel metal2 s 938 23800 994 24600 6 top_width_0_height_0__pin_35_upper
port 65 nsew signal tristate
rlabel metal2 s 20902 23800 20958 24600 6 top_width_0_height_0__pin_36_lower
port 66 nsew signal tristate
rlabel metal2 s 1582 23800 1638 24600 6 top_width_0_height_0__pin_36_upper
port 67 nsew signal tristate
rlabel metal2 s 21546 23800 21602 24600 6 top_width_0_height_0__pin_37_lower
port 68 nsew signal tristate
rlabel metal2 s 2226 23800 2282 24600 6 top_width_0_height_0__pin_37_upper
port 69 nsew signal tristate
rlabel metal2 s 22190 23800 22246 24600 6 top_width_0_height_0__pin_38_lower
port 70 nsew signal tristate
rlabel metal2 s 2870 23800 2926 24600 6 top_width_0_height_0__pin_38_upper
port 71 nsew signal tristate
rlabel metal2 s 22834 23800 22890 24600 6 top_width_0_height_0__pin_39_lower
port 72 nsew signal tristate
rlabel metal2 s 3514 23800 3570 24600 6 top_width_0_height_0__pin_39_upper
port 73 nsew signal tristate
rlabel metal2 s 7378 23800 7434 24600 6 top_width_0_height_0__pin_3_
port 74 nsew signal input
rlabel metal2 s 23478 23800 23534 24600 6 top_width_0_height_0__pin_40_lower
port 75 nsew signal tristate
rlabel metal2 s 4158 23800 4214 24600 6 top_width_0_height_0__pin_40_upper
port 76 nsew signal tristate
rlabel metal2 s 24122 23800 24178 24600 6 top_width_0_height_0__pin_41_lower
port 77 nsew signal tristate
rlabel metal2 s 4802 23800 4858 24600 6 top_width_0_height_0__pin_41_upper
port 78 nsew signal tristate
rlabel metal2 s 8022 23800 8078 24600 6 top_width_0_height_0__pin_4_
port 79 nsew signal input
rlabel metal2 s 8666 23800 8722 24600 6 top_width_0_height_0__pin_5_
port 80 nsew signal input
rlabel metal2 s 9310 23800 9366 24600 6 top_width_0_height_0__pin_6_
port 81 nsew signal input
rlabel metal2 s 9954 23800 10010 24600 6 top_width_0_height_0__pin_7_
port 82 nsew signal input
rlabel metal2 s 10598 23800 10654 24600 6 top_width_0_height_0__pin_8_
port 83 nsew signal input
rlabel metal2 s 11242 23800 11298 24600 6 top_width_0_height_0__pin_9_
port 84 nsew signal input
rlabel metal4 s 19604 2128 19924 22352 6 VPWR
port 85 nsew power bidirectional
rlabel metal4 s 12140 2128 12460 22352 6 VPWR
port 86 nsew power bidirectional
rlabel metal4 s 4676 2128 4996 22352 6 VPWR
port 87 nsew power bidirectional
rlabel metal4 s 15872 2128 16192 22352 6 VGND
port 88 nsew ground bidirectional
rlabel metal4 s 8408 2128 8728 22352 6 VGND
port 89 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 24600 24600
<< end >>
